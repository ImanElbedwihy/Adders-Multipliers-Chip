module alu_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [15:0] A;
   input [15:0] B;
   input CI;
   output [15:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [15:1] carry;

   FA1DHD U1_0 (.S(SUM[0]), 
	.CO(carry[1]), 
	.CI(n1), 
	.B(B[0]), 
	.A(A[0]));
   FA1DHD U1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.CI(carry[1]), 
	.B(B[1]), 
	.A(A[1]));
   FA1DHD U1_13 (.S(SUM[13]), 
	.CO(carry[14]), 
	.CI(carry[13]), 
	.B(B[13]), 
	.A(A[13]));
   FA1DHD U1_11 (.S(SUM[11]), 
	.CO(carry[12]), 
	.CI(carry[11]), 
	.B(B[11]), 
	.A(A[11]));
   FA1DHD U1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.CI(carry[7]), 
	.B(B[7]), 
	.A(A[7]));
   FA1DHD U1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(B[5]), 
	.A(A[5]));
   FA1DHD U1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(B[3]), 
	.A(A[3]));
   FA1DHD U1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(B[2]), 
	.A(A[2]));
   FA1DHD U1_9 (.S(SUM[9]), 
	.CO(carry[10]), 
	.CI(carry[9]), 
	.B(B[9]), 
	.A(A[9]));
   FA1DHD U1_14 (.S(SUM[14]), 
	.CO(carry[15]), 
	.CI(carry[14]), 
	.B(B[14]), 
	.A(A[14]));
   FA1DHD U1_12 (.S(SUM[12]), 
	.CO(carry[13]), 
	.CI(carry[12]), 
	.B(B[12]), 
	.A(A[12]));
   FA1DHD U1_10 (.S(SUM[10]), 
	.CO(carry[11]), 
	.CI(carry[10]), 
	.B(B[10]), 
	.A(A[10]));
   FA1DHD U1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.CI(carry[8]), 
	.B(B[8]), 
	.A(A[8]));
   FA1DHD U1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(B[6]), 
	.A(A[6]));
   FA1DHD U1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(B[4]), 
	.A(A[4]));
   XOR3EHD U1_15 (.O(SUM[15]), 
	.I3(carry[15]), 
	.I2(B[15]), 
	.I1(A[15]));
   TIE0DHD U1 (.O(n1));
endmodule

module alu_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [15:0] A;
   input [15:0] B;
   input CI;
   output [15:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire [16:0] carry;

   FA1DHD U2_0 (.S(DIFF[0]), 
	.CO(carry[1]), 
	.CI(n17), 
	.B(n16), 
	.A(A[0]));
   FA1DHD U2_1 (.S(DIFF[1]), 
	.CO(carry[2]), 
	.CI(carry[1]), 
	.B(n15), 
	.A(A[1]));
   FA1DHD U2_13 (.S(DIFF[13]), 
	.CO(carry[14]), 
	.CI(carry[13]), 
	.B(n3), 
	.A(A[13]));
   FA1DHD U2_11 (.S(DIFF[11]), 
	.CO(carry[12]), 
	.CI(carry[11]), 
	.B(n5), 
	.A(A[11]));
   FA1DHD U2_7 (.S(DIFF[7]), 
	.CO(carry[8]), 
	.CI(carry[7]), 
	.B(n9), 
	.A(A[7]));
   FA1DHD U2_5 (.S(DIFF[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(n11), 
	.A(A[5]));
   FA1DHD U2_3 (.S(DIFF[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(n13), 
	.A(A[3]));
   FA1DHD U2_2 (.S(DIFF[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(n14), 
	.A(A[2]));
   FA1DHD U2_9 (.S(DIFF[9]), 
	.CO(carry[10]), 
	.CI(carry[9]), 
	.B(n7), 
	.A(A[9]));
   FA1DHD U2_14 (.S(DIFF[14]), 
	.CO(carry[15]), 
	.CI(carry[14]), 
	.B(n2), 
	.A(A[14]));
   FA1DHD U2_12 (.S(DIFF[12]), 
	.CO(carry[13]), 
	.CI(carry[12]), 
	.B(n4), 
	.A(A[12]));
   FA1DHD U2_10 (.S(DIFF[10]), 
	.CO(carry[11]), 
	.CI(carry[10]), 
	.B(n6), 
	.A(A[10]));
   FA1DHD U2_8 (.S(DIFF[8]), 
	.CO(carry[9]), 
	.CI(carry[8]), 
	.B(n8), 
	.A(A[8]));
   FA1DHD U2_6 (.S(DIFF[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(n10), 
	.A(A[6]));
   FA1DHD U2_4 (.S(DIFF[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(n12), 
	.A(A[4]));
   XOR3EHD U2_15 (.O(DIFF[15]), 
	.I3(carry[15]), 
	.I2(n1), 
	.I1(A[15]));
   INVDHD U1 (.O(n1), 
	.I(B[15]));
   INVDHD U2 (.O(n12), 
	.I(B[4]));
   INVDHD U3 (.O(n10), 
	.I(B[6]));
   INVDHD U4 (.O(n8), 
	.I(B[8]));
   INVDHD U5 (.O(n6), 
	.I(B[10]));
   INVDHD U6 (.O(n4), 
	.I(B[12]));
   INVDHD U7 (.O(n2), 
	.I(B[14]));
   INVDHD U8 (.O(n7), 
	.I(B[9]));
   INVDHD U9 (.O(n14), 
	.I(B[2]));
   INVDHD U10 (.O(n13), 
	.I(B[3]));
   INVDHD U11 (.O(n11), 
	.I(B[5]));
   INVDHD U12 (.O(n9), 
	.I(B[7]));
   INVDHD U13 (.O(n5), 
	.I(B[11]));
   INVDHD U14 (.O(n3), 
	.I(B[13]));
   INVDHD U15 (.O(n15), 
	.I(B[1]));
   INVDHD U16 (.O(n16), 
	.I(B[0]));
   TIE1DHD U17 (.O(n17));
endmodule

module data_memory (
	clk, 
	mem_access_addr, 
	mem_write_data, 
	mem_write_en, 
	mem_read, 
	mem_read_data, 
	clk_m__L3_N1, 
	clk_m__L3_N10, 
	clk_m__L3_N100, 
	clk_m__L3_N101, 
	clk_m__L3_N102, 
	clk_m__L3_N103, 
	clk_m__L3_N104, 
	clk_m__L3_N105, 
	clk_m__L3_N106, 
	clk_m__L3_N107, 
	clk_m__L3_N108, 
	clk_m__L3_N109, 
	clk_m__L3_N11, 
	clk_m__L3_N110, 
	clk_m__L3_N111, 
	clk_m__L3_N112, 
	clk_m__L3_N113, 
	clk_m__L3_N114, 
	clk_m__L3_N115, 
	clk_m__L3_N116, 
	clk_m__L3_N117, 
	clk_m__L3_N118, 
	clk_m__L3_N119, 
	clk_m__L3_N12, 
	clk_m__L3_N120, 
	clk_m__L3_N121, 
	clk_m__L3_N122, 
	clk_m__L3_N123, 
	clk_m__L3_N124, 
	clk_m__L3_N125, 
	clk_m__L3_N126, 
	clk_m__L3_N127, 
	clk_m__L3_N128, 
	clk_m__L3_N129, 
	clk_m__L3_N13, 
	clk_m__L3_N130, 
	clk_m__L3_N131, 
	clk_m__L3_N132, 
	clk_m__L3_N133, 
	clk_m__L3_N134, 
	clk_m__L3_N135, 
	clk_m__L3_N136, 
	clk_m__L3_N137, 
	clk_m__L3_N138, 
	clk_m__L3_N139, 
	clk_m__L3_N14, 
	clk_m__L3_N140, 
	clk_m__L3_N141, 
	clk_m__L3_N142, 
	clk_m__L3_N143, 
	clk_m__L3_N144, 
	clk_m__L3_N145, 
	clk_m__L3_N146, 
	clk_m__L3_N147, 
	clk_m__L3_N148, 
	clk_m__L3_N149, 
	clk_m__L3_N15, 
	clk_m__L3_N150, 
	clk_m__L3_N151, 
	clk_m__L3_N152, 
	clk_m__L3_N153, 
	clk_m__L3_N154, 
	clk_m__L3_N155, 
	clk_m__L3_N156, 
	clk_m__L3_N157, 
	clk_m__L3_N158, 
	clk_m__L3_N159, 
	clk_m__L3_N16, 
	clk_m__L3_N160, 
	clk_m__L3_N161, 
	clk_m__L3_N162, 
	clk_m__L3_N163, 
	clk_m__L3_N164, 
	clk_m__L3_N165, 
	clk_m__L3_N166, 
	clk_m__L3_N167, 
	clk_m__L3_N168, 
	clk_m__L3_N169, 
	clk_m__L3_N17, 
	clk_m__L3_N170, 
	clk_m__L3_N171, 
	clk_m__L3_N172, 
	clk_m__L3_N173, 
	clk_m__L3_N174, 
	clk_m__L3_N175, 
	clk_m__L3_N176, 
	clk_m__L3_N177, 
	clk_m__L3_N18, 
	clk_m__L3_N19, 
	clk_m__L3_N2, 
	clk_m__L3_N20, 
	clk_m__L3_N21, 
	clk_m__L3_N22, 
	clk_m__L3_N23, 
	clk_m__L3_N24, 
	clk_m__L3_N25, 
	clk_m__L3_N26, 
	clk_m__L3_N27, 
	clk_m__L3_N28, 
	clk_m__L3_N29, 
	clk_m__L3_N3, 
	clk_m__L3_N30, 
	clk_m__L3_N31, 
	clk_m__L3_N32, 
	clk_m__L3_N33, 
	clk_m__L3_N34, 
	clk_m__L3_N35, 
	clk_m__L3_N36, 
	clk_m__L3_N37, 
	clk_m__L3_N38, 
	clk_m__L3_N39, 
	clk_m__L3_N4, 
	clk_m__L3_N40, 
	clk_m__L3_N41, 
	clk_m__L3_N42, 
	clk_m__L3_N43, 
	clk_m__L3_N44, 
	clk_m__L3_N45, 
	clk_m__L3_N46, 
	clk_m__L3_N47, 
	clk_m__L3_N48, 
	clk_m__L3_N49, 
	clk_m__L3_N5, 
	clk_m__L3_N50, 
	clk_m__L3_N52, 
	clk_m__L3_N53, 
	clk_m__L3_N54, 
	clk_m__L3_N55, 
	clk_m__L3_N56, 
	clk_m__L3_N57, 
	clk_m__L3_N58, 
	clk_m__L3_N59, 
	clk_m__L3_N6, 
	clk_m__L3_N60, 
	clk_m__L3_N61, 
	clk_m__L3_N62, 
	clk_m__L3_N63, 
	clk_m__L3_N64, 
	clk_m__L3_N65, 
	clk_m__L3_N66, 
	clk_m__L3_N67, 
	clk_m__L3_N68, 
	clk_m__L3_N69, 
	clk_m__L3_N7, 
	clk_m__L3_N70, 
	clk_m__L3_N71, 
	clk_m__L3_N72, 
	clk_m__L3_N73, 
	clk_m__L3_N74, 
	clk_m__L3_N75, 
	clk_m__L3_N76, 
	clk_m__L3_N77, 
	clk_m__L3_N78, 
	clk_m__L3_N79, 
	clk_m__L3_N8, 
	clk_m__L3_N80, 
	clk_m__L3_N81, 
	clk_m__L3_N82, 
	clk_m__L3_N83, 
	clk_m__L3_N84, 
	clk_m__L3_N85, 
	clk_m__L3_N86, 
	clk_m__L3_N87, 
	clk_m__L3_N88, 
	clk_m__L3_N89, 
	clk_m__L3_N9, 
	clk_m__L3_N90, 
	clk_m__L3_N91, 
	clk_m__L3_N92, 
	clk_m__L3_N93, 
	clk_m__L3_N94, 
	clk_m__L3_N95, 
	clk_m__L3_N96, 
	clk_m__L3_N97, 
	clk_m__L3_N98, 
	clk_m__L3_N99, 
	clk_m__N0);
   input clk;
   input [15:0] mem_access_addr;
   input [15:0] mem_write_data;
   input mem_write_en;
   input mem_read;
   output [15:0] mem_read_data;
   input clk_m__L3_N1;
   input clk_m__L3_N10;
   input clk_m__L3_N100;
   input clk_m__L3_N101;
   input clk_m__L3_N102;
   input clk_m__L3_N103;
   input clk_m__L3_N104;
   input clk_m__L3_N105;
   input clk_m__L3_N106;
   input clk_m__L3_N107;
   input clk_m__L3_N108;
   input clk_m__L3_N109;
   input clk_m__L3_N11;
   input clk_m__L3_N110;
   input clk_m__L3_N111;
   input clk_m__L3_N112;
   input clk_m__L3_N113;
   input clk_m__L3_N114;
   input clk_m__L3_N115;
   input clk_m__L3_N116;
   input clk_m__L3_N117;
   input clk_m__L3_N118;
   input clk_m__L3_N119;
   input clk_m__L3_N12;
   input clk_m__L3_N120;
   input clk_m__L3_N121;
   input clk_m__L3_N122;
   input clk_m__L3_N123;
   input clk_m__L3_N124;
   input clk_m__L3_N125;
   input clk_m__L3_N126;
   input clk_m__L3_N127;
   input clk_m__L3_N128;
   input clk_m__L3_N129;
   input clk_m__L3_N13;
   input clk_m__L3_N130;
   input clk_m__L3_N131;
   input clk_m__L3_N132;
   input clk_m__L3_N133;
   input clk_m__L3_N134;
   input clk_m__L3_N135;
   input clk_m__L3_N136;
   input clk_m__L3_N137;
   input clk_m__L3_N138;
   input clk_m__L3_N139;
   input clk_m__L3_N14;
   input clk_m__L3_N140;
   input clk_m__L3_N141;
   input clk_m__L3_N142;
   input clk_m__L3_N143;
   input clk_m__L3_N144;
   input clk_m__L3_N145;
   input clk_m__L3_N146;
   input clk_m__L3_N147;
   input clk_m__L3_N148;
   input clk_m__L3_N149;
   input clk_m__L3_N15;
   input clk_m__L3_N150;
   input clk_m__L3_N151;
   input clk_m__L3_N152;
   input clk_m__L3_N153;
   input clk_m__L3_N154;
   input clk_m__L3_N155;
   input clk_m__L3_N156;
   input clk_m__L3_N157;
   input clk_m__L3_N158;
   input clk_m__L3_N159;
   input clk_m__L3_N16;
   input clk_m__L3_N160;
   input clk_m__L3_N161;
   input clk_m__L3_N162;
   input clk_m__L3_N163;
   input clk_m__L3_N164;
   input clk_m__L3_N165;
   input clk_m__L3_N166;
   input clk_m__L3_N167;
   input clk_m__L3_N168;
   input clk_m__L3_N169;
   input clk_m__L3_N17;
   input clk_m__L3_N170;
   input clk_m__L3_N171;
   input clk_m__L3_N172;
   input clk_m__L3_N173;
   input clk_m__L3_N174;
   input clk_m__L3_N175;
   input clk_m__L3_N176;
   input clk_m__L3_N177;
   input clk_m__L3_N18;
   input clk_m__L3_N19;
   input clk_m__L3_N2;
   input clk_m__L3_N20;
   input clk_m__L3_N21;
   input clk_m__L3_N22;
   input clk_m__L3_N23;
   input clk_m__L3_N24;
   input clk_m__L3_N25;
   input clk_m__L3_N26;
   input clk_m__L3_N27;
   input clk_m__L3_N28;
   input clk_m__L3_N29;
   input clk_m__L3_N3;
   input clk_m__L3_N30;
   input clk_m__L3_N31;
   input clk_m__L3_N32;
   input clk_m__L3_N33;
   input clk_m__L3_N34;
   input clk_m__L3_N35;
   input clk_m__L3_N36;
   input clk_m__L3_N37;
   input clk_m__L3_N38;
   input clk_m__L3_N39;
   input clk_m__L3_N4;
   input clk_m__L3_N40;
   input clk_m__L3_N41;
   input clk_m__L3_N42;
   input clk_m__L3_N43;
   input clk_m__L3_N44;
   input clk_m__L3_N45;
   input clk_m__L3_N46;
   input clk_m__L3_N47;
   input clk_m__L3_N48;
   input clk_m__L3_N49;
   input clk_m__L3_N5;
   input clk_m__L3_N50;
   input clk_m__L3_N52;
   input clk_m__L3_N53;
   input clk_m__L3_N54;
   input clk_m__L3_N55;
   input clk_m__L3_N56;
   input clk_m__L3_N57;
   input clk_m__L3_N58;
   input clk_m__L3_N59;
   input clk_m__L3_N6;
   input clk_m__L3_N60;
   input clk_m__L3_N61;
   input clk_m__L3_N62;
   input clk_m__L3_N63;
   input clk_m__L3_N64;
   input clk_m__L3_N65;
   input clk_m__L3_N66;
   input clk_m__L3_N67;
   input clk_m__L3_N68;
   input clk_m__L3_N69;
   input clk_m__L3_N7;
   input clk_m__L3_N70;
   input clk_m__L3_N71;
   input clk_m__L3_N72;
   input clk_m__L3_N73;
   input clk_m__L3_N74;
   input clk_m__L3_N75;
   input clk_m__L3_N76;
   input clk_m__L3_N77;
   input clk_m__L3_N78;
   input clk_m__L3_N79;
   input clk_m__L3_N8;
   input clk_m__L3_N80;
   input clk_m__L3_N81;
   input clk_m__L3_N82;
   input clk_m__L3_N83;
   input clk_m__L3_N84;
   input clk_m__L3_N85;
   input clk_m__L3_N86;
   input clk_m__L3_N87;
   input clk_m__L3_N88;
   input clk_m__L3_N89;
   input clk_m__L3_N9;
   input clk_m__L3_N90;
   input clk_m__L3_N91;
   input clk_m__L3_N92;
   input clk_m__L3_N93;
   input clk_m__L3_N94;
   input clk_m__L3_N95;
   input clk_m__L3_N96;
   input clk_m__L3_N97;
   input clk_m__L3_N98;
   input clk_m__L3_N99;
   input clk_m__N0;

   // Internal wires
   wire FE_OFN94_mem_write;
   wire FE_OFN93_mem_write;
   wire FE_OFN92_mem_write;
   wire FE_OFN91_n23;
   wire FE_OFN90_n23;
   wire FE_OFN89_n23;
   wire FE_OFN88_n22;
   wire FE_OFN87_n22;
   wire FE_OFN86_n22;
   wire FE_OFN85_n21;
   wire FE_OFN84_n21;
   wire FE_OFN83_n21;
   wire FE_OFN82_n20;
   wire FE_OFN81_n20;
   wire FE_OFN80_n20;
   wire FE_OFN79_n20;
   wire FE_OFN78_n19;
   wire FE_OFN77_n19;
   wire FE_OFN76_n19;
   wire FE_OFN75_n18;
   wire FE_OFN74_n18;
   wire FE_OFN73_n18;
   wire FE_OFN72_n17;
   wire FE_OFN71_n17;
   wire FE_OFN70_n17;
   wire FE_OFN69_n16;
   wire FE_OFN68_n16;
   wire FE_OFN67_n16;
   wire FE_OFN66_n16;
   wire FE_OFN65_n15;
   wire FE_OFN64_n15;
   wire FE_OFN63_n15;
   wire FE_OFN62_n14;
   wire FE_OFN61_n14;
   wire FE_OFN60_n14;
   wire FE_OFN59_n14;
   wire FE_OFN58_n13;
   wire FE_OFN57_n13;
   wire FE_OFN56_n13;
   wire FE_OFN55_n12;
   wire FE_OFN54_n12;
   wire FE_OFN53_n12;
   wire FE_OFN52_n11;
   wire FE_OFN51_n11;
   wire FE_OFN50_n11;
   wire FE_OFN49_n10;
   wire FE_OFN48_n10;
   wire FE_OFN47_n10;
   wire FE_OFN46_n9;
   wire FE_OFN45_n9;
   wire FE_OFN44_n9;
   wire FE_OFN43_n6;
   wire FE_OFN42_n6;
   wire FE_OFN41_n6;
   wire FE_OFN40_n6459;
   wire FE_OFN39_n6459;
   wire FE_OFN38_n6459;
   wire FE_OFN37_n6459;
   wire FE_OFN36_n6459;
   wire FE_OFN35_n6459;
   wire FE_OFN34_n6459;
   wire FE_OFN33_n6459;
   wire FE_OFN32_n6459;
   wire FE_OFN31_n6459;
   wire FE_OFN30_n6459;
   wire FE_OFN29_n6459;
   wire FE_OFN28_n6459;
   wire FE_OFN27_n6459;
   wire FE_OFN26_n6459;
   wire FE_OFN25_n6459;
   wire FE_OFN24_n6136;
   wire FE_OFN23_n6136;
   wire FE_OFN22_n6136;
   wire FE_OFN21_n7440;
   wire FE_OFN20_n7440;
   wire FE_OFN19_n7440;
   wire FE_OFN18_n7440;
   wire FE_OFN17_n7440;
   wire FE_OFN16_n7440;
   wire FE_OFN15_n7440;
   wire FE_OFN14_n7440;
   wire FE_OFN13_n7440;
   wire FE_OFN12_n7440;
   wire FE_OFN11_n7440;
   wire FE_OFN10_n7440;
   wire FE_OFN9_n7440;
   wire FE_OFN8_n7440;
   wire FE_OFN7_n7440;
   wire FE_OFN6_n7440;
   wire FE_OFN5_n7440;
   wire FE_OFN4_n7442;
   wire FE_OFN3_n7442;
   wire FE_OFN2_n7442;
   wire FE_OFN1_n7442;
   wire FE_OFN0_n7442;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire \ram[255][15] ;
   wire \ram[255][14] ;
   wire \ram[255][13] ;
   wire \ram[255][12] ;
   wire \ram[255][11] ;
   wire \ram[255][10] ;
   wire \ram[255][9] ;
   wire \ram[255][8] ;
   wire \ram[255][7] ;
   wire \ram[255][6] ;
   wire \ram[255][5] ;
   wire \ram[255][4] ;
   wire \ram[255][3] ;
   wire \ram[255][2] ;
   wire \ram[255][1] ;
   wire \ram[255][0] ;
   wire \ram[254][15] ;
   wire \ram[254][14] ;
   wire \ram[254][13] ;
   wire \ram[254][12] ;
   wire \ram[254][11] ;
   wire \ram[254][10] ;
   wire \ram[254][9] ;
   wire \ram[254][8] ;
   wire \ram[254][7] ;
   wire \ram[254][6] ;
   wire \ram[254][5] ;
   wire \ram[254][4] ;
   wire \ram[254][3] ;
   wire \ram[254][2] ;
   wire \ram[254][1] ;
   wire \ram[254][0] ;
   wire \ram[253][15] ;
   wire \ram[253][14] ;
   wire \ram[253][13] ;
   wire \ram[253][12] ;
   wire \ram[253][11] ;
   wire \ram[253][10] ;
   wire \ram[253][9] ;
   wire \ram[253][8] ;
   wire \ram[253][7] ;
   wire \ram[253][6] ;
   wire \ram[253][5] ;
   wire \ram[253][4] ;
   wire \ram[253][3] ;
   wire \ram[253][2] ;
   wire \ram[253][1] ;
   wire \ram[253][0] ;
   wire \ram[252][15] ;
   wire \ram[252][14] ;
   wire \ram[252][13] ;
   wire \ram[252][12] ;
   wire \ram[252][11] ;
   wire \ram[252][10] ;
   wire \ram[252][9] ;
   wire \ram[252][8] ;
   wire \ram[252][7] ;
   wire \ram[252][6] ;
   wire \ram[252][5] ;
   wire \ram[252][4] ;
   wire \ram[252][3] ;
   wire \ram[252][2] ;
   wire \ram[252][1] ;
   wire \ram[252][0] ;
   wire \ram[251][15] ;
   wire \ram[251][14] ;
   wire \ram[251][13] ;
   wire \ram[251][12] ;
   wire \ram[251][11] ;
   wire \ram[251][10] ;
   wire \ram[251][9] ;
   wire \ram[251][8] ;
   wire \ram[251][7] ;
   wire \ram[251][6] ;
   wire \ram[251][5] ;
   wire \ram[251][4] ;
   wire \ram[251][3] ;
   wire \ram[251][2] ;
   wire \ram[251][1] ;
   wire \ram[251][0] ;
   wire \ram[250][15] ;
   wire \ram[250][14] ;
   wire \ram[250][13] ;
   wire \ram[250][12] ;
   wire \ram[250][11] ;
   wire \ram[250][10] ;
   wire \ram[250][9] ;
   wire \ram[250][8] ;
   wire \ram[250][7] ;
   wire \ram[250][6] ;
   wire \ram[250][5] ;
   wire \ram[250][4] ;
   wire \ram[250][3] ;
   wire \ram[250][2] ;
   wire \ram[250][1] ;
   wire \ram[250][0] ;
   wire \ram[249][15] ;
   wire \ram[249][14] ;
   wire \ram[249][13] ;
   wire \ram[249][12] ;
   wire \ram[249][11] ;
   wire \ram[249][10] ;
   wire \ram[249][9] ;
   wire \ram[249][8] ;
   wire \ram[249][7] ;
   wire \ram[249][6] ;
   wire \ram[249][5] ;
   wire \ram[249][4] ;
   wire \ram[249][3] ;
   wire \ram[249][2] ;
   wire \ram[249][1] ;
   wire \ram[249][0] ;
   wire \ram[248][15] ;
   wire \ram[248][14] ;
   wire \ram[248][13] ;
   wire \ram[248][12] ;
   wire \ram[248][11] ;
   wire \ram[248][10] ;
   wire \ram[248][9] ;
   wire \ram[248][8] ;
   wire \ram[248][7] ;
   wire \ram[248][6] ;
   wire \ram[248][5] ;
   wire \ram[248][4] ;
   wire \ram[248][3] ;
   wire \ram[248][2] ;
   wire \ram[248][1] ;
   wire \ram[248][0] ;
   wire \ram[247][15] ;
   wire \ram[247][14] ;
   wire \ram[247][13] ;
   wire \ram[247][12] ;
   wire \ram[247][11] ;
   wire \ram[247][10] ;
   wire \ram[247][9] ;
   wire \ram[247][8] ;
   wire \ram[247][7] ;
   wire \ram[247][6] ;
   wire \ram[247][5] ;
   wire \ram[247][4] ;
   wire \ram[247][3] ;
   wire \ram[247][2] ;
   wire \ram[247][1] ;
   wire \ram[247][0] ;
   wire \ram[246][15] ;
   wire \ram[246][14] ;
   wire \ram[246][13] ;
   wire \ram[246][12] ;
   wire \ram[246][11] ;
   wire \ram[246][10] ;
   wire \ram[246][9] ;
   wire \ram[246][8] ;
   wire \ram[246][7] ;
   wire \ram[246][6] ;
   wire \ram[246][5] ;
   wire \ram[246][4] ;
   wire \ram[246][3] ;
   wire \ram[246][2] ;
   wire \ram[246][1] ;
   wire \ram[246][0] ;
   wire \ram[245][15] ;
   wire \ram[245][14] ;
   wire \ram[245][13] ;
   wire \ram[245][12] ;
   wire \ram[245][11] ;
   wire \ram[245][10] ;
   wire \ram[245][9] ;
   wire \ram[245][8] ;
   wire \ram[245][7] ;
   wire \ram[245][6] ;
   wire \ram[245][5] ;
   wire \ram[245][4] ;
   wire \ram[245][3] ;
   wire \ram[245][2] ;
   wire \ram[245][1] ;
   wire \ram[245][0] ;
   wire \ram[244][15] ;
   wire \ram[244][14] ;
   wire \ram[244][13] ;
   wire \ram[244][12] ;
   wire \ram[244][11] ;
   wire \ram[244][10] ;
   wire \ram[244][9] ;
   wire \ram[244][8] ;
   wire \ram[244][7] ;
   wire \ram[244][6] ;
   wire \ram[244][5] ;
   wire \ram[244][4] ;
   wire \ram[244][3] ;
   wire \ram[244][2] ;
   wire \ram[244][1] ;
   wire \ram[244][0] ;
   wire \ram[243][15] ;
   wire \ram[243][14] ;
   wire \ram[243][13] ;
   wire \ram[243][12] ;
   wire \ram[243][11] ;
   wire \ram[243][10] ;
   wire \ram[243][9] ;
   wire \ram[243][8] ;
   wire \ram[243][7] ;
   wire \ram[243][6] ;
   wire \ram[243][5] ;
   wire \ram[243][4] ;
   wire \ram[243][3] ;
   wire \ram[243][2] ;
   wire \ram[243][1] ;
   wire \ram[243][0] ;
   wire \ram[242][15] ;
   wire \ram[242][14] ;
   wire \ram[242][13] ;
   wire \ram[242][12] ;
   wire \ram[242][11] ;
   wire \ram[242][10] ;
   wire \ram[242][9] ;
   wire \ram[242][8] ;
   wire \ram[242][7] ;
   wire \ram[242][6] ;
   wire \ram[242][5] ;
   wire \ram[242][4] ;
   wire \ram[242][3] ;
   wire \ram[242][2] ;
   wire \ram[242][1] ;
   wire \ram[242][0] ;
   wire \ram[241][15] ;
   wire \ram[241][14] ;
   wire \ram[241][13] ;
   wire \ram[241][12] ;
   wire \ram[241][11] ;
   wire \ram[241][10] ;
   wire \ram[241][9] ;
   wire \ram[241][8] ;
   wire \ram[241][7] ;
   wire \ram[241][6] ;
   wire \ram[241][5] ;
   wire \ram[241][4] ;
   wire \ram[241][3] ;
   wire \ram[241][2] ;
   wire \ram[241][1] ;
   wire \ram[241][0] ;
   wire \ram[240][15] ;
   wire \ram[240][14] ;
   wire \ram[240][13] ;
   wire \ram[240][12] ;
   wire \ram[240][11] ;
   wire \ram[240][10] ;
   wire \ram[240][9] ;
   wire \ram[240][8] ;
   wire \ram[240][7] ;
   wire \ram[240][6] ;
   wire \ram[240][5] ;
   wire \ram[240][4] ;
   wire \ram[240][3] ;
   wire \ram[240][2] ;
   wire \ram[240][1] ;
   wire \ram[240][0] ;
   wire \ram[239][15] ;
   wire \ram[239][14] ;
   wire \ram[239][13] ;
   wire \ram[239][12] ;
   wire \ram[239][11] ;
   wire \ram[239][10] ;
   wire \ram[239][9] ;
   wire \ram[239][8] ;
   wire \ram[239][7] ;
   wire \ram[239][6] ;
   wire \ram[239][5] ;
   wire \ram[239][4] ;
   wire \ram[239][3] ;
   wire \ram[239][2] ;
   wire \ram[239][1] ;
   wire \ram[239][0] ;
   wire \ram[238][15] ;
   wire \ram[238][14] ;
   wire \ram[238][13] ;
   wire \ram[238][12] ;
   wire \ram[238][11] ;
   wire \ram[238][10] ;
   wire \ram[238][9] ;
   wire \ram[238][8] ;
   wire \ram[238][7] ;
   wire \ram[238][6] ;
   wire \ram[238][5] ;
   wire \ram[238][4] ;
   wire \ram[238][3] ;
   wire \ram[238][2] ;
   wire \ram[238][1] ;
   wire \ram[238][0] ;
   wire \ram[237][15] ;
   wire \ram[237][14] ;
   wire \ram[237][13] ;
   wire \ram[237][12] ;
   wire \ram[237][11] ;
   wire \ram[237][10] ;
   wire \ram[237][9] ;
   wire \ram[237][8] ;
   wire \ram[237][7] ;
   wire \ram[237][6] ;
   wire \ram[237][5] ;
   wire \ram[237][4] ;
   wire \ram[237][3] ;
   wire \ram[237][2] ;
   wire \ram[237][1] ;
   wire \ram[237][0] ;
   wire \ram[236][15] ;
   wire \ram[236][14] ;
   wire \ram[236][13] ;
   wire \ram[236][12] ;
   wire \ram[236][11] ;
   wire \ram[236][10] ;
   wire \ram[236][9] ;
   wire \ram[236][8] ;
   wire \ram[236][7] ;
   wire \ram[236][6] ;
   wire \ram[236][5] ;
   wire \ram[236][4] ;
   wire \ram[236][3] ;
   wire \ram[236][2] ;
   wire \ram[236][1] ;
   wire \ram[236][0] ;
   wire \ram[235][15] ;
   wire \ram[235][14] ;
   wire \ram[235][13] ;
   wire \ram[235][12] ;
   wire \ram[235][11] ;
   wire \ram[235][10] ;
   wire \ram[235][9] ;
   wire \ram[235][8] ;
   wire \ram[235][7] ;
   wire \ram[235][6] ;
   wire \ram[235][5] ;
   wire \ram[235][4] ;
   wire \ram[235][3] ;
   wire \ram[235][2] ;
   wire \ram[235][1] ;
   wire \ram[235][0] ;
   wire \ram[234][15] ;
   wire \ram[234][14] ;
   wire \ram[234][13] ;
   wire \ram[234][12] ;
   wire \ram[234][11] ;
   wire \ram[234][10] ;
   wire \ram[234][9] ;
   wire \ram[234][8] ;
   wire \ram[234][7] ;
   wire \ram[234][6] ;
   wire \ram[234][5] ;
   wire \ram[234][4] ;
   wire \ram[234][3] ;
   wire \ram[234][2] ;
   wire \ram[234][1] ;
   wire \ram[234][0] ;
   wire \ram[233][15] ;
   wire \ram[233][14] ;
   wire \ram[233][13] ;
   wire \ram[233][12] ;
   wire \ram[233][11] ;
   wire \ram[233][10] ;
   wire \ram[233][9] ;
   wire \ram[233][8] ;
   wire \ram[233][7] ;
   wire \ram[233][6] ;
   wire \ram[233][5] ;
   wire \ram[233][4] ;
   wire \ram[233][3] ;
   wire \ram[233][2] ;
   wire \ram[233][1] ;
   wire \ram[233][0] ;
   wire \ram[232][15] ;
   wire \ram[232][14] ;
   wire \ram[232][13] ;
   wire \ram[232][12] ;
   wire \ram[232][11] ;
   wire \ram[232][10] ;
   wire \ram[232][9] ;
   wire \ram[232][8] ;
   wire \ram[232][7] ;
   wire \ram[232][6] ;
   wire \ram[232][5] ;
   wire \ram[232][4] ;
   wire \ram[232][3] ;
   wire \ram[232][2] ;
   wire \ram[232][1] ;
   wire \ram[232][0] ;
   wire \ram[231][15] ;
   wire \ram[231][14] ;
   wire \ram[231][13] ;
   wire \ram[231][12] ;
   wire \ram[231][11] ;
   wire \ram[231][10] ;
   wire \ram[231][9] ;
   wire \ram[231][8] ;
   wire \ram[231][7] ;
   wire \ram[231][6] ;
   wire \ram[231][5] ;
   wire \ram[231][4] ;
   wire \ram[231][3] ;
   wire \ram[231][2] ;
   wire \ram[231][1] ;
   wire \ram[231][0] ;
   wire \ram[230][15] ;
   wire \ram[230][14] ;
   wire \ram[230][13] ;
   wire \ram[230][12] ;
   wire \ram[230][11] ;
   wire \ram[230][10] ;
   wire \ram[230][9] ;
   wire \ram[230][8] ;
   wire \ram[230][7] ;
   wire \ram[230][6] ;
   wire \ram[230][5] ;
   wire \ram[230][4] ;
   wire \ram[230][3] ;
   wire \ram[230][2] ;
   wire \ram[230][1] ;
   wire \ram[230][0] ;
   wire \ram[229][15] ;
   wire \ram[229][14] ;
   wire \ram[229][13] ;
   wire \ram[229][12] ;
   wire \ram[229][11] ;
   wire \ram[229][10] ;
   wire \ram[229][9] ;
   wire \ram[229][8] ;
   wire \ram[229][7] ;
   wire \ram[229][6] ;
   wire \ram[229][5] ;
   wire \ram[229][4] ;
   wire \ram[229][3] ;
   wire \ram[229][2] ;
   wire \ram[229][1] ;
   wire \ram[229][0] ;
   wire \ram[228][15] ;
   wire \ram[228][14] ;
   wire \ram[228][13] ;
   wire \ram[228][12] ;
   wire \ram[228][11] ;
   wire \ram[228][10] ;
   wire \ram[228][9] ;
   wire \ram[228][8] ;
   wire \ram[228][7] ;
   wire \ram[228][6] ;
   wire \ram[228][5] ;
   wire \ram[228][4] ;
   wire \ram[228][3] ;
   wire \ram[228][2] ;
   wire \ram[228][1] ;
   wire \ram[228][0] ;
   wire \ram[227][15] ;
   wire \ram[227][14] ;
   wire \ram[227][13] ;
   wire \ram[227][12] ;
   wire \ram[227][11] ;
   wire \ram[227][10] ;
   wire \ram[227][9] ;
   wire \ram[227][8] ;
   wire \ram[227][7] ;
   wire \ram[227][6] ;
   wire \ram[227][5] ;
   wire \ram[227][4] ;
   wire \ram[227][3] ;
   wire \ram[227][2] ;
   wire \ram[227][1] ;
   wire \ram[227][0] ;
   wire \ram[226][15] ;
   wire \ram[226][14] ;
   wire \ram[226][13] ;
   wire \ram[226][12] ;
   wire \ram[226][11] ;
   wire \ram[226][10] ;
   wire \ram[226][9] ;
   wire \ram[226][8] ;
   wire \ram[226][7] ;
   wire \ram[226][6] ;
   wire \ram[226][5] ;
   wire \ram[226][4] ;
   wire \ram[226][3] ;
   wire \ram[226][2] ;
   wire \ram[226][1] ;
   wire \ram[226][0] ;
   wire \ram[225][15] ;
   wire \ram[225][14] ;
   wire \ram[225][13] ;
   wire \ram[225][12] ;
   wire \ram[225][11] ;
   wire \ram[225][10] ;
   wire \ram[225][9] ;
   wire \ram[225][8] ;
   wire \ram[225][7] ;
   wire \ram[225][6] ;
   wire \ram[225][5] ;
   wire \ram[225][4] ;
   wire \ram[225][3] ;
   wire \ram[225][2] ;
   wire \ram[225][1] ;
   wire \ram[225][0] ;
   wire \ram[224][15] ;
   wire \ram[224][14] ;
   wire \ram[224][13] ;
   wire \ram[224][12] ;
   wire \ram[224][11] ;
   wire \ram[224][10] ;
   wire \ram[224][9] ;
   wire \ram[224][8] ;
   wire \ram[224][7] ;
   wire \ram[224][6] ;
   wire \ram[224][5] ;
   wire \ram[224][4] ;
   wire \ram[224][3] ;
   wire \ram[224][2] ;
   wire \ram[224][1] ;
   wire \ram[224][0] ;
   wire \ram[223][15] ;
   wire \ram[223][14] ;
   wire \ram[223][13] ;
   wire \ram[223][12] ;
   wire \ram[223][11] ;
   wire \ram[223][10] ;
   wire \ram[223][9] ;
   wire \ram[223][8] ;
   wire \ram[223][7] ;
   wire \ram[223][6] ;
   wire \ram[223][5] ;
   wire \ram[223][4] ;
   wire \ram[223][3] ;
   wire \ram[223][2] ;
   wire \ram[223][1] ;
   wire \ram[223][0] ;
   wire \ram[222][15] ;
   wire \ram[222][14] ;
   wire \ram[222][13] ;
   wire \ram[222][12] ;
   wire \ram[222][11] ;
   wire \ram[222][10] ;
   wire \ram[222][9] ;
   wire \ram[222][8] ;
   wire \ram[222][7] ;
   wire \ram[222][6] ;
   wire \ram[222][5] ;
   wire \ram[222][4] ;
   wire \ram[222][3] ;
   wire \ram[222][2] ;
   wire \ram[222][1] ;
   wire \ram[222][0] ;
   wire \ram[221][15] ;
   wire \ram[221][14] ;
   wire \ram[221][13] ;
   wire \ram[221][12] ;
   wire \ram[221][11] ;
   wire \ram[221][10] ;
   wire \ram[221][9] ;
   wire \ram[221][8] ;
   wire \ram[221][7] ;
   wire \ram[221][6] ;
   wire \ram[221][5] ;
   wire \ram[221][4] ;
   wire \ram[221][3] ;
   wire \ram[221][2] ;
   wire \ram[221][1] ;
   wire \ram[221][0] ;
   wire \ram[220][15] ;
   wire \ram[220][14] ;
   wire \ram[220][13] ;
   wire \ram[220][12] ;
   wire \ram[220][11] ;
   wire \ram[220][10] ;
   wire \ram[220][9] ;
   wire \ram[220][8] ;
   wire \ram[220][7] ;
   wire \ram[220][6] ;
   wire \ram[220][5] ;
   wire \ram[220][4] ;
   wire \ram[220][3] ;
   wire \ram[220][2] ;
   wire \ram[220][1] ;
   wire \ram[220][0] ;
   wire \ram[219][15] ;
   wire \ram[219][14] ;
   wire \ram[219][13] ;
   wire \ram[219][12] ;
   wire \ram[219][11] ;
   wire \ram[219][10] ;
   wire \ram[219][9] ;
   wire \ram[219][8] ;
   wire \ram[219][7] ;
   wire \ram[219][6] ;
   wire \ram[219][5] ;
   wire \ram[219][4] ;
   wire \ram[219][3] ;
   wire \ram[219][2] ;
   wire \ram[219][1] ;
   wire \ram[219][0] ;
   wire \ram[218][15] ;
   wire \ram[218][14] ;
   wire \ram[218][13] ;
   wire \ram[218][12] ;
   wire \ram[218][11] ;
   wire \ram[218][10] ;
   wire \ram[218][9] ;
   wire \ram[218][8] ;
   wire \ram[218][7] ;
   wire \ram[218][6] ;
   wire \ram[218][5] ;
   wire \ram[218][4] ;
   wire \ram[218][3] ;
   wire \ram[218][2] ;
   wire \ram[218][1] ;
   wire \ram[218][0] ;
   wire \ram[217][15] ;
   wire \ram[217][14] ;
   wire \ram[217][13] ;
   wire \ram[217][12] ;
   wire \ram[217][11] ;
   wire \ram[217][10] ;
   wire \ram[217][9] ;
   wire \ram[217][8] ;
   wire \ram[217][7] ;
   wire \ram[217][6] ;
   wire \ram[217][5] ;
   wire \ram[217][4] ;
   wire \ram[217][3] ;
   wire \ram[217][2] ;
   wire \ram[217][1] ;
   wire \ram[217][0] ;
   wire \ram[216][15] ;
   wire \ram[216][14] ;
   wire \ram[216][13] ;
   wire \ram[216][12] ;
   wire \ram[216][11] ;
   wire \ram[216][10] ;
   wire \ram[216][9] ;
   wire \ram[216][8] ;
   wire \ram[216][7] ;
   wire \ram[216][6] ;
   wire \ram[216][5] ;
   wire \ram[216][4] ;
   wire \ram[216][3] ;
   wire \ram[216][2] ;
   wire \ram[216][1] ;
   wire \ram[216][0] ;
   wire \ram[215][15] ;
   wire \ram[215][14] ;
   wire \ram[215][13] ;
   wire \ram[215][12] ;
   wire \ram[215][11] ;
   wire \ram[215][10] ;
   wire \ram[215][9] ;
   wire \ram[215][8] ;
   wire \ram[215][7] ;
   wire \ram[215][6] ;
   wire \ram[215][5] ;
   wire \ram[215][4] ;
   wire \ram[215][3] ;
   wire \ram[215][2] ;
   wire \ram[215][1] ;
   wire \ram[215][0] ;
   wire \ram[214][15] ;
   wire \ram[214][14] ;
   wire \ram[214][13] ;
   wire \ram[214][12] ;
   wire \ram[214][11] ;
   wire \ram[214][10] ;
   wire \ram[214][9] ;
   wire \ram[214][8] ;
   wire \ram[214][7] ;
   wire \ram[214][6] ;
   wire \ram[214][5] ;
   wire \ram[214][4] ;
   wire \ram[214][3] ;
   wire \ram[214][2] ;
   wire \ram[214][1] ;
   wire \ram[214][0] ;
   wire \ram[213][15] ;
   wire \ram[213][14] ;
   wire \ram[213][13] ;
   wire \ram[213][12] ;
   wire \ram[213][11] ;
   wire \ram[213][10] ;
   wire \ram[213][9] ;
   wire \ram[213][8] ;
   wire \ram[213][7] ;
   wire \ram[213][6] ;
   wire \ram[213][5] ;
   wire \ram[213][4] ;
   wire \ram[213][3] ;
   wire \ram[213][2] ;
   wire \ram[213][1] ;
   wire \ram[213][0] ;
   wire \ram[212][15] ;
   wire \ram[212][14] ;
   wire \ram[212][13] ;
   wire \ram[212][12] ;
   wire \ram[212][11] ;
   wire \ram[212][10] ;
   wire \ram[212][9] ;
   wire \ram[212][8] ;
   wire \ram[212][7] ;
   wire \ram[212][6] ;
   wire \ram[212][5] ;
   wire \ram[212][4] ;
   wire \ram[212][3] ;
   wire \ram[212][2] ;
   wire \ram[212][1] ;
   wire \ram[212][0] ;
   wire \ram[211][15] ;
   wire \ram[211][14] ;
   wire \ram[211][13] ;
   wire \ram[211][12] ;
   wire \ram[211][11] ;
   wire \ram[211][10] ;
   wire \ram[211][9] ;
   wire \ram[211][8] ;
   wire \ram[211][7] ;
   wire \ram[211][6] ;
   wire \ram[211][5] ;
   wire \ram[211][4] ;
   wire \ram[211][3] ;
   wire \ram[211][2] ;
   wire \ram[211][1] ;
   wire \ram[211][0] ;
   wire \ram[210][15] ;
   wire \ram[210][14] ;
   wire \ram[210][13] ;
   wire \ram[210][12] ;
   wire \ram[210][11] ;
   wire \ram[210][10] ;
   wire \ram[210][9] ;
   wire \ram[210][8] ;
   wire \ram[210][7] ;
   wire \ram[210][6] ;
   wire \ram[210][5] ;
   wire \ram[210][4] ;
   wire \ram[210][3] ;
   wire \ram[210][2] ;
   wire \ram[210][1] ;
   wire \ram[210][0] ;
   wire \ram[209][15] ;
   wire \ram[209][14] ;
   wire \ram[209][13] ;
   wire \ram[209][12] ;
   wire \ram[209][11] ;
   wire \ram[209][10] ;
   wire \ram[209][9] ;
   wire \ram[209][8] ;
   wire \ram[209][7] ;
   wire \ram[209][6] ;
   wire \ram[209][5] ;
   wire \ram[209][4] ;
   wire \ram[209][3] ;
   wire \ram[209][2] ;
   wire \ram[209][1] ;
   wire \ram[209][0] ;
   wire \ram[208][15] ;
   wire \ram[208][14] ;
   wire \ram[208][13] ;
   wire \ram[208][12] ;
   wire \ram[208][11] ;
   wire \ram[208][10] ;
   wire \ram[208][9] ;
   wire \ram[208][8] ;
   wire \ram[208][7] ;
   wire \ram[208][6] ;
   wire \ram[208][5] ;
   wire \ram[208][4] ;
   wire \ram[208][3] ;
   wire \ram[208][2] ;
   wire \ram[208][1] ;
   wire \ram[208][0] ;
   wire \ram[207][15] ;
   wire \ram[207][14] ;
   wire \ram[207][13] ;
   wire \ram[207][12] ;
   wire \ram[207][11] ;
   wire \ram[207][10] ;
   wire \ram[207][9] ;
   wire \ram[207][8] ;
   wire \ram[207][7] ;
   wire \ram[207][6] ;
   wire \ram[207][5] ;
   wire \ram[207][4] ;
   wire \ram[207][3] ;
   wire \ram[207][2] ;
   wire \ram[207][1] ;
   wire \ram[207][0] ;
   wire \ram[206][15] ;
   wire \ram[206][14] ;
   wire \ram[206][13] ;
   wire \ram[206][12] ;
   wire \ram[206][11] ;
   wire \ram[206][10] ;
   wire \ram[206][9] ;
   wire \ram[206][8] ;
   wire \ram[206][7] ;
   wire \ram[206][6] ;
   wire \ram[206][5] ;
   wire \ram[206][4] ;
   wire \ram[206][3] ;
   wire \ram[206][2] ;
   wire \ram[206][1] ;
   wire \ram[206][0] ;
   wire \ram[205][15] ;
   wire \ram[205][14] ;
   wire \ram[205][13] ;
   wire \ram[205][12] ;
   wire \ram[205][11] ;
   wire \ram[205][10] ;
   wire \ram[205][9] ;
   wire \ram[205][8] ;
   wire \ram[205][7] ;
   wire \ram[205][6] ;
   wire \ram[205][5] ;
   wire \ram[205][4] ;
   wire \ram[205][3] ;
   wire \ram[205][2] ;
   wire \ram[205][1] ;
   wire \ram[205][0] ;
   wire \ram[204][15] ;
   wire \ram[204][14] ;
   wire \ram[204][13] ;
   wire \ram[204][12] ;
   wire \ram[204][11] ;
   wire \ram[204][10] ;
   wire \ram[204][9] ;
   wire \ram[204][8] ;
   wire \ram[204][7] ;
   wire \ram[204][6] ;
   wire \ram[204][5] ;
   wire \ram[204][4] ;
   wire \ram[204][3] ;
   wire \ram[204][2] ;
   wire \ram[204][1] ;
   wire \ram[204][0] ;
   wire \ram[203][15] ;
   wire \ram[203][14] ;
   wire \ram[203][13] ;
   wire \ram[203][12] ;
   wire \ram[203][11] ;
   wire \ram[203][10] ;
   wire \ram[203][9] ;
   wire \ram[203][8] ;
   wire \ram[203][7] ;
   wire \ram[203][6] ;
   wire \ram[203][5] ;
   wire \ram[203][4] ;
   wire \ram[203][3] ;
   wire \ram[203][2] ;
   wire \ram[203][1] ;
   wire \ram[203][0] ;
   wire \ram[202][15] ;
   wire \ram[202][14] ;
   wire \ram[202][13] ;
   wire \ram[202][12] ;
   wire \ram[202][11] ;
   wire \ram[202][10] ;
   wire \ram[202][9] ;
   wire \ram[202][8] ;
   wire \ram[202][7] ;
   wire \ram[202][6] ;
   wire \ram[202][5] ;
   wire \ram[202][4] ;
   wire \ram[202][3] ;
   wire \ram[202][2] ;
   wire \ram[202][1] ;
   wire \ram[202][0] ;
   wire \ram[201][15] ;
   wire \ram[201][14] ;
   wire \ram[201][13] ;
   wire \ram[201][12] ;
   wire \ram[201][11] ;
   wire \ram[201][10] ;
   wire \ram[201][9] ;
   wire \ram[201][8] ;
   wire \ram[201][7] ;
   wire \ram[201][6] ;
   wire \ram[201][5] ;
   wire \ram[201][4] ;
   wire \ram[201][3] ;
   wire \ram[201][2] ;
   wire \ram[201][1] ;
   wire \ram[201][0] ;
   wire \ram[200][15] ;
   wire \ram[200][14] ;
   wire \ram[200][13] ;
   wire \ram[200][12] ;
   wire \ram[200][11] ;
   wire \ram[200][10] ;
   wire \ram[200][9] ;
   wire \ram[200][8] ;
   wire \ram[200][7] ;
   wire \ram[200][6] ;
   wire \ram[200][5] ;
   wire \ram[200][4] ;
   wire \ram[200][3] ;
   wire \ram[200][2] ;
   wire \ram[200][1] ;
   wire \ram[200][0] ;
   wire \ram[199][15] ;
   wire \ram[199][14] ;
   wire \ram[199][13] ;
   wire \ram[199][12] ;
   wire \ram[199][11] ;
   wire \ram[199][10] ;
   wire \ram[199][9] ;
   wire \ram[199][8] ;
   wire \ram[199][7] ;
   wire \ram[199][6] ;
   wire \ram[199][5] ;
   wire \ram[199][4] ;
   wire \ram[199][3] ;
   wire \ram[199][2] ;
   wire \ram[199][1] ;
   wire \ram[199][0] ;
   wire \ram[198][15] ;
   wire \ram[198][14] ;
   wire \ram[198][13] ;
   wire \ram[198][12] ;
   wire \ram[198][11] ;
   wire \ram[198][10] ;
   wire \ram[198][9] ;
   wire \ram[198][8] ;
   wire \ram[198][7] ;
   wire \ram[198][6] ;
   wire \ram[198][5] ;
   wire \ram[198][4] ;
   wire \ram[198][3] ;
   wire \ram[198][2] ;
   wire \ram[198][1] ;
   wire \ram[198][0] ;
   wire \ram[197][15] ;
   wire \ram[197][14] ;
   wire \ram[197][13] ;
   wire \ram[197][12] ;
   wire \ram[197][11] ;
   wire \ram[197][10] ;
   wire \ram[197][9] ;
   wire \ram[197][8] ;
   wire \ram[197][7] ;
   wire \ram[197][6] ;
   wire \ram[197][5] ;
   wire \ram[197][4] ;
   wire \ram[197][3] ;
   wire \ram[197][2] ;
   wire \ram[197][1] ;
   wire \ram[197][0] ;
   wire \ram[196][15] ;
   wire \ram[196][14] ;
   wire \ram[196][13] ;
   wire \ram[196][12] ;
   wire \ram[196][11] ;
   wire \ram[196][10] ;
   wire \ram[196][9] ;
   wire \ram[196][8] ;
   wire \ram[196][7] ;
   wire \ram[196][6] ;
   wire \ram[196][5] ;
   wire \ram[196][4] ;
   wire \ram[196][3] ;
   wire \ram[196][2] ;
   wire \ram[196][1] ;
   wire \ram[196][0] ;
   wire \ram[195][15] ;
   wire \ram[195][14] ;
   wire \ram[195][13] ;
   wire \ram[195][12] ;
   wire \ram[195][11] ;
   wire \ram[195][10] ;
   wire \ram[195][9] ;
   wire \ram[195][8] ;
   wire \ram[195][7] ;
   wire \ram[195][6] ;
   wire \ram[195][5] ;
   wire \ram[195][4] ;
   wire \ram[195][3] ;
   wire \ram[195][2] ;
   wire \ram[195][1] ;
   wire \ram[195][0] ;
   wire \ram[194][15] ;
   wire \ram[194][14] ;
   wire \ram[194][13] ;
   wire \ram[194][12] ;
   wire \ram[194][11] ;
   wire \ram[194][10] ;
   wire \ram[194][9] ;
   wire \ram[194][8] ;
   wire \ram[194][7] ;
   wire \ram[194][6] ;
   wire \ram[194][5] ;
   wire \ram[194][4] ;
   wire \ram[194][3] ;
   wire \ram[194][2] ;
   wire \ram[194][1] ;
   wire \ram[194][0] ;
   wire \ram[193][15] ;
   wire \ram[193][14] ;
   wire \ram[193][13] ;
   wire \ram[193][12] ;
   wire \ram[193][11] ;
   wire \ram[193][10] ;
   wire \ram[193][9] ;
   wire \ram[193][8] ;
   wire \ram[193][7] ;
   wire \ram[193][6] ;
   wire \ram[193][5] ;
   wire \ram[193][4] ;
   wire \ram[193][3] ;
   wire \ram[193][2] ;
   wire \ram[193][1] ;
   wire \ram[193][0] ;
   wire \ram[192][15] ;
   wire \ram[192][14] ;
   wire \ram[192][13] ;
   wire \ram[192][12] ;
   wire \ram[192][11] ;
   wire \ram[192][10] ;
   wire \ram[192][9] ;
   wire \ram[192][8] ;
   wire \ram[192][7] ;
   wire \ram[192][6] ;
   wire \ram[192][5] ;
   wire \ram[192][4] ;
   wire \ram[192][3] ;
   wire \ram[192][2] ;
   wire \ram[192][1] ;
   wire \ram[192][0] ;
   wire \ram[191][15] ;
   wire \ram[191][14] ;
   wire \ram[191][13] ;
   wire \ram[191][12] ;
   wire \ram[191][11] ;
   wire \ram[191][10] ;
   wire \ram[191][9] ;
   wire \ram[191][8] ;
   wire \ram[191][7] ;
   wire \ram[191][6] ;
   wire \ram[191][5] ;
   wire \ram[191][4] ;
   wire \ram[191][3] ;
   wire \ram[191][2] ;
   wire \ram[191][1] ;
   wire \ram[191][0] ;
   wire \ram[190][15] ;
   wire \ram[190][14] ;
   wire \ram[190][13] ;
   wire \ram[190][12] ;
   wire \ram[190][11] ;
   wire \ram[190][10] ;
   wire \ram[190][9] ;
   wire \ram[190][8] ;
   wire \ram[190][7] ;
   wire \ram[190][6] ;
   wire \ram[190][5] ;
   wire \ram[190][4] ;
   wire \ram[190][3] ;
   wire \ram[190][2] ;
   wire \ram[190][1] ;
   wire \ram[190][0] ;
   wire \ram[189][15] ;
   wire \ram[189][14] ;
   wire \ram[189][13] ;
   wire \ram[189][12] ;
   wire \ram[189][11] ;
   wire \ram[189][10] ;
   wire \ram[189][9] ;
   wire \ram[189][8] ;
   wire \ram[189][7] ;
   wire \ram[189][6] ;
   wire \ram[189][5] ;
   wire \ram[189][4] ;
   wire \ram[189][3] ;
   wire \ram[189][2] ;
   wire \ram[189][1] ;
   wire \ram[189][0] ;
   wire \ram[188][15] ;
   wire \ram[188][14] ;
   wire \ram[188][13] ;
   wire \ram[188][12] ;
   wire \ram[188][11] ;
   wire \ram[188][10] ;
   wire \ram[188][9] ;
   wire \ram[188][8] ;
   wire \ram[188][7] ;
   wire \ram[188][6] ;
   wire \ram[188][5] ;
   wire \ram[188][4] ;
   wire \ram[188][3] ;
   wire \ram[188][2] ;
   wire \ram[188][1] ;
   wire \ram[188][0] ;
   wire \ram[187][15] ;
   wire \ram[187][14] ;
   wire \ram[187][13] ;
   wire \ram[187][12] ;
   wire \ram[187][11] ;
   wire \ram[187][10] ;
   wire \ram[187][9] ;
   wire \ram[187][8] ;
   wire \ram[187][7] ;
   wire \ram[187][6] ;
   wire \ram[187][5] ;
   wire \ram[187][4] ;
   wire \ram[187][3] ;
   wire \ram[187][2] ;
   wire \ram[187][1] ;
   wire \ram[187][0] ;
   wire \ram[186][15] ;
   wire \ram[186][14] ;
   wire \ram[186][13] ;
   wire \ram[186][12] ;
   wire \ram[186][11] ;
   wire \ram[186][10] ;
   wire \ram[186][9] ;
   wire \ram[186][8] ;
   wire \ram[186][7] ;
   wire \ram[186][6] ;
   wire \ram[186][5] ;
   wire \ram[186][4] ;
   wire \ram[186][3] ;
   wire \ram[186][2] ;
   wire \ram[186][1] ;
   wire \ram[186][0] ;
   wire \ram[185][15] ;
   wire \ram[185][14] ;
   wire \ram[185][13] ;
   wire \ram[185][12] ;
   wire \ram[185][11] ;
   wire \ram[185][10] ;
   wire \ram[185][9] ;
   wire \ram[185][8] ;
   wire \ram[185][7] ;
   wire \ram[185][6] ;
   wire \ram[185][5] ;
   wire \ram[185][4] ;
   wire \ram[185][3] ;
   wire \ram[185][2] ;
   wire \ram[185][1] ;
   wire \ram[185][0] ;
   wire \ram[184][15] ;
   wire \ram[184][14] ;
   wire \ram[184][13] ;
   wire \ram[184][12] ;
   wire \ram[184][11] ;
   wire \ram[184][10] ;
   wire \ram[184][9] ;
   wire \ram[184][8] ;
   wire \ram[184][7] ;
   wire \ram[184][6] ;
   wire \ram[184][5] ;
   wire \ram[184][4] ;
   wire \ram[184][3] ;
   wire \ram[184][2] ;
   wire \ram[184][1] ;
   wire \ram[184][0] ;
   wire \ram[183][15] ;
   wire \ram[183][14] ;
   wire \ram[183][13] ;
   wire \ram[183][12] ;
   wire \ram[183][11] ;
   wire \ram[183][10] ;
   wire \ram[183][9] ;
   wire \ram[183][8] ;
   wire \ram[183][7] ;
   wire \ram[183][6] ;
   wire \ram[183][5] ;
   wire \ram[183][4] ;
   wire \ram[183][3] ;
   wire \ram[183][2] ;
   wire \ram[183][1] ;
   wire \ram[183][0] ;
   wire \ram[182][15] ;
   wire \ram[182][14] ;
   wire \ram[182][13] ;
   wire \ram[182][12] ;
   wire \ram[182][11] ;
   wire \ram[182][10] ;
   wire \ram[182][9] ;
   wire \ram[182][8] ;
   wire \ram[182][7] ;
   wire \ram[182][6] ;
   wire \ram[182][5] ;
   wire \ram[182][4] ;
   wire \ram[182][3] ;
   wire \ram[182][2] ;
   wire \ram[182][1] ;
   wire \ram[182][0] ;
   wire \ram[181][15] ;
   wire \ram[181][14] ;
   wire \ram[181][13] ;
   wire \ram[181][12] ;
   wire \ram[181][11] ;
   wire \ram[181][10] ;
   wire \ram[181][9] ;
   wire \ram[181][8] ;
   wire \ram[181][7] ;
   wire \ram[181][6] ;
   wire \ram[181][5] ;
   wire \ram[181][4] ;
   wire \ram[181][3] ;
   wire \ram[181][2] ;
   wire \ram[181][1] ;
   wire \ram[181][0] ;
   wire \ram[180][15] ;
   wire \ram[180][14] ;
   wire \ram[180][13] ;
   wire \ram[180][12] ;
   wire \ram[180][11] ;
   wire \ram[180][10] ;
   wire \ram[180][9] ;
   wire \ram[180][8] ;
   wire \ram[180][7] ;
   wire \ram[180][6] ;
   wire \ram[180][5] ;
   wire \ram[180][4] ;
   wire \ram[180][3] ;
   wire \ram[180][2] ;
   wire \ram[180][1] ;
   wire \ram[180][0] ;
   wire \ram[179][15] ;
   wire \ram[179][14] ;
   wire \ram[179][13] ;
   wire \ram[179][12] ;
   wire \ram[179][11] ;
   wire \ram[179][10] ;
   wire \ram[179][9] ;
   wire \ram[179][8] ;
   wire \ram[179][7] ;
   wire \ram[179][6] ;
   wire \ram[179][5] ;
   wire \ram[179][4] ;
   wire \ram[179][3] ;
   wire \ram[179][2] ;
   wire \ram[179][1] ;
   wire \ram[179][0] ;
   wire \ram[178][15] ;
   wire \ram[178][14] ;
   wire \ram[178][13] ;
   wire \ram[178][12] ;
   wire \ram[178][11] ;
   wire \ram[178][10] ;
   wire \ram[178][9] ;
   wire \ram[178][8] ;
   wire \ram[178][7] ;
   wire \ram[178][6] ;
   wire \ram[178][5] ;
   wire \ram[178][4] ;
   wire \ram[178][3] ;
   wire \ram[178][2] ;
   wire \ram[178][1] ;
   wire \ram[178][0] ;
   wire \ram[177][15] ;
   wire \ram[177][14] ;
   wire \ram[177][13] ;
   wire \ram[177][12] ;
   wire \ram[177][11] ;
   wire \ram[177][10] ;
   wire \ram[177][9] ;
   wire \ram[177][8] ;
   wire \ram[177][7] ;
   wire \ram[177][6] ;
   wire \ram[177][5] ;
   wire \ram[177][4] ;
   wire \ram[177][3] ;
   wire \ram[177][2] ;
   wire \ram[177][1] ;
   wire \ram[177][0] ;
   wire \ram[176][15] ;
   wire \ram[176][14] ;
   wire \ram[176][13] ;
   wire \ram[176][12] ;
   wire \ram[176][11] ;
   wire \ram[176][10] ;
   wire \ram[176][9] ;
   wire \ram[176][8] ;
   wire \ram[176][7] ;
   wire \ram[176][6] ;
   wire \ram[176][5] ;
   wire \ram[176][4] ;
   wire \ram[176][3] ;
   wire \ram[176][2] ;
   wire \ram[176][1] ;
   wire \ram[176][0] ;
   wire \ram[175][15] ;
   wire \ram[175][14] ;
   wire \ram[175][13] ;
   wire \ram[175][12] ;
   wire \ram[175][11] ;
   wire \ram[175][10] ;
   wire \ram[175][9] ;
   wire \ram[175][8] ;
   wire \ram[175][7] ;
   wire \ram[175][6] ;
   wire \ram[175][5] ;
   wire \ram[175][4] ;
   wire \ram[175][3] ;
   wire \ram[175][2] ;
   wire \ram[175][1] ;
   wire \ram[175][0] ;
   wire \ram[174][15] ;
   wire \ram[174][14] ;
   wire \ram[174][13] ;
   wire \ram[174][12] ;
   wire \ram[174][11] ;
   wire \ram[174][10] ;
   wire \ram[174][9] ;
   wire \ram[174][8] ;
   wire \ram[174][7] ;
   wire \ram[174][6] ;
   wire \ram[174][5] ;
   wire \ram[174][4] ;
   wire \ram[174][3] ;
   wire \ram[174][2] ;
   wire \ram[174][1] ;
   wire \ram[174][0] ;
   wire \ram[173][15] ;
   wire \ram[173][14] ;
   wire \ram[173][13] ;
   wire \ram[173][12] ;
   wire \ram[173][11] ;
   wire \ram[173][10] ;
   wire \ram[173][9] ;
   wire \ram[173][8] ;
   wire \ram[173][7] ;
   wire \ram[173][6] ;
   wire \ram[173][5] ;
   wire \ram[173][4] ;
   wire \ram[173][3] ;
   wire \ram[173][2] ;
   wire \ram[173][1] ;
   wire \ram[173][0] ;
   wire \ram[172][15] ;
   wire \ram[172][14] ;
   wire \ram[172][13] ;
   wire \ram[172][12] ;
   wire \ram[172][11] ;
   wire \ram[172][10] ;
   wire \ram[172][9] ;
   wire \ram[172][8] ;
   wire \ram[172][7] ;
   wire \ram[172][6] ;
   wire \ram[172][5] ;
   wire \ram[172][4] ;
   wire \ram[172][3] ;
   wire \ram[172][2] ;
   wire \ram[172][1] ;
   wire \ram[172][0] ;
   wire \ram[171][15] ;
   wire \ram[171][14] ;
   wire \ram[171][13] ;
   wire \ram[171][12] ;
   wire \ram[171][11] ;
   wire \ram[171][10] ;
   wire \ram[171][9] ;
   wire \ram[171][8] ;
   wire \ram[171][7] ;
   wire \ram[171][6] ;
   wire \ram[171][5] ;
   wire \ram[171][4] ;
   wire \ram[171][3] ;
   wire \ram[171][2] ;
   wire \ram[171][1] ;
   wire \ram[171][0] ;
   wire \ram[170][15] ;
   wire \ram[170][14] ;
   wire \ram[170][13] ;
   wire \ram[170][12] ;
   wire \ram[170][11] ;
   wire \ram[170][10] ;
   wire \ram[170][9] ;
   wire \ram[170][8] ;
   wire \ram[170][7] ;
   wire \ram[170][6] ;
   wire \ram[170][5] ;
   wire \ram[170][4] ;
   wire \ram[170][3] ;
   wire \ram[170][2] ;
   wire \ram[170][1] ;
   wire \ram[170][0] ;
   wire \ram[169][15] ;
   wire \ram[169][14] ;
   wire \ram[169][13] ;
   wire \ram[169][12] ;
   wire \ram[169][11] ;
   wire \ram[169][10] ;
   wire \ram[169][9] ;
   wire \ram[169][8] ;
   wire \ram[169][7] ;
   wire \ram[169][6] ;
   wire \ram[169][5] ;
   wire \ram[169][4] ;
   wire \ram[169][3] ;
   wire \ram[169][2] ;
   wire \ram[169][1] ;
   wire \ram[169][0] ;
   wire \ram[168][15] ;
   wire \ram[168][14] ;
   wire \ram[168][13] ;
   wire \ram[168][12] ;
   wire \ram[168][11] ;
   wire \ram[168][10] ;
   wire \ram[168][9] ;
   wire \ram[168][8] ;
   wire \ram[168][7] ;
   wire \ram[168][6] ;
   wire \ram[168][5] ;
   wire \ram[168][4] ;
   wire \ram[168][3] ;
   wire \ram[168][2] ;
   wire \ram[168][1] ;
   wire \ram[168][0] ;
   wire \ram[167][15] ;
   wire \ram[167][14] ;
   wire \ram[167][13] ;
   wire \ram[167][12] ;
   wire \ram[167][11] ;
   wire \ram[167][10] ;
   wire \ram[167][9] ;
   wire \ram[167][8] ;
   wire \ram[167][7] ;
   wire \ram[167][6] ;
   wire \ram[167][5] ;
   wire \ram[167][4] ;
   wire \ram[167][3] ;
   wire \ram[167][2] ;
   wire \ram[167][1] ;
   wire \ram[167][0] ;
   wire \ram[166][15] ;
   wire \ram[166][14] ;
   wire \ram[166][13] ;
   wire \ram[166][12] ;
   wire \ram[166][11] ;
   wire \ram[166][10] ;
   wire \ram[166][9] ;
   wire \ram[166][8] ;
   wire \ram[166][7] ;
   wire \ram[166][6] ;
   wire \ram[166][5] ;
   wire \ram[166][4] ;
   wire \ram[166][3] ;
   wire \ram[166][2] ;
   wire \ram[166][1] ;
   wire \ram[166][0] ;
   wire \ram[165][15] ;
   wire \ram[165][14] ;
   wire \ram[165][13] ;
   wire \ram[165][12] ;
   wire \ram[165][11] ;
   wire \ram[165][10] ;
   wire \ram[165][9] ;
   wire \ram[165][8] ;
   wire \ram[165][7] ;
   wire \ram[165][6] ;
   wire \ram[165][5] ;
   wire \ram[165][4] ;
   wire \ram[165][3] ;
   wire \ram[165][2] ;
   wire \ram[165][1] ;
   wire \ram[165][0] ;
   wire \ram[164][15] ;
   wire \ram[164][14] ;
   wire \ram[164][13] ;
   wire \ram[164][12] ;
   wire \ram[164][11] ;
   wire \ram[164][10] ;
   wire \ram[164][9] ;
   wire \ram[164][8] ;
   wire \ram[164][7] ;
   wire \ram[164][6] ;
   wire \ram[164][5] ;
   wire \ram[164][4] ;
   wire \ram[164][3] ;
   wire \ram[164][2] ;
   wire \ram[164][1] ;
   wire \ram[164][0] ;
   wire \ram[163][15] ;
   wire \ram[163][14] ;
   wire \ram[163][13] ;
   wire \ram[163][12] ;
   wire \ram[163][11] ;
   wire \ram[163][10] ;
   wire \ram[163][9] ;
   wire \ram[163][8] ;
   wire \ram[163][7] ;
   wire \ram[163][6] ;
   wire \ram[163][5] ;
   wire \ram[163][4] ;
   wire \ram[163][3] ;
   wire \ram[163][2] ;
   wire \ram[163][1] ;
   wire \ram[163][0] ;
   wire \ram[162][15] ;
   wire \ram[162][14] ;
   wire \ram[162][13] ;
   wire \ram[162][12] ;
   wire \ram[162][11] ;
   wire \ram[162][10] ;
   wire \ram[162][9] ;
   wire \ram[162][8] ;
   wire \ram[162][7] ;
   wire \ram[162][6] ;
   wire \ram[162][5] ;
   wire \ram[162][4] ;
   wire \ram[162][3] ;
   wire \ram[162][2] ;
   wire \ram[162][1] ;
   wire \ram[162][0] ;
   wire \ram[161][15] ;
   wire \ram[161][14] ;
   wire \ram[161][13] ;
   wire \ram[161][12] ;
   wire \ram[161][11] ;
   wire \ram[161][10] ;
   wire \ram[161][9] ;
   wire \ram[161][8] ;
   wire \ram[161][7] ;
   wire \ram[161][6] ;
   wire \ram[161][5] ;
   wire \ram[161][4] ;
   wire \ram[161][3] ;
   wire \ram[161][2] ;
   wire \ram[161][1] ;
   wire \ram[161][0] ;
   wire \ram[160][15] ;
   wire \ram[160][14] ;
   wire \ram[160][13] ;
   wire \ram[160][12] ;
   wire \ram[160][11] ;
   wire \ram[160][10] ;
   wire \ram[160][9] ;
   wire \ram[160][8] ;
   wire \ram[160][7] ;
   wire \ram[160][6] ;
   wire \ram[160][5] ;
   wire \ram[160][4] ;
   wire \ram[160][3] ;
   wire \ram[160][2] ;
   wire \ram[160][1] ;
   wire \ram[160][0] ;
   wire \ram[159][15] ;
   wire \ram[159][14] ;
   wire \ram[159][13] ;
   wire \ram[159][12] ;
   wire \ram[159][11] ;
   wire \ram[159][10] ;
   wire \ram[159][9] ;
   wire \ram[159][8] ;
   wire \ram[159][7] ;
   wire \ram[159][6] ;
   wire \ram[159][5] ;
   wire \ram[159][4] ;
   wire \ram[159][3] ;
   wire \ram[159][2] ;
   wire \ram[159][1] ;
   wire \ram[159][0] ;
   wire \ram[158][15] ;
   wire \ram[158][14] ;
   wire \ram[158][13] ;
   wire \ram[158][12] ;
   wire \ram[158][11] ;
   wire \ram[158][10] ;
   wire \ram[158][9] ;
   wire \ram[158][8] ;
   wire \ram[158][7] ;
   wire \ram[158][6] ;
   wire \ram[158][5] ;
   wire \ram[158][4] ;
   wire \ram[158][3] ;
   wire \ram[158][2] ;
   wire \ram[158][1] ;
   wire \ram[158][0] ;
   wire \ram[157][15] ;
   wire \ram[157][14] ;
   wire \ram[157][13] ;
   wire \ram[157][12] ;
   wire \ram[157][11] ;
   wire \ram[157][10] ;
   wire \ram[157][9] ;
   wire \ram[157][8] ;
   wire \ram[157][7] ;
   wire \ram[157][6] ;
   wire \ram[157][5] ;
   wire \ram[157][4] ;
   wire \ram[157][3] ;
   wire \ram[157][2] ;
   wire \ram[157][1] ;
   wire \ram[157][0] ;
   wire \ram[156][15] ;
   wire \ram[156][14] ;
   wire \ram[156][13] ;
   wire \ram[156][12] ;
   wire \ram[156][11] ;
   wire \ram[156][10] ;
   wire \ram[156][9] ;
   wire \ram[156][8] ;
   wire \ram[156][7] ;
   wire \ram[156][6] ;
   wire \ram[156][5] ;
   wire \ram[156][4] ;
   wire \ram[156][3] ;
   wire \ram[156][2] ;
   wire \ram[156][1] ;
   wire \ram[156][0] ;
   wire \ram[155][15] ;
   wire \ram[155][14] ;
   wire \ram[155][13] ;
   wire \ram[155][12] ;
   wire \ram[155][11] ;
   wire \ram[155][10] ;
   wire \ram[155][9] ;
   wire \ram[155][8] ;
   wire \ram[155][7] ;
   wire \ram[155][6] ;
   wire \ram[155][5] ;
   wire \ram[155][4] ;
   wire \ram[155][3] ;
   wire \ram[155][2] ;
   wire \ram[155][1] ;
   wire \ram[155][0] ;
   wire \ram[154][15] ;
   wire \ram[154][14] ;
   wire \ram[154][13] ;
   wire \ram[154][12] ;
   wire \ram[154][11] ;
   wire \ram[154][10] ;
   wire \ram[154][9] ;
   wire \ram[154][8] ;
   wire \ram[154][7] ;
   wire \ram[154][6] ;
   wire \ram[154][5] ;
   wire \ram[154][4] ;
   wire \ram[154][3] ;
   wire \ram[154][2] ;
   wire \ram[154][1] ;
   wire \ram[154][0] ;
   wire \ram[153][15] ;
   wire \ram[153][14] ;
   wire \ram[153][13] ;
   wire \ram[153][12] ;
   wire \ram[153][11] ;
   wire \ram[153][10] ;
   wire \ram[153][9] ;
   wire \ram[153][8] ;
   wire \ram[153][7] ;
   wire \ram[153][6] ;
   wire \ram[153][5] ;
   wire \ram[153][4] ;
   wire \ram[153][3] ;
   wire \ram[153][2] ;
   wire \ram[153][1] ;
   wire \ram[153][0] ;
   wire \ram[152][15] ;
   wire \ram[152][14] ;
   wire \ram[152][13] ;
   wire \ram[152][12] ;
   wire \ram[152][11] ;
   wire \ram[152][10] ;
   wire \ram[152][9] ;
   wire \ram[152][8] ;
   wire \ram[152][7] ;
   wire \ram[152][6] ;
   wire \ram[152][5] ;
   wire \ram[152][4] ;
   wire \ram[152][3] ;
   wire \ram[152][2] ;
   wire \ram[152][1] ;
   wire \ram[152][0] ;
   wire \ram[151][15] ;
   wire \ram[151][14] ;
   wire \ram[151][13] ;
   wire \ram[151][12] ;
   wire \ram[151][11] ;
   wire \ram[151][10] ;
   wire \ram[151][9] ;
   wire \ram[151][8] ;
   wire \ram[151][7] ;
   wire \ram[151][6] ;
   wire \ram[151][5] ;
   wire \ram[151][4] ;
   wire \ram[151][3] ;
   wire \ram[151][2] ;
   wire \ram[151][1] ;
   wire \ram[151][0] ;
   wire \ram[150][15] ;
   wire \ram[150][14] ;
   wire \ram[150][13] ;
   wire \ram[150][12] ;
   wire \ram[150][11] ;
   wire \ram[150][10] ;
   wire \ram[150][9] ;
   wire \ram[150][8] ;
   wire \ram[150][7] ;
   wire \ram[150][6] ;
   wire \ram[150][5] ;
   wire \ram[150][4] ;
   wire \ram[150][3] ;
   wire \ram[150][2] ;
   wire \ram[150][1] ;
   wire \ram[150][0] ;
   wire \ram[149][15] ;
   wire \ram[149][14] ;
   wire \ram[149][13] ;
   wire \ram[149][12] ;
   wire \ram[149][11] ;
   wire \ram[149][10] ;
   wire \ram[149][9] ;
   wire \ram[149][8] ;
   wire \ram[149][7] ;
   wire \ram[149][6] ;
   wire \ram[149][5] ;
   wire \ram[149][4] ;
   wire \ram[149][3] ;
   wire \ram[149][2] ;
   wire \ram[149][1] ;
   wire \ram[149][0] ;
   wire \ram[148][15] ;
   wire \ram[148][14] ;
   wire \ram[148][13] ;
   wire \ram[148][12] ;
   wire \ram[148][11] ;
   wire \ram[148][10] ;
   wire \ram[148][9] ;
   wire \ram[148][8] ;
   wire \ram[148][7] ;
   wire \ram[148][6] ;
   wire \ram[148][5] ;
   wire \ram[148][4] ;
   wire \ram[148][3] ;
   wire \ram[148][2] ;
   wire \ram[148][1] ;
   wire \ram[148][0] ;
   wire \ram[147][15] ;
   wire \ram[147][14] ;
   wire \ram[147][13] ;
   wire \ram[147][12] ;
   wire \ram[147][11] ;
   wire \ram[147][10] ;
   wire \ram[147][9] ;
   wire \ram[147][8] ;
   wire \ram[147][7] ;
   wire \ram[147][6] ;
   wire \ram[147][5] ;
   wire \ram[147][4] ;
   wire \ram[147][3] ;
   wire \ram[147][2] ;
   wire \ram[147][1] ;
   wire \ram[147][0] ;
   wire \ram[146][15] ;
   wire \ram[146][14] ;
   wire \ram[146][13] ;
   wire \ram[146][12] ;
   wire \ram[146][11] ;
   wire \ram[146][10] ;
   wire \ram[146][9] ;
   wire \ram[146][8] ;
   wire \ram[146][7] ;
   wire \ram[146][6] ;
   wire \ram[146][5] ;
   wire \ram[146][4] ;
   wire \ram[146][3] ;
   wire \ram[146][2] ;
   wire \ram[146][1] ;
   wire \ram[146][0] ;
   wire \ram[145][15] ;
   wire \ram[145][14] ;
   wire \ram[145][13] ;
   wire \ram[145][12] ;
   wire \ram[145][11] ;
   wire \ram[145][10] ;
   wire \ram[145][9] ;
   wire \ram[145][8] ;
   wire \ram[145][7] ;
   wire \ram[145][6] ;
   wire \ram[145][5] ;
   wire \ram[145][4] ;
   wire \ram[145][3] ;
   wire \ram[145][2] ;
   wire \ram[145][1] ;
   wire \ram[145][0] ;
   wire \ram[144][15] ;
   wire \ram[144][14] ;
   wire \ram[144][13] ;
   wire \ram[144][12] ;
   wire \ram[144][11] ;
   wire \ram[144][10] ;
   wire \ram[144][9] ;
   wire \ram[144][8] ;
   wire \ram[144][7] ;
   wire \ram[144][6] ;
   wire \ram[144][5] ;
   wire \ram[144][4] ;
   wire \ram[144][3] ;
   wire \ram[144][2] ;
   wire \ram[144][1] ;
   wire \ram[144][0] ;
   wire \ram[143][15] ;
   wire \ram[143][14] ;
   wire \ram[143][13] ;
   wire \ram[143][12] ;
   wire \ram[143][11] ;
   wire \ram[143][10] ;
   wire \ram[143][9] ;
   wire \ram[143][8] ;
   wire \ram[143][7] ;
   wire \ram[143][6] ;
   wire \ram[143][5] ;
   wire \ram[143][4] ;
   wire \ram[143][3] ;
   wire \ram[143][2] ;
   wire \ram[143][1] ;
   wire \ram[143][0] ;
   wire \ram[142][15] ;
   wire \ram[142][14] ;
   wire \ram[142][13] ;
   wire \ram[142][12] ;
   wire \ram[142][11] ;
   wire \ram[142][10] ;
   wire \ram[142][9] ;
   wire \ram[142][8] ;
   wire \ram[142][7] ;
   wire \ram[142][6] ;
   wire \ram[142][5] ;
   wire \ram[142][4] ;
   wire \ram[142][3] ;
   wire \ram[142][2] ;
   wire \ram[142][1] ;
   wire \ram[142][0] ;
   wire \ram[141][15] ;
   wire \ram[141][14] ;
   wire \ram[141][13] ;
   wire \ram[141][12] ;
   wire \ram[141][11] ;
   wire \ram[141][10] ;
   wire \ram[141][9] ;
   wire \ram[141][8] ;
   wire \ram[141][7] ;
   wire \ram[141][6] ;
   wire \ram[141][5] ;
   wire \ram[141][4] ;
   wire \ram[141][3] ;
   wire \ram[141][2] ;
   wire \ram[141][1] ;
   wire \ram[141][0] ;
   wire \ram[140][15] ;
   wire \ram[140][14] ;
   wire \ram[140][13] ;
   wire \ram[140][12] ;
   wire \ram[140][11] ;
   wire \ram[140][10] ;
   wire \ram[140][9] ;
   wire \ram[140][8] ;
   wire \ram[140][7] ;
   wire \ram[140][6] ;
   wire \ram[140][5] ;
   wire \ram[140][4] ;
   wire \ram[140][3] ;
   wire \ram[140][2] ;
   wire \ram[140][1] ;
   wire \ram[140][0] ;
   wire \ram[139][15] ;
   wire \ram[139][14] ;
   wire \ram[139][13] ;
   wire \ram[139][12] ;
   wire \ram[139][11] ;
   wire \ram[139][10] ;
   wire \ram[139][9] ;
   wire \ram[139][8] ;
   wire \ram[139][7] ;
   wire \ram[139][6] ;
   wire \ram[139][5] ;
   wire \ram[139][4] ;
   wire \ram[139][3] ;
   wire \ram[139][2] ;
   wire \ram[139][1] ;
   wire \ram[139][0] ;
   wire \ram[138][15] ;
   wire \ram[138][14] ;
   wire \ram[138][13] ;
   wire \ram[138][12] ;
   wire \ram[138][11] ;
   wire \ram[138][10] ;
   wire \ram[138][9] ;
   wire \ram[138][8] ;
   wire \ram[138][7] ;
   wire \ram[138][6] ;
   wire \ram[138][5] ;
   wire \ram[138][4] ;
   wire \ram[138][3] ;
   wire \ram[138][2] ;
   wire \ram[138][1] ;
   wire \ram[138][0] ;
   wire \ram[137][15] ;
   wire \ram[137][14] ;
   wire \ram[137][13] ;
   wire \ram[137][12] ;
   wire \ram[137][11] ;
   wire \ram[137][10] ;
   wire \ram[137][9] ;
   wire \ram[137][8] ;
   wire \ram[137][7] ;
   wire \ram[137][6] ;
   wire \ram[137][5] ;
   wire \ram[137][4] ;
   wire \ram[137][3] ;
   wire \ram[137][2] ;
   wire \ram[137][1] ;
   wire \ram[137][0] ;
   wire \ram[136][15] ;
   wire \ram[136][14] ;
   wire \ram[136][13] ;
   wire \ram[136][12] ;
   wire \ram[136][11] ;
   wire \ram[136][10] ;
   wire \ram[136][9] ;
   wire \ram[136][8] ;
   wire \ram[136][7] ;
   wire \ram[136][6] ;
   wire \ram[136][5] ;
   wire \ram[136][4] ;
   wire \ram[136][3] ;
   wire \ram[136][2] ;
   wire \ram[136][1] ;
   wire \ram[136][0] ;
   wire \ram[135][15] ;
   wire \ram[135][14] ;
   wire \ram[135][13] ;
   wire \ram[135][12] ;
   wire \ram[135][11] ;
   wire \ram[135][10] ;
   wire \ram[135][9] ;
   wire \ram[135][8] ;
   wire \ram[135][7] ;
   wire \ram[135][6] ;
   wire \ram[135][5] ;
   wire \ram[135][4] ;
   wire \ram[135][3] ;
   wire \ram[135][2] ;
   wire \ram[135][1] ;
   wire \ram[135][0] ;
   wire \ram[134][15] ;
   wire \ram[134][14] ;
   wire \ram[134][13] ;
   wire \ram[134][12] ;
   wire \ram[134][11] ;
   wire \ram[134][10] ;
   wire \ram[134][9] ;
   wire \ram[134][8] ;
   wire \ram[134][7] ;
   wire \ram[134][6] ;
   wire \ram[134][5] ;
   wire \ram[134][4] ;
   wire \ram[134][3] ;
   wire \ram[134][2] ;
   wire \ram[134][1] ;
   wire \ram[134][0] ;
   wire \ram[133][15] ;
   wire \ram[133][14] ;
   wire \ram[133][13] ;
   wire \ram[133][12] ;
   wire \ram[133][11] ;
   wire \ram[133][10] ;
   wire \ram[133][9] ;
   wire \ram[133][8] ;
   wire \ram[133][7] ;
   wire \ram[133][6] ;
   wire \ram[133][5] ;
   wire \ram[133][4] ;
   wire \ram[133][3] ;
   wire \ram[133][2] ;
   wire \ram[133][1] ;
   wire \ram[133][0] ;
   wire \ram[132][15] ;
   wire \ram[132][14] ;
   wire \ram[132][13] ;
   wire \ram[132][12] ;
   wire \ram[132][11] ;
   wire \ram[132][10] ;
   wire \ram[132][9] ;
   wire \ram[132][8] ;
   wire \ram[132][7] ;
   wire \ram[132][6] ;
   wire \ram[132][5] ;
   wire \ram[132][4] ;
   wire \ram[132][3] ;
   wire \ram[132][2] ;
   wire \ram[132][1] ;
   wire \ram[132][0] ;
   wire \ram[131][15] ;
   wire \ram[131][14] ;
   wire \ram[131][13] ;
   wire \ram[131][12] ;
   wire \ram[131][11] ;
   wire \ram[131][10] ;
   wire \ram[131][9] ;
   wire \ram[131][8] ;
   wire \ram[131][7] ;
   wire \ram[131][6] ;
   wire \ram[131][5] ;
   wire \ram[131][4] ;
   wire \ram[131][3] ;
   wire \ram[131][2] ;
   wire \ram[131][1] ;
   wire \ram[131][0] ;
   wire \ram[130][15] ;
   wire \ram[130][14] ;
   wire \ram[130][13] ;
   wire \ram[130][12] ;
   wire \ram[130][11] ;
   wire \ram[130][10] ;
   wire \ram[130][9] ;
   wire \ram[130][8] ;
   wire \ram[130][7] ;
   wire \ram[130][6] ;
   wire \ram[130][5] ;
   wire \ram[130][4] ;
   wire \ram[130][3] ;
   wire \ram[130][2] ;
   wire \ram[130][1] ;
   wire \ram[130][0] ;
   wire \ram[129][15] ;
   wire \ram[129][14] ;
   wire \ram[129][13] ;
   wire \ram[129][12] ;
   wire \ram[129][11] ;
   wire \ram[129][10] ;
   wire \ram[129][9] ;
   wire \ram[129][8] ;
   wire \ram[129][7] ;
   wire \ram[129][6] ;
   wire \ram[129][5] ;
   wire \ram[129][4] ;
   wire \ram[129][3] ;
   wire \ram[129][2] ;
   wire \ram[129][1] ;
   wire \ram[129][0] ;
   wire \ram[128][15] ;
   wire \ram[128][14] ;
   wire \ram[128][13] ;
   wire \ram[128][12] ;
   wire \ram[128][11] ;
   wire \ram[128][10] ;
   wire \ram[128][9] ;
   wire \ram[128][8] ;
   wire \ram[128][7] ;
   wire \ram[128][6] ;
   wire \ram[128][5] ;
   wire \ram[128][4] ;
   wire \ram[128][3] ;
   wire \ram[128][2] ;
   wire \ram[128][1] ;
   wire \ram[128][0] ;
   wire \ram[127][15] ;
   wire \ram[127][14] ;
   wire \ram[127][13] ;
   wire \ram[127][12] ;
   wire \ram[127][11] ;
   wire \ram[127][10] ;
   wire \ram[127][9] ;
   wire \ram[127][8] ;
   wire \ram[127][7] ;
   wire \ram[127][6] ;
   wire \ram[127][5] ;
   wire \ram[127][4] ;
   wire \ram[127][3] ;
   wire \ram[127][2] ;
   wire \ram[127][1] ;
   wire \ram[127][0] ;
   wire \ram[126][15] ;
   wire \ram[126][14] ;
   wire \ram[126][13] ;
   wire \ram[126][12] ;
   wire \ram[126][11] ;
   wire \ram[126][10] ;
   wire \ram[126][9] ;
   wire \ram[126][8] ;
   wire \ram[126][7] ;
   wire \ram[126][6] ;
   wire \ram[126][5] ;
   wire \ram[126][4] ;
   wire \ram[126][3] ;
   wire \ram[126][2] ;
   wire \ram[126][1] ;
   wire \ram[126][0] ;
   wire \ram[125][15] ;
   wire \ram[125][14] ;
   wire \ram[125][13] ;
   wire \ram[125][12] ;
   wire \ram[125][11] ;
   wire \ram[125][10] ;
   wire \ram[125][9] ;
   wire \ram[125][8] ;
   wire \ram[125][7] ;
   wire \ram[125][6] ;
   wire \ram[125][5] ;
   wire \ram[125][4] ;
   wire \ram[125][3] ;
   wire \ram[125][2] ;
   wire \ram[125][1] ;
   wire \ram[125][0] ;
   wire \ram[124][15] ;
   wire \ram[124][14] ;
   wire \ram[124][13] ;
   wire \ram[124][12] ;
   wire \ram[124][11] ;
   wire \ram[124][10] ;
   wire \ram[124][9] ;
   wire \ram[124][8] ;
   wire \ram[124][7] ;
   wire \ram[124][6] ;
   wire \ram[124][5] ;
   wire \ram[124][4] ;
   wire \ram[124][3] ;
   wire \ram[124][2] ;
   wire \ram[124][1] ;
   wire \ram[124][0] ;
   wire \ram[123][15] ;
   wire \ram[123][14] ;
   wire \ram[123][13] ;
   wire \ram[123][12] ;
   wire \ram[123][11] ;
   wire \ram[123][10] ;
   wire \ram[123][9] ;
   wire \ram[123][8] ;
   wire \ram[123][7] ;
   wire \ram[123][6] ;
   wire \ram[123][5] ;
   wire \ram[123][4] ;
   wire \ram[123][3] ;
   wire \ram[123][2] ;
   wire \ram[123][1] ;
   wire \ram[123][0] ;
   wire \ram[122][15] ;
   wire \ram[122][14] ;
   wire \ram[122][13] ;
   wire \ram[122][12] ;
   wire \ram[122][11] ;
   wire \ram[122][10] ;
   wire \ram[122][9] ;
   wire \ram[122][8] ;
   wire \ram[122][7] ;
   wire \ram[122][6] ;
   wire \ram[122][5] ;
   wire \ram[122][4] ;
   wire \ram[122][3] ;
   wire \ram[122][2] ;
   wire \ram[122][1] ;
   wire \ram[122][0] ;
   wire \ram[121][15] ;
   wire \ram[121][14] ;
   wire \ram[121][13] ;
   wire \ram[121][12] ;
   wire \ram[121][11] ;
   wire \ram[121][10] ;
   wire \ram[121][9] ;
   wire \ram[121][8] ;
   wire \ram[121][7] ;
   wire \ram[121][6] ;
   wire \ram[121][5] ;
   wire \ram[121][4] ;
   wire \ram[121][3] ;
   wire \ram[121][2] ;
   wire \ram[121][1] ;
   wire \ram[121][0] ;
   wire \ram[120][15] ;
   wire \ram[120][14] ;
   wire \ram[120][13] ;
   wire \ram[120][12] ;
   wire \ram[120][11] ;
   wire \ram[120][10] ;
   wire \ram[120][9] ;
   wire \ram[120][8] ;
   wire \ram[120][7] ;
   wire \ram[120][6] ;
   wire \ram[120][5] ;
   wire \ram[120][4] ;
   wire \ram[120][3] ;
   wire \ram[120][2] ;
   wire \ram[120][1] ;
   wire \ram[120][0] ;
   wire \ram[119][15] ;
   wire \ram[119][14] ;
   wire \ram[119][13] ;
   wire \ram[119][12] ;
   wire \ram[119][11] ;
   wire \ram[119][10] ;
   wire \ram[119][9] ;
   wire \ram[119][8] ;
   wire \ram[119][7] ;
   wire \ram[119][6] ;
   wire \ram[119][5] ;
   wire \ram[119][4] ;
   wire \ram[119][3] ;
   wire \ram[119][2] ;
   wire \ram[119][1] ;
   wire \ram[119][0] ;
   wire \ram[118][15] ;
   wire \ram[118][14] ;
   wire \ram[118][13] ;
   wire \ram[118][12] ;
   wire \ram[118][11] ;
   wire \ram[118][10] ;
   wire \ram[118][9] ;
   wire \ram[118][8] ;
   wire \ram[118][7] ;
   wire \ram[118][6] ;
   wire \ram[118][5] ;
   wire \ram[118][4] ;
   wire \ram[118][3] ;
   wire \ram[118][2] ;
   wire \ram[118][1] ;
   wire \ram[118][0] ;
   wire \ram[117][15] ;
   wire \ram[117][14] ;
   wire \ram[117][13] ;
   wire \ram[117][12] ;
   wire \ram[117][11] ;
   wire \ram[117][10] ;
   wire \ram[117][9] ;
   wire \ram[117][8] ;
   wire \ram[117][7] ;
   wire \ram[117][6] ;
   wire \ram[117][5] ;
   wire \ram[117][4] ;
   wire \ram[117][3] ;
   wire \ram[117][2] ;
   wire \ram[117][1] ;
   wire \ram[117][0] ;
   wire \ram[116][15] ;
   wire \ram[116][14] ;
   wire \ram[116][13] ;
   wire \ram[116][12] ;
   wire \ram[116][11] ;
   wire \ram[116][10] ;
   wire \ram[116][9] ;
   wire \ram[116][8] ;
   wire \ram[116][7] ;
   wire \ram[116][6] ;
   wire \ram[116][5] ;
   wire \ram[116][4] ;
   wire \ram[116][3] ;
   wire \ram[116][2] ;
   wire \ram[116][1] ;
   wire \ram[116][0] ;
   wire \ram[115][15] ;
   wire \ram[115][14] ;
   wire \ram[115][13] ;
   wire \ram[115][12] ;
   wire \ram[115][11] ;
   wire \ram[115][10] ;
   wire \ram[115][9] ;
   wire \ram[115][8] ;
   wire \ram[115][7] ;
   wire \ram[115][6] ;
   wire \ram[115][5] ;
   wire \ram[115][4] ;
   wire \ram[115][3] ;
   wire \ram[115][2] ;
   wire \ram[115][1] ;
   wire \ram[115][0] ;
   wire \ram[114][15] ;
   wire \ram[114][14] ;
   wire \ram[114][13] ;
   wire \ram[114][12] ;
   wire \ram[114][11] ;
   wire \ram[114][10] ;
   wire \ram[114][9] ;
   wire \ram[114][8] ;
   wire \ram[114][7] ;
   wire \ram[114][6] ;
   wire \ram[114][5] ;
   wire \ram[114][4] ;
   wire \ram[114][3] ;
   wire \ram[114][2] ;
   wire \ram[114][1] ;
   wire \ram[114][0] ;
   wire \ram[113][15] ;
   wire \ram[113][14] ;
   wire \ram[113][13] ;
   wire \ram[113][12] ;
   wire \ram[113][11] ;
   wire \ram[113][10] ;
   wire \ram[113][9] ;
   wire \ram[113][8] ;
   wire \ram[113][7] ;
   wire \ram[113][6] ;
   wire \ram[113][5] ;
   wire \ram[113][4] ;
   wire \ram[113][3] ;
   wire \ram[113][2] ;
   wire \ram[113][1] ;
   wire \ram[113][0] ;
   wire \ram[112][15] ;
   wire \ram[112][14] ;
   wire \ram[112][13] ;
   wire \ram[112][12] ;
   wire \ram[112][11] ;
   wire \ram[112][10] ;
   wire \ram[112][9] ;
   wire \ram[112][8] ;
   wire \ram[112][7] ;
   wire \ram[112][6] ;
   wire \ram[112][5] ;
   wire \ram[112][4] ;
   wire \ram[112][3] ;
   wire \ram[112][2] ;
   wire \ram[112][1] ;
   wire \ram[112][0] ;
   wire \ram[111][15] ;
   wire \ram[111][14] ;
   wire \ram[111][13] ;
   wire \ram[111][12] ;
   wire \ram[111][11] ;
   wire \ram[111][10] ;
   wire \ram[111][9] ;
   wire \ram[111][8] ;
   wire \ram[111][7] ;
   wire \ram[111][6] ;
   wire \ram[111][5] ;
   wire \ram[111][4] ;
   wire \ram[111][3] ;
   wire \ram[111][2] ;
   wire \ram[111][1] ;
   wire \ram[111][0] ;
   wire \ram[110][15] ;
   wire \ram[110][14] ;
   wire \ram[110][13] ;
   wire \ram[110][12] ;
   wire \ram[110][11] ;
   wire \ram[110][10] ;
   wire \ram[110][9] ;
   wire \ram[110][8] ;
   wire \ram[110][7] ;
   wire \ram[110][6] ;
   wire \ram[110][5] ;
   wire \ram[110][4] ;
   wire \ram[110][3] ;
   wire \ram[110][2] ;
   wire \ram[110][1] ;
   wire \ram[110][0] ;
   wire \ram[109][15] ;
   wire \ram[109][14] ;
   wire \ram[109][13] ;
   wire \ram[109][12] ;
   wire \ram[109][11] ;
   wire \ram[109][10] ;
   wire \ram[109][9] ;
   wire \ram[109][8] ;
   wire \ram[109][7] ;
   wire \ram[109][6] ;
   wire \ram[109][5] ;
   wire \ram[109][4] ;
   wire \ram[109][3] ;
   wire \ram[109][2] ;
   wire \ram[109][1] ;
   wire \ram[109][0] ;
   wire \ram[108][15] ;
   wire \ram[108][14] ;
   wire \ram[108][13] ;
   wire \ram[108][12] ;
   wire \ram[108][11] ;
   wire \ram[108][10] ;
   wire \ram[108][9] ;
   wire \ram[108][8] ;
   wire \ram[108][7] ;
   wire \ram[108][6] ;
   wire \ram[108][5] ;
   wire \ram[108][4] ;
   wire \ram[108][3] ;
   wire \ram[108][2] ;
   wire \ram[108][1] ;
   wire \ram[108][0] ;
   wire \ram[107][15] ;
   wire \ram[107][14] ;
   wire \ram[107][13] ;
   wire \ram[107][12] ;
   wire \ram[107][11] ;
   wire \ram[107][10] ;
   wire \ram[107][9] ;
   wire \ram[107][8] ;
   wire \ram[107][7] ;
   wire \ram[107][6] ;
   wire \ram[107][5] ;
   wire \ram[107][4] ;
   wire \ram[107][3] ;
   wire \ram[107][2] ;
   wire \ram[107][1] ;
   wire \ram[107][0] ;
   wire \ram[106][15] ;
   wire \ram[106][14] ;
   wire \ram[106][13] ;
   wire \ram[106][12] ;
   wire \ram[106][11] ;
   wire \ram[106][10] ;
   wire \ram[106][9] ;
   wire \ram[106][8] ;
   wire \ram[106][7] ;
   wire \ram[106][6] ;
   wire \ram[106][5] ;
   wire \ram[106][4] ;
   wire \ram[106][3] ;
   wire \ram[106][2] ;
   wire \ram[106][1] ;
   wire \ram[106][0] ;
   wire \ram[105][15] ;
   wire \ram[105][14] ;
   wire \ram[105][13] ;
   wire \ram[105][12] ;
   wire \ram[105][11] ;
   wire \ram[105][10] ;
   wire \ram[105][9] ;
   wire \ram[105][8] ;
   wire \ram[105][7] ;
   wire \ram[105][6] ;
   wire \ram[105][5] ;
   wire \ram[105][4] ;
   wire \ram[105][3] ;
   wire \ram[105][2] ;
   wire \ram[105][1] ;
   wire \ram[105][0] ;
   wire \ram[104][15] ;
   wire \ram[104][14] ;
   wire \ram[104][13] ;
   wire \ram[104][12] ;
   wire \ram[104][11] ;
   wire \ram[104][10] ;
   wire \ram[104][9] ;
   wire \ram[104][8] ;
   wire \ram[104][7] ;
   wire \ram[104][6] ;
   wire \ram[104][5] ;
   wire \ram[104][4] ;
   wire \ram[104][3] ;
   wire \ram[104][2] ;
   wire \ram[104][1] ;
   wire \ram[104][0] ;
   wire \ram[103][15] ;
   wire \ram[103][14] ;
   wire \ram[103][13] ;
   wire \ram[103][12] ;
   wire \ram[103][11] ;
   wire \ram[103][10] ;
   wire \ram[103][9] ;
   wire \ram[103][8] ;
   wire \ram[103][7] ;
   wire \ram[103][6] ;
   wire \ram[103][5] ;
   wire \ram[103][4] ;
   wire \ram[103][3] ;
   wire \ram[103][2] ;
   wire \ram[103][1] ;
   wire \ram[103][0] ;
   wire \ram[102][15] ;
   wire \ram[102][14] ;
   wire \ram[102][13] ;
   wire \ram[102][12] ;
   wire \ram[102][11] ;
   wire \ram[102][10] ;
   wire \ram[102][9] ;
   wire \ram[102][8] ;
   wire \ram[102][7] ;
   wire \ram[102][6] ;
   wire \ram[102][5] ;
   wire \ram[102][4] ;
   wire \ram[102][3] ;
   wire \ram[102][2] ;
   wire \ram[102][1] ;
   wire \ram[102][0] ;
   wire \ram[101][15] ;
   wire \ram[101][14] ;
   wire \ram[101][13] ;
   wire \ram[101][12] ;
   wire \ram[101][11] ;
   wire \ram[101][10] ;
   wire \ram[101][9] ;
   wire \ram[101][8] ;
   wire \ram[101][7] ;
   wire \ram[101][6] ;
   wire \ram[101][5] ;
   wire \ram[101][4] ;
   wire \ram[101][3] ;
   wire \ram[101][2] ;
   wire \ram[101][1] ;
   wire \ram[101][0] ;
   wire \ram[100][15] ;
   wire \ram[100][14] ;
   wire \ram[100][13] ;
   wire \ram[100][12] ;
   wire \ram[100][11] ;
   wire \ram[100][10] ;
   wire \ram[100][9] ;
   wire \ram[100][8] ;
   wire \ram[100][7] ;
   wire \ram[100][6] ;
   wire \ram[100][5] ;
   wire \ram[100][4] ;
   wire \ram[100][3] ;
   wire \ram[100][2] ;
   wire \ram[100][1] ;
   wire \ram[100][0] ;
   wire \ram[99][15] ;
   wire \ram[99][14] ;
   wire \ram[99][13] ;
   wire \ram[99][12] ;
   wire \ram[99][11] ;
   wire \ram[99][10] ;
   wire \ram[99][9] ;
   wire \ram[99][8] ;
   wire \ram[99][7] ;
   wire \ram[99][6] ;
   wire \ram[99][5] ;
   wire \ram[99][4] ;
   wire \ram[99][3] ;
   wire \ram[99][2] ;
   wire \ram[99][1] ;
   wire \ram[99][0] ;
   wire \ram[98][15] ;
   wire \ram[98][14] ;
   wire \ram[98][13] ;
   wire \ram[98][12] ;
   wire \ram[98][11] ;
   wire \ram[98][10] ;
   wire \ram[98][9] ;
   wire \ram[98][8] ;
   wire \ram[98][7] ;
   wire \ram[98][6] ;
   wire \ram[98][5] ;
   wire \ram[98][4] ;
   wire \ram[98][3] ;
   wire \ram[98][2] ;
   wire \ram[98][1] ;
   wire \ram[98][0] ;
   wire \ram[97][15] ;
   wire \ram[97][14] ;
   wire \ram[97][13] ;
   wire \ram[97][12] ;
   wire \ram[97][11] ;
   wire \ram[97][10] ;
   wire \ram[97][9] ;
   wire \ram[97][8] ;
   wire \ram[97][7] ;
   wire \ram[97][6] ;
   wire \ram[97][5] ;
   wire \ram[97][4] ;
   wire \ram[97][3] ;
   wire \ram[97][2] ;
   wire \ram[97][1] ;
   wire \ram[97][0] ;
   wire \ram[96][15] ;
   wire \ram[96][14] ;
   wire \ram[96][13] ;
   wire \ram[96][12] ;
   wire \ram[96][11] ;
   wire \ram[96][10] ;
   wire \ram[96][9] ;
   wire \ram[96][8] ;
   wire \ram[96][7] ;
   wire \ram[96][6] ;
   wire \ram[96][5] ;
   wire \ram[96][4] ;
   wire \ram[96][3] ;
   wire \ram[96][2] ;
   wire \ram[96][1] ;
   wire \ram[96][0] ;
   wire \ram[95][15] ;
   wire \ram[95][14] ;
   wire \ram[95][13] ;
   wire \ram[95][12] ;
   wire \ram[95][11] ;
   wire \ram[95][10] ;
   wire \ram[95][9] ;
   wire \ram[95][8] ;
   wire \ram[95][7] ;
   wire \ram[95][6] ;
   wire \ram[95][5] ;
   wire \ram[95][4] ;
   wire \ram[95][3] ;
   wire \ram[95][2] ;
   wire \ram[95][1] ;
   wire \ram[95][0] ;
   wire \ram[94][15] ;
   wire \ram[94][14] ;
   wire \ram[94][13] ;
   wire \ram[94][12] ;
   wire \ram[94][11] ;
   wire \ram[94][10] ;
   wire \ram[94][9] ;
   wire \ram[94][8] ;
   wire \ram[94][7] ;
   wire \ram[94][6] ;
   wire \ram[94][5] ;
   wire \ram[94][4] ;
   wire \ram[94][3] ;
   wire \ram[94][2] ;
   wire \ram[94][1] ;
   wire \ram[94][0] ;
   wire \ram[93][15] ;
   wire \ram[93][14] ;
   wire \ram[93][13] ;
   wire \ram[93][12] ;
   wire \ram[93][11] ;
   wire \ram[93][10] ;
   wire \ram[93][9] ;
   wire \ram[93][8] ;
   wire \ram[93][7] ;
   wire \ram[93][6] ;
   wire \ram[93][5] ;
   wire \ram[93][4] ;
   wire \ram[93][3] ;
   wire \ram[93][2] ;
   wire \ram[93][1] ;
   wire \ram[93][0] ;
   wire \ram[92][15] ;
   wire \ram[92][14] ;
   wire \ram[92][13] ;
   wire \ram[92][12] ;
   wire \ram[92][11] ;
   wire \ram[92][10] ;
   wire \ram[92][9] ;
   wire \ram[92][8] ;
   wire \ram[92][7] ;
   wire \ram[92][6] ;
   wire \ram[92][5] ;
   wire \ram[92][4] ;
   wire \ram[92][3] ;
   wire \ram[92][2] ;
   wire \ram[92][1] ;
   wire \ram[92][0] ;
   wire \ram[91][15] ;
   wire \ram[91][14] ;
   wire \ram[91][13] ;
   wire \ram[91][12] ;
   wire \ram[91][11] ;
   wire \ram[91][10] ;
   wire \ram[91][9] ;
   wire \ram[91][8] ;
   wire \ram[91][7] ;
   wire \ram[91][6] ;
   wire \ram[91][5] ;
   wire \ram[91][4] ;
   wire \ram[91][3] ;
   wire \ram[91][2] ;
   wire \ram[91][1] ;
   wire \ram[91][0] ;
   wire \ram[90][15] ;
   wire \ram[90][14] ;
   wire \ram[90][13] ;
   wire \ram[90][12] ;
   wire \ram[90][11] ;
   wire \ram[90][10] ;
   wire \ram[90][9] ;
   wire \ram[90][8] ;
   wire \ram[90][7] ;
   wire \ram[90][6] ;
   wire \ram[90][5] ;
   wire \ram[90][4] ;
   wire \ram[90][3] ;
   wire \ram[90][2] ;
   wire \ram[90][1] ;
   wire \ram[90][0] ;
   wire \ram[89][15] ;
   wire \ram[89][14] ;
   wire \ram[89][13] ;
   wire \ram[89][12] ;
   wire \ram[89][11] ;
   wire \ram[89][10] ;
   wire \ram[89][9] ;
   wire \ram[89][8] ;
   wire \ram[89][7] ;
   wire \ram[89][6] ;
   wire \ram[89][5] ;
   wire \ram[89][4] ;
   wire \ram[89][3] ;
   wire \ram[89][2] ;
   wire \ram[89][1] ;
   wire \ram[89][0] ;
   wire \ram[88][15] ;
   wire \ram[88][14] ;
   wire \ram[88][13] ;
   wire \ram[88][12] ;
   wire \ram[88][11] ;
   wire \ram[88][10] ;
   wire \ram[88][9] ;
   wire \ram[88][8] ;
   wire \ram[88][7] ;
   wire \ram[88][6] ;
   wire \ram[88][5] ;
   wire \ram[88][4] ;
   wire \ram[88][3] ;
   wire \ram[88][2] ;
   wire \ram[88][1] ;
   wire \ram[88][0] ;
   wire \ram[87][15] ;
   wire \ram[87][14] ;
   wire \ram[87][13] ;
   wire \ram[87][12] ;
   wire \ram[87][11] ;
   wire \ram[87][10] ;
   wire \ram[87][9] ;
   wire \ram[87][8] ;
   wire \ram[87][7] ;
   wire \ram[87][6] ;
   wire \ram[87][5] ;
   wire \ram[87][4] ;
   wire \ram[87][3] ;
   wire \ram[87][2] ;
   wire \ram[87][1] ;
   wire \ram[87][0] ;
   wire \ram[86][15] ;
   wire \ram[86][14] ;
   wire \ram[86][13] ;
   wire \ram[86][12] ;
   wire \ram[86][11] ;
   wire \ram[86][10] ;
   wire \ram[86][9] ;
   wire \ram[86][8] ;
   wire \ram[86][7] ;
   wire \ram[86][6] ;
   wire \ram[86][5] ;
   wire \ram[86][4] ;
   wire \ram[86][3] ;
   wire \ram[86][2] ;
   wire \ram[86][1] ;
   wire \ram[86][0] ;
   wire \ram[85][15] ;
   wire \ram[85][14] ;
   wire \ram[85][13] ;
   wire \ram[85][12] ;
   wire \ram[85][11] ;
   wire \ram[85][10] ;
   wire \ram[85][9] ;
   wire \ram[85][8] ;
   wire \ram[85][7] ;
   wire \ram[85][6] ;
   wire \ram[85][5] ;
   wire \ram[85][4] ;
   wire \ram[85][3] ;
   wire \ram[85][2] ;
   wire \ram[85][1] ;
   wire \ram[85][0] ;
   wire \ram[84][15] ;
   wire \ram[84][14] ;
   wire \ram[84][13] ;
   wire \ram[84][12] ;
   wire \ram[84][11] ;
   wire \ram[84][10] ;
   wire \ram[84][9] ;
   wire \ram[84][8] ;
   wire \ram[84][7] ;
   wire \ram[84][6] ;
   wire \ram[84][5] ;
   wire \ram[84][4] ;
   wire \ram[84][3] ;
   wire \ram[84][2] ;
   wire \ram[84][1] ;
   wire \ram[84][0] ;
   wire \ram[83][15] ;
   wire \ram[83][14] ;
   wire \ram[83][13] ;
   wire \ram[83][12] ;
   wire \ram[83][11] ;
   wire \ram[83][10] ;
   wire \ram[83][9] ;
   wire \ram[83][8] ;
   wire \ram[83][7] ;
   wire \ram[83][6] ;
   wire \ram[83][5] ;
   wire \ram[83][4] ;
   wire \ram[83][3] ;
   wire \ram[83][2] ;
   wire \ram[83][1] ;
   wire \ram[83][0] ;
   wire \ram[82][15] ;
   wire \ram[82][14] ;
   wire \ram[82][13] ;
   wire \ram[82][12] ;
   wire \ram[82][11] ;
   wire \ram[82][10] ;
   wire \ram[82][9] ;
   wire \ram[82][8] ;
   wire \ram[82][7] ;
   wire \ram[82][6] ;
   wire \ram[82][5] ;
   wire \ram[82][4] ;
   wire \ram[82][3] ;
   wire \ram[82][2] ;
   wire \ram[82][1] ;
   wire \ram[82][0] ;
   wire \ram[81][15] ;
   wire \ram[81][14] ;
   wire \ram[81][13] ;
   wire \ram[81][12] ;
   wire \ram[81][11] ;
   wire \ram[81][10] ;
   wire \ram[81][9] ;
   wire \ram[81][8] ;
   wire \ram[81][7] ;
   wire \ram[81][6] ;
   wire \ram[81][5] ;
   wire \ram[81][4] ;
   wire \ram[81][3] ;
   wire \ram[81][2] ;
   wire \ram[81][1] ;
   wire \ram[81][0] ;
   wire \ram[80][15] ;
   wire \ram[80][14] ;
   wire \ram[80][13] ;
   wire \ram[80][12] ;
   wire \ram[80][11] ;
   wire \ram[80][10] ;
   wire \ram[80][9] ;
   wire \ram[80][8] ;
   wire \ram[80][7] ;
   wire \ram[80][6] ;
   wire \ram[80][5] ;
   wire \ram[80][4] ;
   wire \ram[80][3] ;
   wire \ram[80][2] ;
   wire \ram[80][1] ;
   wire \ram[80][0] ;
   wire \ram[79][15] ;
   wire \ram[79][14] ;
   wire \ram[79][13] ;
   wire \ram[79][12] ;
   wire \ram[79][11] ;
   wire \ram[79][10] ;
   wire \ram[79][9] ;
   wire \ram[79][8] ;
   wire \ram[79][7] ;
   wire \ram[79][6] ;
   wire \ram[79][5] ;
   wire \ram[79][4] ;
   wire \ram[79][3] ;
   wire \ram[79][2] ;
   wire \ram[79][1] ;
   wire \ram[79][0] ;
   wire \ram[78][15] ;
   wire \ram[78][14] ;
   wire \ram[78][13] ;
   wire \ram[78][12] ;
   wire \ram[78][11] ;
   wire \ram[78][10] ;
   wire \ram[78][9] ;
   wire \ram[78][8] ;
   wire \ram[78][7] ;
   wire \ram[78][6] ;
   wire \ram[78][5] ;
   wire \ram[78][4] ;
   wire \ram[78][3] ;
   wire \ram[78][2] ;
   wire \ram[78][1] ;
   wire \ram[78][0] ;
   wire \ram[77][15] ;
   wire \ram[77][14] ;
   wire \ram[77][13] ;
   wire \ram[77][12] ;
   wire \ram[77][11] ;
   wire \ram[77][10] ;
   wire \ram[77][9] ;
   wire \ram[77][8] ;
   wire \ram[77][7] ;
   wire \ram[77][6] ;
   wire \ram[77][5] ;
   wire \ram[77][4] ;
   wire \ram[77][3] ;
   wire \ram[77][2] ;
   wire \ram[77][1] ;
   wire \ram[77][0] ;
   wire \ram[76][15] ;
   wire \ram[76][14] ;
   wire \ram[76][13] ;
   wire \ram[76][12] ;
   wire \ram[76][11] ;
   wire \ram[76][10] ;
   wire \ram[76][9] ;
   wire \ram[76][8] ;
   wire \ram[76][7] ;
   wire \ram[76][6] ;
   wire \ram[76][5] ;
   wire \ram[76][4] ;
   wire \ram[76][3] ;
   wire \ram[76][2] ;
   wire \ram[76][1] ;
   wire \ram[76][0] ;
   wire \ram[75][15] ;
   wire \ram[75][14] ;
   wire \ram[75][13] ;
   wire \ram[75][12] ;
   wire \ram[75][11] ;
   wire \ram[75][10] ;
   wire \ram[75][9] ;
   wire \ram[75][8] ;
   wire \ram[75][7] ;
   wire \ram[75][6] ;
   wire \ram[75][5] ;
   wire \ram[75][4] ;
   wire \ram[75][3] ;
   wire \ram[75][2] ;
   wire \ram[75][1] ;
   wire \ram[75][0] ;
   wire \ram[74][15] ;
   wire \ram[74][14] ;
   wire \ram[74][13] ;
   wire \ram[74][12] ;
   wire \ram[74][11] ;
   wire \ram[74][10] ;
   wire \ram[74][9] ;
   wire \ram[74][8] ;
   wire \ram[74][7] ;
   wire \ram[74][6] ;
   wire \ram[74][5] ;
   wire \ram[74][4] ;
   wire \ram[74][3] ;
   wire \ram[74][2] ;
   wire \ram[74][1] ;
   wire \ram[74][0] ;
   wire \ram[73][15] ;
   wire \ram[73][14] ;
   wire \ram[73][13] ;
   wire \ram[73][12] ;
   wire \ram[73][11] ;
   wire \ram[73][10] ;
   wire \ram[73][9] ;
   wire \ram[73][8] ;
   wire \ram[73][7] ;
   wire \ram[73][6] ;
   wire \ram[73][5] ;
   wire \ram[73][4] ;
   wire \ram[73][3] ;
   wire \ram[73][2] ;
   wire \ram[73][1] ;
   wire \ram[73][0] ;
   wire \ram[72][15] ;
   wire \ram[72][14] ;
   wire \ram[72][13] ;
   wire \ram[72][12] ;
   wire \ram[72][11] ;
   wire \ram[72][10] ;
   wire \ram[72][9] ;
   wire \ram[72][8] ;
   wire \ram[72][7] ;
   wire \ram[72][6] ;
   wire \ram[72][5] ;
   wire \ram[72][4] ;
   wire \ram[72][3] ;
   wire \ram[72][2] ;
   wire \ram[72][1] ;
   wire \ram[72][0] ;
   wire \ram[71][15] ;
   wire \ram[71][14] ;
   wire \ram[71][13] ;
   wire \ram[71][12] ;
   wire \ram[71][11] ;
   wire \ram[71][10] ;
   wire \ram[71][9] ;
   wire \ram[71][8] ;
   wire \ram[71][7] ;
   wire \ram[71][6] ;
   wire \ram[71][5] ;
   wire \ram[71][4] ;
   wire \ram[71][3] ;
   wire \ram[71][2] ;
   wire \ram[71][1] ;
   wire \ram[71][0] ;
   wire \ram[70][15] ;
   wire \ram[70][14] ;
   wire \ram[70][13] ;
   wire \ram[70][12] ;
   wire \ram[70][11] ;
   wire \ram[70][10] ;
   wire \ram[70][9] ;
   wire \ram[70][8] ;
   wire \ram[70][7] ;
   wire \ram[70][6] ;
   wire \ram[70][5] ;
   wire \ram[70][4] ;
   wire \ram[70][3] ;
   wire \ram[70][2] ;
   wire \ram[70][1] ;
   wire \ram[70][0] ;
   wire \ram[69][15] ;
   wire \ram[69][14] ;
   wire \ram[69][13] ;
   wire \ram[69][12] ;
   wire \ram[69][11] ;
   wire \ram[69][10] ;
   wire \ram[69][9] ;
   wire \ram[69][8] ;
   wire \ram[69][7] ;
   wire \ram[69][6] ;
   wire \ram[69][5] ;
   wire \ram[69][4] ;
   wire \ram[69][3] ;
   wire \ram[69][2] ;
   wire \ram[69][1] ;
   wire \ram[69][0] ;
   wire \ram[68][15] ;
   wire \ram[68][14] ;
   wire \ram[68][13] ;
   wire \ram[68][12] ;
   wire \ram[68][11] ;
   wire \ram[68][10] ;
   wire \ram[68][9] ;
   wire \ram[68][8] ;
   wire \ram[68][7] ;
   wire \ram[68][6] ;
   wire \ram[68][5] ;
   wire \ram[68][4] ;
   wire \ram[68][3] ;
   wire \ram[68][2] ;
   wire \ram[68][1] ;
   wire \ram[68][0] ;
   wire \ram[67][15] ;
   wire \ram[67][14] ;
   wire \ram[67][13] ;
   wire \ram[67][12] ;
   wire \ram[67][11] ;
   wire \ram[67][10] ;
   wire \ram[67][9] ;
   wire \ram[67][8] ;
   wire \ram[67][7] ;
   wire \ram[67][6] ;
   wire \ram[67][5] ;
   wire \ram[67][4] ;
   wire \ram[67][3] ;
   wire \ram[67][2] ;
   wire \ram[67][1] ;
   wire \ram[67][0] ;
   wire \ram[66][15] ;
   wire \ram[66][14] ;
   wire \ram[66][13] ;
   wire \ram[66][12] ;
   wire \ram[66][11] ;
   wire \ram[66][10] ;
   wire \ram[66][9] ;
   wire \ram[66][8] ;
   wire \ram[66][7] ;
   wire \ram[66][6] ;
   wire \ram[66][5] ;
   wire \ram[66][4] ;
   wire \ram[66][3] ;
   wire \ram[66][2] ;
   wire \ram[66][1] ;
   wire \ram[66][0] ;
   wire \ram[65][15] ;
   wire \ram[65][14] ;
   wire \ram[65][13] ;
   wire \ram[65][12] ;
   wire \ram[65][11] ;
   wire \ram[65][10] ;
   wire \ram[65][9] ;
   wire \ram[65][8] ;
   wire \ram[65][7] ;
   wire \ram[65][6] ;
   wire \ram[65][5] ;
   wire \ram[65][4] ;
   wire \ram[65][3] ;
   wire \ram[65][2] ;
   wire \ram[65][1] ;
   wire \ram[65][0] ;
   wire \ram[64][15] ;
   wire \ram[64][14] ;
   wire \ram[64][13] ;
   wire \ram[64][12] ;
   wire \ram[64][11] ;
   wire \ram[64][10] ;
   wire \ram[64][9] ;
   wire \ram[64][8] ;
   wire \ram[64][7] ;
   wire \ram[64][6] ;
   wire \ram[64][5] ;
   wire \ram[64][4] ;
   wire \ram[64][3] ;
   wire \ram[64][2] ;
   wire \ram[64][1] ;
   wire \ram[64][0] ;
   wire \ram[63][15] ;
   wire \ram[63][14] ;
   wire \ram[63][13] ;
   wire \ram[63][12] ;
   wire \ram[63][11] ;
   wire \ram[63][10] ;
   wire \ram[63][9] ;
   wire \ram[63][8] ;
   wire \ram[63][7] ;
   wire \ram[63][6] ;
   wire \ram[63][5] ;
   wire \ram[63][4] ;
   wire \ram[63][3] ;
   wire \ram[63][2] ;
   wire \ram[63][1] ;
   wire \ram[63][0] ;
   wire \ram[62][15] ;
   wire \ram[62][14] ;
   wire \ram[62][13] ;
   wire \ram[62][12] ;
   wire \ram[62][11] ;
   wire \ram[62][10] ;
   wire \ram[62][9] ;
   wire \ram[62][8] ;
   wire \ram[62][7] ;
   wire \ram[62][6] ;
   wire \ram[62][5] ;
   wire \ram[62][4] ;
   wire \ram[62][3] ;
   wire \ram[62][2] ;
   wire \ram[62][1] ;
   wire \ram[62][0] ;
   wire \ram[61][15] ;
   wire \ram[61][14] ;
   wire \ram[61][13] ;
   wire \ram[61][12] ;
   wire \ram[61][11] ;
   wire \ram[61][10] ;
   wire \ram[61][9] ;
   wire \ram[61][8] ;
   wire \ram[61][7] ;
   wire \ram[61][6] ;
   wire \ram[61][5] ;
   wire \ram[61][4] ;
   wire \ram[61][3] ;
   wire \ram[61][2] ;
   wire \ram[61][1] ;
   wire \ram[61][0] ;
   wire \ram[60][15] ;
   wire \ram[60][14] ;
   wire \ram[60][13] ;
   wire \ram[60][12] ;
   wire \ram[60][11] ;
   wire \ram[60][10] ;
   wire \ram[60][9] ;
   wire \ram[60][8] ;
   wire \ram[60][7] ;
   wire \ram[60][6] ;
   wire \ram[60][5] ;
   wire \ram[60][4] ;
   wire \ram[60][3] ;
   wire \ram[60][2] ;
   wire \ram[60][1] ;
   wire \ram[60][0] ;
   wire \ram[59][15] ;
   wire \ram[59][14] ;
   wire \ram[59][13] ;
   wire \ram[59][12] ;
   wire \ram[59][11] ;
   wire \ram[59][10] ;
   wire \ram[59][9] ;
   wire \ram[59][8] ;
   wire \ram[59][7] ;
   wire \ram[59][6] ;
   wire \ram[59][5] ;
   wire \ram[59][4] ;
   wire \ram[59][3] ;
   wire \ram[59][2] ;
   wire \ram[59][1] ;
   wire \ram[59][0] ;
   wire \ram[58][15] ;
   wire \ram[58][14] ;
   wire \ram[58][13] ;
   wire \ram[58][12] ;
   wire \ram[58][11] ;
   wire \ram[58][10] ;
   wire \ram[58][9] ;
   wire \ram[58][8] ;
   wire \ram[58][7] ;
   wire \ram[58][6] ;
   wire \ram[58][5] ;
   wire \ram[58][4] ;
   wire \ram[58][3] ;
   wire \ram[58][2] ;
   wire \ram[58][1] ;
   wire \ram[58][0] ;
   wire \ram[57][15] ;
   wire \ram[57][14] ;
   wire \ram[57][13] ;
   wire \ram[57][12] ;
   wire \ram[57][11] ;
   wire \ram[57][10] ;
   wire \ram[57][9] ;
   wire \ram[57][8] ;
   wire \ram[57][7] ;
   wire \ram[57][6] ;
   wire \ram[57][5] ;
   wire \ram[57][4] ;
   wire \ram[57][3] ;
   wire \ram[57][2] ;
   wire \ram[57][1] ;
   wire \ram[57][0] ;
   wire \ram[56][15] ;
   wire \ram[56][14] ;
   wire \ram[56][13] ;
   wire \ram[56][12] ;
   wire \ram[56][11] ;
   wire \ram[56][10] ;
   wire \ram[56][9] ;
   wire \ram[56][8] ;
   wire \ram[56][7] ;
   wire \ram[56][6] ;
   wire \ram[56][5] ;
   wire \ram[56][4] ;
   wire \ram[56][3] ;
   wire \ram[56][2] ;
   wire \ram[56][1] ;
   wire \ram[56][0] ;
   wire \ram[55][15] ;
   wire \ram[55][14] ;
   wire \ram[55][13] ;
   wire \ram[55][12] ;
   wire \ram[55][11] ;
   wire \ram[55][10] ;
   wire \ram[55][9] ;
   wire \ram[55][8] ;
   wire \ram[55][7] ;
   wire \ram[55][6] ;
   wire \ram[55][5] ;
   wire \ram[55][4] ;
   wire \ram[55][3] ;
   wire \ram[55][2] ;
   wire \ram[55][1] ;
   wire \ram[55][0] ;
   wire \ram[54][15] ;
   wire \ram[54][14] ;
   wire \ram[54][13] ;
   wire \ram[54][12] ;
   wire \ram[54][11] ;
   wire \ram[54][10] ;
   wire \ram[54][9] ;
   wire \ram[54][8] ;
   wire \ram[54][7] ;
   wire \ram[54][6] ;
   wire \ram[54][5] ;
   wire \ram[54][4] ;
   wire \ram[54][3] ;
   wire \ram[54][2] ;
   wire \ram[54][1] ;
   wire \ram[54][0] ;
   wire \ram[53][15] ;
   wire \ram[53][14] ;
   wire \ram[53][13] ;
   wire \ram[53][12] ;
   wire \ram[53][11] ;
   wire \ram[53][10] ;
   wire \ram[53][9] ;
   wire \ram[53][8] ;
   wire \ram[53][7] ;
   wire \ram[53][6] ;
   wire \ram[53][5] ;
   wire \ram[53][4] ;
   wire \ram[53][3] ;
   wire \ram[53][2] ;
   wire \ram[53][1] ;
   wire \ram[53][0] ;
   wire \ram[52][15] ;
   wire \ram[52][14] ;
   wire \ram[52][13] ;
   wire \ram[52][12] ;
   wire \ram[52][11] ;
   wire \ram[52][10] ;
   wire \ram[52][9] ;
   wire \ram[52][8] ;
   wire \ram[52][7] ;
   wire \ram[52][6] ;
   wire \ram[52][5] ;
   wire \ram[52][4] ;
   wire \ram[52][3] ;
   wire \ram[52][2] ;
   wire \ram[52][1] ;
   wire \ram[52][0] ;
   wire \ram[51][15] ;
   wire \ram[51][14] ;
   wire \ram[51][13] ;
   wire \ram[51][12] ;
   wire \ram[51][11] ;
   wire \ram[51][10] ;
   wire \ram[51][9] ;
   wire \ram[51][8] ;
   wire \ram[51][7] ;
   wire \ram[51][6] ;
   wire \ram[51][5] ;
   wire \ram[51][4] ;
   wire \ram[51][3] ;
   wire \ram[51][2] ;
   wire \ram[51][1] ;
   wire \ram[51][0] ;
   wire \ram[50][15] ;
   wire \ram[50][14] ;
   wire \ram[50][13] ;
   wire \ram[50][12] ;
   wire \ram[50][11] ;
   wire \ram[50][10] ;
   wire \ram[50][9] ;
   wire \ram[50][8] ;
   wire \ram[50][7] ;
   wire \ram[50][6] ;
   wire \ram[50][5] ;
   wire \ram[50][4] ;
   wire \ram[50][3] ;
   wire \ram[50][2] ;
   wire \ram[50][1] ;
   wire \ram[50][0] ;
   wire \ram[49][15] ;
   wire \ram[49][14] ;
   wire \ram[49][13] ;
   wire \ram[49][12] ;
   wire \ram[49][11] ;
   wire \ram[49][10] ;
   wire \ram[49][9] ;
   wire \ram[49][8] ;
   wire \ram[49][7] ;
   wire \ram[49][6] ;
   wire \ram[49][5] ;
   wire \ram[49][4] ;
   wire \ram[49][3] ;
   wire \ram[49][2] ;
   wire \ram[49][1] ;
   wire \ram[49][0] ;
   wire \ram[48][15] ;
   wire \ram[48][14] ;
   wire \ram[48][13] ;
   wire \ram[48][12] ;
   wire \ram[48][11] ;
   wire \ram[48][10] ;
   wire \ram[48][9] ;
   wire \ram[48][8] ;
   wire \ram[48][7] ;
   wire \ram[48][6] ;
   wire \ram[48][5] ;
   wire \ram[48][4] ;
   wire \ram[48][3] ;
   wire \ram[48][2] ;
   wire \ram[48][1] ;
   wire \ram[48][0] ;
   wire \ram[47][15] ;
   wire \ram[47][14] ;
   wire \ram[47][13] ;
   wire \ram[47][12] ;
   wire \ram[47][11] ;
   wire \ram[47][10] ;
   wire \ram[47][9] ;
   wire \ram[47][8] ;
   wire \ram[47][7] ;
   wire \ram[47][6] ;
   wire \ram[47][5] ;
   wire \ram[47][4] ;
   wire \ram[47][3] ;
   wire \ram[47][2] ;
   wire \ram[47][1] ;
   wire \ram[47][0] ;
   wire \ram[46][15] ;
   wire \ram[46][14] ;
   wire \ram[46][13] ;
   wire \ram[46][12] ;
   wire \ram[46][11] ;
   wire \ram[46][10] ;
   wire \ram[46][9] ;
   wire \ram[46][8] ;
   wire \ram[46][7] ;
   wire \ram[46][6] ;
   wire \ram[46][5] ;
   wire \ram[46][4] ;
   wire \ram[46][3] ;
   wire \ram[46][2] ;
   wire \ram[46][1] ;
   wire \ram[46][0] ;
   wire \ram[45][15] ;
   wire \ram[45][14] ;
   wire \ram[45][13] ;
   wire \ram[45][12] ;
   wire \ram[45][11] ;
   wire \ram[45][10] ;
   wire \ram[45][9] ;
   wire \ram[45][8] ;
   wire \ram[45][7] ;
   wire \ram[45][6] ;
   wire \ram[45][5] ;
   wire \ram[45][4] ;
   wire \ram[45][3] ;
   wire \ram[45][2] ;
   wire \ram[45][1] ;
   wire \ram[45][0] ;
   wire \ram[44][15] ;
   wire \ram[44][14] ;
   wire \ram[44][13] ;
   wire \ram[44][12] ;
   wire \ram[44][11] ;
   wire \ram[44][10] ;
   wire \ram[44][9] ;
   wire \ram[44][8] ;
   wire \ram[44][7] ;
   wire \ram[44][6] ;
   wire \ram[44][5] ;
   wire \ram[44][4] ;
   wire \ram[44][3] ;
   wire \ram[44][2] ;
   wire \ram[44][1] ;
   wire \ram[44][0] ;
   wire \ram[43][15] ;
   wire \ram[43][14] ;
   wire \ram[43][13] ;
   wire \ram[43][12] ;
   wire \ram[43][11] ;
   wire \ram[43][10] ;
   wire \ram[43][9] ;
   wire \ram[43][8] ;
   wire \ram[43][7] ;
   wire \ram[43][6] ;
   wire \ram[43][5] ;
   wire \ram[43][4] ;
   wire \ram[43][3] ;
   wire \ram[43][2] ;
   wire \ram[43][1] ;
   wire \ram[43][0] ;
   wire \ram[42][15] ;
   wire \ram[42][14] ;
   wire \ram[42][13] ;
   wire \ram[42][12] ;
   wire \ram[42][11] ;
   wire \ram[42][10] ;
   wire \ram[42][9] ;
   wire \ram[42][8] ;
   wire \ram[42][7] ;
   wire \ram[42][6] ;
   wire \ram[42][5] ;
   wire \ram[42][4] ;
   wire \ram[42][3] ;
   wire \ram[42][2] ;
   wire \ram[42][1] ;
   wire \ram[42][0] ;
   wire \ram[41][15] ;
   wire \ram[41][14] ;
   wire \ram[41][13] ;
   wire \ram[41][12] ;
   wire \ram[41][11] ;
   wire \ram[41][10] ;
   wire \ram[41][9] ;
   wire \ram[41][8] ;
   wire \ram[41][7] ;
   wire \ram[41][6] ;
   wire \ram[41][5] ;
   wire \ram[41][4] ;
   wire \ram[41][3] ;
   wire \ram[41][2] ;
   wire \ram[41][1] ;
   wire \ram[41][0] ;
   wire \ram[40][15] ;
   wire \ram[40][14] ;
   wire \ram[40][13] ;
   wire \ram[40][12] ;
   wire \ram[40][11] ;
   wire \ram[40][10] ;
   wire \ram[40][9] ;
   wire \ram[40][8] ;
   wire \ram[40][7] ;
   wire \ram[40][6] ;
   wire \ram[40][5] ;
   wire \ram[40][4] ;
   wire \ram[40][3] ;
   wire \ram[40][2] ;
   wire \ram[40][1] ;
   wire \ram[40][0] ;
   wire \ram[39][15] ;
   wire \ram[39][14] ;
   wire \ram[39][13] ;
   wire \ram[39][12] ;
   wire \ram[39][11] ;
   wire \ram[39][10] ;
   wire \ram[39][9] ;
   wire \ram[39][8] ;
   wire \ram[39][7] ;
   wire \ram[39][6] ;
   wire \ram[39][5] ;
   wire \ram[39][4] ;
   wire \ram[39][3] ;
   wire \ram[39][2] ;
   wire \ram[39][1] ;
   wire \ram[39][0] ;
   wire \ram[38][15] ;
   wire \ram[38][14] ;
   wire \ram[38][13] ;
   wire \ram[38][12] ;
   wire \ram[38][11] ;
   wire \ram[38][10] ;
   wire \ram[38][9] ;
   wire \ram[38][8] ;
   wire \ram[38][7] ;
   wire \ram[38][6] ;
   wire \ram[38][5] ;
   wire \ram[38][4] ;
   wire \ram[38][3] ;
   wire \ram[38][2] ;
   wire \ram[38][1] ;
   wire \ram[38][0] ;
   wire \ram[37][15] ;
   wire \ram[37][14] ;
   wire \ram[37][13] ;
   wire \ram[37][12] ;
   wire \ram[37][11] ;
   wire \ram[37][10] ;
   wire \ram[37][9] ;
   wire \ram[37][8] ;
   wire \ram[37][7] ;
   wire \ram[37][6] ;
   wire \ram[37][5] ;
   wire \ram[37][4] ;
   wire \ram[37][3] ;
   wire \ram[37][2] ;
   wire \ram[37][1] ;
   wire \ram[37][0] ;
   wire \ram[36][15] ;
   wire \ram[36][14] ;
   wire \ram[36][13] ;
   wire \ram[36][12] ;
   wire \ram[36][11] ;
   wire \ram[36][10] ;
   wire \ram[36][9] ;
   wire \ram[36][8] ;
   wire \ram[36][7] ;
   wire \ram[36][6] ;
   wire \ram[36][5] ;
   wire \ram[36][4] ;
   wire \ram[36][3] ;
   wire \ram[36][2] ;
   wire \ram[36][1] ;
   wire \ram[36][0] ;
   wire \ram[35][15] ;
   wire \ram[35][14] ;
   wire \ram[35][13] ;
   wire \ram[35][12] ;
   wire \ram[35][11] ;
   wire \ram[35][10] ;
   wire \ram[35][9] ;
   wire \ram[35][8] ;
   wire \ram[35][7] ;
   wire \ram[35][6] ;
   wire \ram[35][5] ;
   wire \ram[35][4] ;
   wire \ram[35][3] ;
   wire \ram[35][2] ;
   wire \ram[35][1] ;
   wire \ram[35][0] ;
   wire \ram[34][15] ;
   wire \ram[34][14] ;
   wire \ram[34][13] ;
   wire \ram[34][12] ;
   wire \ram[34][11] ;
   wire \ram[34][10] ;
   wire \ram[34][9] ;
   wire \ram[34][8] ;
   wire \ram[34][7] ;
   wire \ram[34][6] ;
   wire \ram[34][5] ;
   wire \ram[34][4] ;
   wire \ram[34][3] ;
   wire \ram[34][2] ;
   wire \ram[34][1] ;
   wire \ram[34][0] ;
   wire \ram[33][15] ;
   wire \ram[33][14] ;
   wire \ram[33][13] ;
   wire \ram[33][12] ;
   wire \ram[33][11] ;
   wire \ram[33][10] ;
   wire \ram[33][9] ;
   wire \ram[33][8] ;
   wire \ram[33][7] ;
   wire \ram[33][6] ;
   wire \ram[33][5] ;
   wire \ram[33][4] ;
   wire \ram[33][3] ;
   wire \ram[33][2] ;
   wire \ram[33][1] ;
   wire \ram[33][0] ;
   wire \ram[32][15] ;
   wire \ram[32][14] ;
   wire \ram[32][13] ;
   wire \ram[32][12] ;
   wire \ram[32][11] ;
   wire \ram[32][10] ;
   wire \ram[32][9] ;
   wire \ram[32][8] ;
   wire \ram[32][7] ;
   wire \ram[32][6] ;
   wire \ram[32][5] ;
   wire \ram[32][4] ;
   wire \ram[32][3] ;
   wire \ram[32][2] ;
   wire \ram[32][1] ;
   wire \ram[32][0] ;
   wire \ram[31][15] ;
   wire \ram[31][14] ;
   wire \ram[31][13] ;
   wire \ram[31][12] ;
   wire \ram[31][11] ;
   wire \ram[31][10] ;
   wire \ram[31][9] ;
   wire \ram[31][8] ;
   wire \ram[31][7] ;
   wire \ram[31][6] ;
   wire \ram[31][5] ;
   wire \ram[31][4] ;
   wire \ram[31][3] ;
   wire \ram[31][2] ;
   wire \ram[31][1] ;
   wire \ram[31][0] ;
   wire \ram[30][15] ;
   wire \ram[30][14] ;
   wire \ram[30][13] ;
   wire \ram[30][12] ;
   wire \ram[30][11] ;
   wire \ram[30][10] ;
   wire \ram[30][9] ;
   wire \ram[30][8] ;
   wire \ram[30][7] ;
   wire \ram[30][6] ;
   wire \ram[30][5] ;
   wire \ram[30][4] ;
   wire \ram[30][3] ;
   wire \ram[30][2] ;
   wire \ram[30][1] ;
   wire \ram[30][0] ;
   wire \ram[29][15] ;
   wire \ram[29][14] ;
   wire \ram[29][13] ;
   wire \ram[29][12] ;
   wire \ram[29][11] ;
   wire \ram[29][10] ;
   wire \ram[29][9] ;
   wire \ram[29][8] ;
   wire \ram[29][7] ;
   wire \ram[29][6] ;
   wire \ram[29][5] ;
   wire \ram[29][4] ;
   wire \ram[29][3] ;
   wire \ram[29][2] ;
   wire \ram[29][1] ;
   wire \ram[29][0] ;
   wire \ram[28][15] ;
   wire \ram[28][14] ;
   wire \ram[28][13] ;
   wire \ram[28][12] ;
   wire \ram[28][11] ;
   wire \ram[28][10] ;
   wire \ram[28][9] ;
   wire \ram[28][8] ;
   wire \ram[28][7] ;
   wire \ram[28][6] ;
   wire \ram[28][5] ;
   wire \ram[28][4] ;
   wire \ram[28][3] ;
   wire \ram[28][2] ;
   wire \ram[28][1] ;
   wire \ram[28][0] ;
   wire \ram[27][15] ;
   wire \ram[27][14] ;
   wire \ram[27][13] ;
   wire \ram[27][12] ;
   wire \ram[27][11] ;
   wire \ram[27][10] ;
   wire \ram[27][9] ;
   wire \ram[27][8] ;
   wire \ram[27][7] ;
   wire \ram[27][6] ;
   wire \ram[27][5] ;
   wire \ram[27][4] ;
   wire \ram[27][3] ;
   wire \ram[27][2] ;
   wire \ram[27][1] ;
   wire \ram[27][0] ;
   wire \ram[26][15] ;
   wire \ram[26][14] ;
   wire \ram[26][13] ;
   wire \ram[26][12] ;
   wire \ram[26][11] ;
   wire \ram[26][10] ;
   wire \ram[26][9] ;
   wire \ram[26][8] ;
   wire \ram[26][7] ;
   wire \ram[26][6] ;
   wire \ram[26][5] ;
   wire \ram[26][4] ;
   wire \ram[26][3] ;
   wire \ram[26][2] ;
   wire \ram[26][1] ;
   wire \ram[26][0] ;
   wire \ram[25][15] ;
   wire \ram[25][14] ;
   wire \ram[25][13] ;
   wire \ram[25][12] ;
   wire \ram[25][11] ;
   wire \ram[25][10] ;
   wire \ram[25][9] ;
   wire \ram[25][8] ;
   wire \ram[25][7] ;
   wire \ram[25][6] ;
   wire \ram[25][5] ;
   wire \ram[25][4] ;
   wire \ram[25][3] ;
   wire \ram[25][2] ;
   wire \ram[25][1] ;
   wire \ram[25][0] ;
   wire \ram[24][15] ;
   wire \ram[24][14] ;
   wire \ram[24][13] ;
   wire \ram[24][12] ;
   wire \ram[24][11] ;
   wire \ram[24][10] ;
   wire \ram[24][9] ;
   wire \ram[24][8] ;
   wire \ram[24][7] ;
   wire \ram[24][6] ;
   wire \ram[24][5] ;
   wire \ram[24][4] ;
   wire \ram[24][3] ;
   wire \ram[24][2] ;
   wire \ram[24][1] ;
   wire \ram[24][0] ;
   wire \ram[23][15] ;
   wire \ram[23][14] ;
   wire \ram[23][13] ;
   wire \ram[23][12] ;
   wire \ram[23][11] ;
   wire \ram[23][10] ;
   wire \ram[23][9] ;
   wire \ram[23][8] ;
   wire \ram[23][7] ;
   wire \ram[23][6] ;
   wire \ram[23][5] ;
   wire \ram[23][4] ;
   wire \ram[23][3] ;
   wire \ram[23][2] ;
   wire \ram[23][1] ;
   wire \ram[23][0] ;
   wire \ram[22][15] ;
   wire \ram[22][14] ;
   wire \ram[22][13] ;
   wire \ram[22][12] ;
   wire \ram[22][11] ;
   wire \ram[22][10] ;
   wire \ram[22][9] ;
   wire \ram[22][8] ;
   wire \ram[22][7] ;
   wire \ram[22][6] ;
   wire \ram[22][5] ;
   wire \ram[22][4] ;
   wire \ram[22][3] ;
   wire \ram[22][2] ;
   wire \ram[22][1] ;
   wire \ram[22][0] ;
   wire \ram[21][15] ;
   wire \ram[21][14] ;
   wire \ram[21][13] ;
   wire \ram[21][12] ;
   wire \ram[21][11] ;
   wire \ram[21][10] ;
   wire \ram[21][9] ;
   wire \ram[21][8] ;
   wire \ram[21][7] ;
   wire \ram[21][6] ;
   wire \ram[21][5] ;
   wire \ram[21][4] ;
   wire \ram[21][3] ;
   wire \ram[21][2] ;
   wire \ram[21][1] ;
   wire \ram[21][0] ;
   wire \ram[20][15] ;
   wire \ram[20][14] ;
   wire \ram[20][13] ;
   wire \ram[20][12] ;
   wire \ram[20][11] ;
   wire \ram[20][10] ;
   wire \ram[20][9] ;
   wire \ram[20][8] ;
   wire \ram[20][7] ;
   wire \ram[20][6] ;
   wire \ram[20][5] ;
   wire \ram[20][4] ;
   wire \ram[20][3] ;
   wire \ram[20][2] ;
   wire \ram[20][1] ;
   wire \ram[20][0] ;
   wire \ram[19][15] ;
   wire \ram[19][14] ;
   wire \ram[19][13] ;
   wire \ram[19][12] ;
   wire \ram[19][11] ;
   wire \ram[19][10] ;
   wire \ram[19][9] ;
   wire \ram[19][8] ;
   wire \ram[19][7] ;
   wire \ram[19][6] ;
   wire \ram[19][5] ;
   wire \ram[19][4] ;
   wire \ram[19][3] ;
   wire \ram[19][2] ;
   wire \ram[19][1] ;
   wire \ram[19][0] ;
   wire \ram[18][15] ;
   wire \ram[18][14] ;
   wire \ram[18][13] ;
   wire \ram[18][12] ;
   wire \ram[18][11] ;
   wire \ram[18][10] ;
   wire \ram[18][9] ;
   wire \ram[18][8] ;
   wire \ram[18][7] ;
   wire \ram[18][6] ;
   wire \ram[18][5] ;
   wire \ram[18][4] ;
   wire \ram[18][3] ;
   wire \ram[18][2] ;
   wire \ram[18][1] ;
   wire \ram[18][0] ;
   wire \ram[17][15] ;
   wire \ram[17][14] ;
   wire \ram[17][13] ;
   wire \ram[17][12] ;
   wire \ram[17][11] ;
   wire \ram[17][10] ;
   wire \ram[17][9] ;
   wire \ram[17][8] ;
   wire \ram[17][7] ;
   wire \ram[17][6] ;
   wire \ram[17][5] ;
   wire \ram[17][4] ;
   wire \ram[17][3] ;
   wire \ram[17][2] ;
   wire \ram[17][1] ;
   wire \ram[17][0] ;
   wire \ram[16][15] ;
   wire \ram[16][14] ;
   wire \ram[16][13] ;
   wire \ram[16][12] ;
   wire \ram[16][11] ;
   wire \ram[16][10] ;
   wire \ram[16][9] ;
   wire \ram[16][8] ;
   wire \ram[16][7] ;
   wire \ram[16][6] ;
   wire \ram[16][5] ;
   wire \ram[16][4] ;
   wire \ram[16][3] ;
   wire \ram[16][2] ;
   wire \ram[16][1] ;
   wire \ram[16][0] ;
   wire \ram[15][15] ;
   wire \ram[15][14] ;
   wire \ram[15][13] ;
   wire \ram[15][12] ;
   wire \ram[15][11] ;
   wire \ram[15][10] ;
   wire \ram[15][9] ;
   wire \ram[15][8] ;
   wire \ram[15][7] ;
   wire \ram[15][6] ;
   wire \ram[15][5] ;
   wire \ram[15][4] ;
   wire \ram[15][3] ;
   wire \ram[15][2] ;
   wire \ram[15][1] ;
   wire \ram[15][0] ;
   wire \ram[14][15] ;
   wire \ram[14][14] ;
   wire \ram[14][13] ;
   wire \ram[14][12] ;
   wire \ram[14][11] ;
   wire \ram[14][10] ;
   wire \ram[14][9] ;
   wire \ram[14][8] ;
   wire \ram[14][7] ;
   wire \ram[14][6] ;
   wire \ram[14][5] ;
   wire \ram[14][4] ;
   wire \ram[14][3] ;
   wire \ram[14][2] ;
   wire \ram[14][1] ;
   wire \ram[14][0] ;
   wire \ram[13][15] ;
   wire \ram[13][14] ;
   wire \ram[13][13] ;
   wire \ram[13][12] ;
   wire \ram[13][11] ;
   wire \ram[13][10] ;
   wire \ram[13][9] ;
   wire \ram[13][8] ;
   wire \ram[13][7] ;
   wire \ram[13][6] ;
   wire \ram[13][5] ;
   wire \ram[13][4] ;
   wire \ram[13][3] ;
   wire \ram[13][2] ;
   wire \ram[13][1] ;
   wire \ram[13][0] ;
   wire \ram[12][15] ;
   wire \ram[12][14] ;
   wire \ram[12][13] ;
   wire \ram[12][12] ;
   wire \ram[12][11] ;
   wire \ram[12][10] ;
   wire \ram[12][9] ;
   wire \ram[12][8] ;
   wire \ram[12][7] ;
   wire \ram[12][6] ;
   wire \ram[12][5] ;
   wire \ram[12][4] ;
   wire \ram[12][3] ;
   wire \ram[12][2] ;
   wire \ram[12][1] ;
   wire \ram[12][0] ;
   wire \ram[11][15] ;
   wire \ram[11][14] ;
   wire \ram[11][13] ;
   wire \ram[11][12] ;
   wire \ram[11][11] ;
   wire \ram[11][10] ;
   wire \ram[11][9] ;
   wire \ram[11][8] ;
   wire \ram[11][7] ;
   wire \ram[11][6] ;
   wire \ram[11][5] ;
   wire \ram[11][4] ;
   wire \ram[11][3] ;
   wire \ram[11][2] ;
   wire \ram[11][1] ;
   wire \ram[11][0] ;
   wire \ram[10][15] ;
   wire \ram[10][14] ;
   wire \ram[10][13] ;
   wire \ram[10][12] ;
   wire \ram[10][11] ;
   wire \ram[10][10] ;
   wire \ram[10][9] ;
   wire \ram[10][8] ;
   wire \ram[10][7] ;
   wire \ram[10][6] ;
   wire \ram[10][5] ;
   wire \ram[10][4] ;
   wire \ram[10][3] ;
   wire \ram[10][2] ;
   wire \ram[10][1] ;
   wire \ram[10][0] ;
   wire \ram[9][15] ;
   wire \ram[9][14] ;
   wire \ram[9][13] ;
   wire \ram[9][12] ;
   wire \ram[9][11] ;
   wire \ram[9][10] ;
   wire \ram[9][9] ;
   wire \ram[9][8] ;
   wire \ram[9][7] ;
   wire \ram[9][6] ;
   wire \ram[9][5] ;
   wire \ram[9][4] ;
   wire \ram[9][3] ;
   wire \ram[9][2] ;
   wire \ram[9][1] ;
   wire \ram[9][0] ;
   wire \ram[8][15] ;
   wire \ram[8][14] ;
   wire \ram[8][13] ;
   wire \ram[8][12] ;
   wire \ram[8][11] ;
   wire \ram[8][10] ;
   wire \ram[8][9] ;
   wire \ram[8][8] ;
   wire \ram[8][7] ;
   wire \ram[8][6] ;
   wire \ram[8][5] ;
   wire \ram[8][4] ;
   wire \ram[8][3] ;
   wire \ram[8][2] ;
   wire \ram[8][1] ;
   wire \ram[8][0] ;
   wire \ram[7][15] ;
   wire \ram[7][14] ;
   wire \ram[7][13] ;
   wire \ram[7][12] ;
   wire \ram[7][11] ;
   wire \ram[7][10] ;
   wire \ram[7][9] ;
   wire \ram[7][8] ;
   wire \ram[7][7] ;
   wire \ram[7][6] ;
   wire \ram[7][5] ;
   wire \ram[7][4] ;
   wire \ram[7][3] ;
   wire \ram[7][2] ;
   wire \ram[7][1] ;
   wire \ram[7][0] ;
   wire \ram[6][15] ;
   wire \ram[6][14] ;
   wire \ram[6][13] ;
   wire \ram[6][12] ;
   wire \ram[6][11] ;
   wire \ram[6][10] ;
   wire \ram[6][9] ;
   wire \ram[6][8] ;
   wire \ram[6][7] ;
   wire \ram[6][6] ;
   wire \ram[6][5] ;
   wire \ram[6][4] ;
   wire \ram[6][3] ;
   wire \ram[6][2] ;
   wire \ram[6][1] ;
   wire \ram[6][0] ;
   wire \ram[5][15] ;
   wire \ram[5][14] ;
   wire \ram[5][13] ;
   wire \ram[5][12] ;
   wire \ram[5][11] ;
   wire \ram[5][10] ;
   wire \ram[5][9] ;
   wire \ram[5][8] ;
   wire \ram[5][7] ;
   wire \ram[5][6] ;
   wire \ram[5][5] ;
   wire \ram[5][4] ;
   wire \ram[5][3] ;
   wire \ram[5][2] ;
   wire \ram[5][1] ;
   wire \ram[5][0] ;
   wire \ram[4][15] ;
   wire \ram[4][14] ;
   wire \ram[4][13] ;
   wire \ram[4][12] ;
   wire \ram[4][11] ;
   wire \ram[4][10] ;
   wire \ram[4][9] ;
   wire \ram[4][8] ;
   wire \ram[4][7] ;
   wire \ram[4][6] ;
   wire \ram[4][5] ;
   wire \ram[4][4] ;
   wire \ram[4][3] ;
   wire \ram[4][2] ;
   wire \ram[4][1] ;
   wire \ram[4][0] ;
   wire \ram[3][15] ;
   wire \ram[3][14] ;
   wire \ram[3][13] ;
   wire \ram[3][12] ;
   wire \ram[3][11] ;
   wire \ram[3][10] ;
   wire \ram[3][9] ;
   wire \ram[3][8] ;
   wire \ram[3][7] ;
   wire \ram[3][6] ;
   wire \ram[3][5] ;
   wire \ram[3][4] ;
   wire \ram[3][3] ;
   wire \ram[3][2] ;
   wire \ram[3][1] ;
   wire \ram[3][0] ;
   wire \ram[2][15] ;
   wire \ram[2][14] ;
   wire \ram[2][13] ;
   wire \ram[2][12] ;
   wire \ram[2][11] ;
   wire \ram[2][10] ;
   wire \ram[2][9] ;
   wire \ram[2][8] ;
   wire \ram[2][7] ;
   wire \ram[2][6] ;
   wire \ram[2][5] ;
   wire \ram[2][4] ;
   wire \ram[2][3] ;
   wire \ram[2][2] ;
   wire \ram[2][1] ;
   wire \ram[2][0] ;
   wire \ram[1][15] ;
   wire \ram[1][14] ;
   wire \ram[1][13] ;
   wire \ram[1][12] ;
   wire \ram[1][11] ;
   wire \ram[1][10] ;
   wire \ram[1][9] ;
   wire \ram[1][8] ;
   wire \ram[1][7] ;
   wire \ram[1][6] ;
   wire \ram[1][5] ;
   wire \ram[1][4] ;
   wire \ram[1][3] ;
   wire \ram[1][2] ;
   wire \ram[1][1] ;
   wire \ram[1][0] ;
   wire \ram[0][15] ;
   wire \ram[0][14] ;
   wire \ram[0][13] ;
   wire \ram[0][12] ;
   wire \ram[0][11] ;
   wire \ram[0][10] ;
   wire \ram[0][9] ;
   wire \ram[0][8] ;
   wire \ram[0][7] ;
   wire \ram[0][6] ;
   wire \ram[0][5] ;
   wire \ram[0][4] ;
   wire \ram[0][3] ;
   wire \ram[0][2] ;
   wire \ram[0][1] ;
   wire \ram[0][0] ;
   wire N4126;
   wire N4127;
   wire N4128;
   wire N4129;
   wire N4130;
   wire N4131;
   wire N4132;
   wire N4133;
   wire N4134;
   wire N4135;
   wire N4136;
   wire N4137;
   wire N4138;
   wire N4139;
   wire N4140;
   wire N4141;
   wire n6;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n27;
   wire n30;
   wire n33;
   wire n36;
   wire n39;
   wire n42;
   wire n45;
   wire n48;
   wire n51;
   wire n54;
   wire n57;
   wire n60;
   wire n63;
   wire n66;
   wire n69;
   wire n71;
   wire n72;
   wire n74;
   wire n77;
   wire n79;
   wire n81;
   wire n83;
   wire n85;
   wire n87;
   wire n89;
   wire n91;
   wire n93;
   wire n95;
   wire n97;
   wire n99;
   wire n101;
   wire n103;
   wire n105;
   wire n106;
   wire n108;
   wire n111;
   wire n113;
   wire n115;
   wire n117;
   wire n119;
   wire n121;
   wire n123;
   wire n125;
   wire n127;
   wire n129;
   wire n131;
   wire n133;
   wire n135;
   wire n137;
   wire n139;
   wire n140;
   wire n142;
   wire n145;
   wire n147;
   wire n149;
   wire n151;
   wire n153;
   wire n155;
   wire n157;
   wire n159;
   wire n161;
   wire n163;
   wire n165;
   wire n167;
   wire n169;
   wire n171;
   wire n173;
   wire n174;
   wire n176;
   wire n179;
   wire n181;
   wire n183;
   wire n185;
   wire n187;
   wire n189;
   wire n191;
   wire n193;
   wire n195;
   wire n197;
   wire n199;
   wire n201;
   wire n203;
   wire n205;
   wire n207;
   wire n208;
   wire n210;
   wire n213;
   wire n215;
   wire n217;
   wire n219;
   wire n221;
   wire n223;
   wire n225;
   wire n227;
   wire n229;
   wire n231;
   wire n233;
   wire n235;
   wire n237;
   wire n239;
   wire n241;
   wire n243;
   wire n246;
   wire n248;
   wire n250;
   wire n252;
   wire n254;
   wire n256;
   wire n258;
   wire n260;
   wire n262;
   wire n264;
   wire n266;
   wire n268;
   wire n270;
   wire n272;
   wire n274;
   wire n276;
   wire n279;
   wire n281;
   wire n283;
   wire n285;
   wire n287;
   wire n289;
   wire n291;
   wire n293;
   wire n295;
   wire n297;
   wire n299;
   wire n301;
   wire n303;
   wire n305;
   wire n307;
   wire n309;
   wire n312;
   wire n314;
   wire n316;
   wire n318;
   wire n320;
   wire n322;
   wire n324;
   wire n326;
   wire n328;
   wire n330;
   wire n332;
   wire n334;
   wire n336;
   wire n338;
   wire n340;
   wire n341;
   wire n343;
   wire n346;
   wire n348;
   wire n350;
   wire n352;
   wire n354;
   wire n356;
   wire n358;
   wire n360;
   wire n362;
   wire n364;
   wire n366;
   wire n368;
   wire n370;
   wire n372;
   wire n374;
   wire n376;
   wire n379;
   wire n381;
   wire n383;
   wire n385;
   wire n387;
   wire n389;
   wire n391;
   wire n393;
   wire n395;
   wire n397;
   wire n399;
   wire n401;
   wire n403;
   wire n405;
   wire n407;
   wire n409;
   wire n412;
   wire n414;
   wire n416;
   wire n418;
   wire n420;
   wire n422;
   wire n424;
   wire n426;
   wire n428;
   wire n430;
   wire n432;
   wire n434;
   wire n436;
   wire n438;
   wire n440;
   wire n442;
   wire n445;
   wire n447;
   wire n449;
   wire n451;
   wire n453;
   wire n455;
   wire n457;
   wire n459;
   wire n461;
   wire n463;
   wire n465;
   wire n467;
   wire n469;
   wire n471;
   wire n473;
   wire n474;
   wire n476;
   wire n479;
   wire n481;
   wire n483;
   wire n485;
   wire n487;
   wire n489;
   wire n491;
   wire n493;
   wire n495;
   wire n497;
   wire n499;
   wire n501;
   wire n503;
   wire n505;
   wire n507;
   wire n509;
   wire n512;
   wire n514;
   wire n516;
   wire n518;
   wire n520;
   wire n522;
   wire n524;
   wire n526;
   wire n528;
   wire n530;
   wire n532;
   wire n534;
   wire n536;
   wire n538;
   wire n540;
   wire n542;
   wire n544;
   wire n545;
   wire n547;
   wire n548;
   wire n550;
   wire n551;
   wire n553;
   wire n554;
   wire n556;
   wire n557;
   wire n559;
   wire n561;
   wire n563;
   wire n565;
   wire n566;
   wire n568;
   wire n570;
   wire n572;
   wire n574;
   wire n575;
   wire n577;
   wire n579;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3297;
   wire n3298;
   wire n3299;
   wire n3300;
   wire n3301;
   wire n3302;
   wire n3303;
   wire n3304;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire n3330;
   wire n3331;
   wire n3332;
   wire n3333;
   wire n3334;
   wire n3335;
   wire n3336;
   wire n3337;
   wire n3338;
   wire n3339;
   wire n3340;
   wire n3341;
   wire n3342;
   wire n3343;
   wire n3344;
   wire n3345;
   wire n3346;
   wire n3347;
   wire n3348;
   wire n3349;
   wire n3350;
   wire n3351;
   wire n3352;
   wire n3353;
   wire n3354;
   wire n3355;
   wire n3356;
   wire n3357;
   wire n3358;
   wire n3359;
   wire n3360;
   wire n3361;
   wire n3362;
   wire n3363;
   wire n3364;
   wire n3365;
   wire n3366;
   wire n3367;
   wire n3368;
   wire n3369;
   wire n3370;
   wire n3371;
   wire n3372;
   wire n3373;
   wire n3374;
   wire n3375;
   wire n3376;
   wire n3377;
   wire n3378;
   wire n3379;
   wire n3380;
   wire n3381;
   wire n3382;
   wire n3383;
   wire n3384;
   wire n3385;
   wire n3386;
   wire n3387;
   wire n3388;
   wire n3389;
   wire n3390;
   wire n3391;
   wire n3392;
   wire n3393;
   wire n3394;
   wire n3395;
   wire n3396;
   wire n3397;
   wire n3398;
   wire n3399;
   wire n3400;
   wire n3401;
   wire n3402;
   wire n3403;
   wire n3404;
   wire n3405;
   wire n3406;
   wire n3407;
   wire n3408;
   wire n3409;
   wire n3410;
   wire n3411;
   wire n3412;
   wire n3413;
   wire n3414;
   wire n3415;
   wire n3416;
   wire n3417;
   wire n3418;
   wire n3419;
   wire n3420;
   wire n3421;
   wire n3422;
   wire n3423;
   wire n3424;
   wire n3425;
   wire n3426;
   wire n3427;
   wire n3428;
   wire n3429;
   wire n3430;
   wire n3431;
   wire n3432;
   wire n3433;
   wire n3434;
   wire n3435;
   wire n3436;
   wire n3437;
   wire n3438;
   wire n3439;
   wire n3440;
   wire n3441;
   wire n3442;
   wire n3443;
   wire n3444;
   wire n3445;
   wire n3446;
   wire n3447;
   wire n3448;
   wire n3449;
   wire n3450;
   wire n3451;
   wire n3452;
   wire n3453;
   wire n3454;
   wire n3455;
   wire n3456;
   wire n3457;
   wire n3458;
   wire n3459;
   wire n3460;
   wire n3461;
   wire n3462;
   wire n3463;
   wire n3464;
   wire n3465;
   wire n3466;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3475;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3485;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3589;
   wire n3590;
   wire n3591;
   wire n3592;
   wire n3593;
   wire n3594;
   wire n3595;
   wire n3596;
   wire n3597;
   wire n3598;
   wire n3599;
   wire n3600;
   wire n3601;
   wire n3602;
   wire n3603;
   wire n3604;
   wire n3605;
   wire n3606;
   wire n3607;
   wire n3608;
   wire n3609;
   wire n3610;
   wire n3611;
   wire n3612;
   wire n3613;
   wire n3614;
   wire n3615;
   wire n3616;
   wire n3617;
   wire n3618;
   wire n3619;
   wire n3620;
   wire n3621;
   wire n3622;
   wire n3623;
   wire n3624;
   wire n3625;
   wire n3626;
   wire n3627;
   wire n3628;
   wire n3629;
   wire n3630;
   wire n3631;
   wire n3632;
   wire n3633;
   wire n3634;
   wire n3635;
   wire n3636;
   wire n3637;
   wire n3638;
   wire n3639;
   wire n3640;
   wire n3641;
   wire n3642;
   wire n3643;
   wire n3644;
   wire n3645;
   wire n3646;
   wire n3647;
   wire n3648;
   wire n3649;
   wire n3650;
   wire n3651;
   wire n3652;
   wire n3653;
   wire n3654;
   wire n3655;
   wire n3656;
   wire n3657;
   wire n3658;
   wire n3659;
   wire n3660;
   wire n3661;
   wire n3662;
   wire n3663;
   wire n3664;
   wire n3665;
   wire n3666;
   wire n3667;
   wire n3668;
   wire n3669;
   wire n3670;
   wire n3671;
   wire n3672;
   wire n3673;
   wire n3674;
   wire n3675;
   wire n3676;
   wire n3677;
   wire n3678;
   wire n3679;
   wire n3680;
   wire n3681;
   wire n3682;
   wire n3683;
   wire n3684;
   wire n3685;
   wire n3686;
   wire n3687;
   wire n3688;
   wire n3689;
   wire n3690;
   wire n3691;
   wire n3692;
   wire n3693;
   wire n3694;
   wire n3695;
   wire n3696;
   wire n3697;
   wire n3698;
   wire n3699;
   wire n3700;
   wire n3701;
   wire n3702;
   wire n3703;
   wire n3704;
   wire n3705;
   wire n3706;
   wire n3707;
   wire n3708;
   wire n3709;
   wire n3710;
   wire n3711;
   wire n3712;
   wire n3713;
   wire n3714;
   wire n3715;
   wire n3716;
   wire n3717;
   wire n3718;
   wire n3719;
   wire n3720;
   wire n3721;
   wire n3722;
   wire n3723;
   wire n3724;
   wire n3725;
   wire n3726;
   wire n3727;
   wire n3728;
   wire n3729;
   wire n3730;
   wire n3731;
   wire n3732;
   wire n3733;
   wire n3734;
   wire n3735;
   wire n3736;
   wire n3737;
   wire n3738;
   wire n3739;
   wire n3740;
   wire n3741;
   wire n3742;
   wire n3743;
   wire n3744;
   wire n3745;
   wire n3746;
   wire n3747;
   wire n3748;
   wire n3749;
   wire n3750;
   wire n3751;
   wire n3752;
   wire n3753;
   wire n3754;
   wire n3755;
   wire n3756;
   wire n3757;
   wire n3758;
   wire n3759;
   wire n3760;
   wire n3761;
   wire n3762;
   wire n3763;
   wire n3764;
   wire n3765;
   wire n3766;
   wire n3767;
   wire n3768;
   wire n3769;
   wire n3770;
   wire n3771;
   wire n3772;
   wire n3773;
   wire n3774;
   wire n3775;
   wire n3776;
   wire n3777;
   wire n3778;
   wire n3779;
   wire n3780;
   wire n3781;
   wire n3782;
   wire n3783;
   wire n3784;
   wire n3785;
   wire n3786;
   wire n3787;
   wire n3788;
   wire n3789;
   wire n3790;
   wire n3791;
   wire n3792;
   wire n3793;
   wire n3794;
   wire n3795;
   wire n3796;
   wire n3797;
   wire n3798;
   wire n3799;
   wire n3800;
   wire n3801;
   wire n3802;
   wire n3803;
   wire n3804;
   wire n3805;
   wire n3806;
   wire n3807;
   wire n3808;
   wire n3809;
   wire n3810;
   wire n3811;
   wire n3812;
   wire n3813;
   wire n3814;
   wire n3815;
   wire n3816;
   wire n3817;
   wire n3818;
   wire n3819;
   wire n3820;
   wire n3821;
   wire n3822;
   wire n3823;
   wire n3824;
   wire n3825;
   wire n3826;
   wire n3827;
   wire n3828;
   wire n3829;
   wire n3830;
   wire n3831;
   wire n3832;
   wire n3833;
   wire n3834;
   wire n3835;
   wire n3836;
   wire n3837;
   wire n3838;
   wire n3839;
   wire n3840;
   wire n3841;
   wire n3842;
   wire n3843;
   wire n3844;
   wire n3845;
   wire n3846;
   wire n3847;
   wire n3848;
   wire n3849;
   wire n3850;
   wire n3851;
   wire n3852;
   wire n3853;
   wire n3854;
   wire n3855;
   wire n3856;
   wire n3857;
   wire n3858;
   wire n3859;
   wire n3860;
   wire n3861;
   wire n3862;
   wire n3863;
   wire n3864;
   wire n3865;
   wire n3866;
   wire n3867;
   wire n3868;
   wire n3869;
   wire n3870;
   wire n3871;
   wire n3872;
   wire n3873;
   wire n3874;
   wire n3875;
   wire n3876;
   wire n3877;
   wire n3878;
   wire n3879;
   wire n3880;
   wire n3881;
   wire n3882;
   wire n3883;
   wire n3884;
   wire n3885;
   wire n3886;
   wire n3887;
   wire n3888;
   wire n3889;
   wire n3890;
   wire n3891;
   wire n3892;
   wire n3893;
   wire n3894;
   wire n3895;
   wire n3896;
   wire n3897;
   wire n3898;
   wire n3899;
   wire n3900;
   wire n3901;
   wire n3902;
   wire n3903;
   wire n3904;
   wire n3905;
   wire n3906;
   wire n3907;
   wire n3908;
   wire n3909;
   wire n3910;
   wire n3911;
   wire n3912;
   wire n3913;
   wire n3914;
   wire n3915;
   wire n3916;
   wire n3917;
   wire n3918;
   wire n3919;
   wire n3920;
   wire n3921;
   wire n3922;
   wire n3923;
   wire n3924;
   wire n3925;
   wire n3926;
   wire n3927;
   wire n3928;
   wire n3929;
   wire n3930;
   wire n3931;
   wire n3932;
   wire n3933;
   wire n3934;
   wire n3935;
   wire n3936;
   wire n3937;
   wire n3938;
   wire n3939;
   wire n3940;
   wire n3941;
   wire n3942;
   wire n3943;
   wire n3944;
   wire n3945;
   wire n3946;
   wire n3947;
   wire n3948;
   wire n3949;
   wire n3950;
   wire n3951;
   wire n3952;
   wire n3953;
   wire n3954;
   wire n3955;
   wire n3956;
   wire n3957;
   wire n3958;
   wire n3959;
   wire n3960;
   wire n3961;
   wire n3962;
   wire n3963;
   wire n3964;
   wire n3965;
   wire n3966;
   wire n3967;
   wire n3968;
   wire n3969;
   wire n3970;
   wire n3971;
   wire n3972;
   wire n3973;
   wire n3974;
   wire n3975;
   wire n3976;
   wire n3977;
   wire n3978;
   wire n3979;
   wire n3980;
   wire n3981;
   wire n3982;
   wire n3983;
   wire n3984;
   wire n3985;
   wire n3986;
   wire n3987;
   wire n3988;
   wire n3989;
   wire n3990;
   wire n3991;
   wire n3992;
   wire n3993;
   wire n3994;
   wire n3995;
   wire n3996;
   wire n3997;
   wire n3998;
   wire n3999;
   wire n4000;
   wire n4001;
   wire n4002;
   wire n4003;
   wire n4004;
   wire n4005;
   wire n4006;
   wire n4007;
   wire n4008;
   wire n4009;
   wire n4010;
   wire n4011;
   wire n4012;
   wire n4013;
   wire n4014;
   wire n4015;
   wire n4016;
   wire n4017;
   wire n4018;
   wire n4019;
   wire n4020;
   wire n4021;
   wire n4022;
   wire n4023;
   wire n4024;
   wire n4025;
   wire n4026;
   wire n4027;
   wire n4028;
   wire n4029;
   wire n4030;
   wire n4031;
   wire n4032;
   wire n4033;
   wire n4034;
   wire n4035;
   wire n4036;
   wire n4037;
   wire n4038;
   wire n4039;
   wire n4040;
   wire n4041;
   wire n4042;
   wire n4043;
   wire n4044;
   wire n4045;
   wire n4046;
   wire n4047;
   wire n4048;
   wire n4049;
   wire n4050;
   wire n4051;
   wire n4052;
   wire n4053;
   wire n4054;
   wire n4055;
   wire n4056;
   wire n4057;
   wire n4058;
   wire n4059;
   wire n4060;
   wire n4061;
   wire n4062;
   wire n4063;
   wire n4064;
   wire n4065;
   wire n4066;
   wire n4067;
   wire n4068;
   wire n4069;
   wire n4070;
   wire n4071;
   wire n4072;
   wire n4073;
   wire n4074;
   wire n4075;
   wire n4076;
   wire n4077;
   wire n4078;
   wire n4079;
   wire n4080;
   wire n4081;
   wire n4082;
   wire n4083;
   wire n4084;
   wire n4085;
   wire n4086;
   wire n4087;
   wire n4088;
   wire n4089;
   wire n4090;
   wire n4091;
   wire n4092;
   wire n4093;
   wire n4094;
   wire n4095;
   wire n4096;
   wire n4097;
   wire n4098;
   wire n4099;
   wire n4100;
   wire n4101;
   wire n4102;
   wire n4103;
   wire n4104;
   wire n4105;
   wire n4106;
   wire n4107;
   wire n4108;
   wire n4109;
   wire n4110;
   wire n4111;
   wire n4112;
   wire n4113;
   wire n4114;
   wire n4115;
   wire n4116;
   wire n4117;
   wire n4118;
   wire n4119;
   wire n4120;
   wire n4121;
   wire n4122;
   wire n4123;
   wire n4124;
   wire n4125;
   wire n4126;
   wire n4127;
   wire n4128;
   wire n4129;
   wire n4130;
   wire n4131;
   wire n4132;
   wire n4133;
   wire n4134;
   wire n4135;
   wire n4136;
   wire n4137;
   wire n4138;
   wire n4139;
   wire n4140;
   wire n4141;
   wire n4142;
   wire n4143;
   wire n4144;
   wire n4145;
   wire n4146;
   wire n4147;
   wire n4148;
   wire n4149;
   wire n4150;
   wire n4151;
   wire n4152;
   wire n4153;
   wire n4154;
   wire n4155;
   wire n4156;
   wire n4157;
   wire n4158;
   wire n4159;
   wire n4160;
   wire n4161;
   wire n4162;
   wire n4163;
   wire n4164;
   wire n4165;
   wire n4166;
   wire n4167;
   wire n4168;
   wire n4169;
   wire n4170;
   wire n4171;
   wire n4172;
   wire n4173;
   wire n4174;
   wire n4175;
   wire n4176;
   wire n4177;
   wire n4178;
   wire n4179;
   wire n4180;
   wire n4181;
   wire n4182;
   wire n4183;
   wire n4184;
   wire n4185;
   wire n4186;
   wire n4187;
   wire n4188;
   wire n4189;
   wire n4190;
   wire n4191;
   wire n4192;
   wire n4193;
   wire n4194;
   wire n4195;
   wire n4196;
   wire n4197;
   wire n4198;
   wire n4199;
   wire n4200;
   wire n4201;
   wire n4202;
   wire n4203;
   wire n4204;
   wire n4205;
   wire n4206;
   wire n4207;
   wire n4208;
   wire n4209;
   wire n4210;
   wire n4211;
   wire n4212;
   wire n4213;
   wire n4214;
   wire n4215;
   wire n4216;
   wire n4217;
   wire n4218;
   wire n4219;
   wire n4220;
   wire n4221;
   wire n4222;
   wire n4223;
   wire n4224;
   wire n4225;
   wire n4226;
   wire n4227;
   wire n4228;
   wire n4229;
   wire n4230;
   wire n4231;
   wire n4232;
   wire n4233;
   wire n4234;
   wire n4235;
   wire n4236;
   wire n4237;
   wire n4238;
   wire n4239;
   wire n4240;
   wire n4241;
   wire n4242;
   wire n4243;
   wire n4244;
   wire n4245;
   wire n4246;
   wire n4247;
   wire n4248;
   wire n4249;
   wire n4250;
   wire n4251;
   wire n4252;
   wire n4253;
   wire n4254;
   wire n4255;
   wire n4256;
   wire n4257;
   wire n4258;
   wire n4259;
   wire n4260;
   wire n4261;
   wire n4262;
   wire n4263;
   wire n4264;
   wire n4265;
   wire n4266;
   wire n4267;
   wire n4268;
   wire n4269;
   wire n4270;
   wire n4271;
   wire n4272;
   wire n4273;
   wire n4274;
   wire n4275;
   wire n4276;
   wire n4277;
   wire n4278;
   wire n4279;
   wire n4280;
   wire n4281;
   wire n4282;
   wire n4283;
   wire n4284;
   wire n4285;
   wire n4286;
   wire n4287;
   wire n4288;
   wire n4289;
   wire n4290;
   wire n4291;
   wire n4292;
   wire n4293;
   wire n4294;
   wire n4295;
   wire n4296;
   wire n4297;
   wire n4298;
   wire n4299;
   wire n4300;
   wire n4301;
   wire n4302;
   wire n4303;
   wire n4304;
   wire n4305;
   wire n4306;
   wire n4307;
   wire n4308;
   wire n4309;
   wire n4310;
   wire n4311;
   wire n4312;
   wire n4313;
   wire n4314;
   wire n4315;
   wire n4316;
   wire n4317;
   wire n4318;
   wire n4319;
   wire n4320;
   wire n4321;
   wire n4322;
   wire n4323;
   wire n4324;
   wire n4325;
   wire n4326;
   wire n4327;
   wire n4328;
   wire n4329;
   wire n4330;
   wire n4331;
   wire n4332;
   wire n4333;
   wire n4334;
   wire n4335;
   wire n4336;
   wire n4337;
   wire n4338;
   wire n4339;
   wire n4340;
   wire n4341;
   wire n4342;
   wire n4343;
   wire n4344;
   wire n4345;
   wire n4346;
   wire n4347;
   wire n4348;
   wire n4349;
   wire n4350;
   wire n4351;
   wire n4352;
   wire n4353;
   wire n4354;
   wire n4355;
   wire n4356;
   wire n4357;
   wire n4358;
   wire n4359;
   wire n4360;
   wire n4361;
   wire n4362;
   wire n4363;
   wire n4364;
   wire n4365;
   wire n4366;
   wire n4367;
   wire n4368;
   wire n4369;
   wire n4370;
   wire n4371;
   wire n4372;
   wire n4373;
   wire n4374;
   wire n4375;
   wire n4376;
   wire n4377;
   wire n4378;
   wire n4379;
   wire n4380;
   wire n4381;
   wire n4382;
   wire n4383;
   wire n4384;
   wire n4385;
   wire n4386;
   wire n4387;
   wire n4388;
   wire n4389;
   wire n4390;
   wire n4391;
   wire n4392;
   wire n4393;
   wire n4394;
   wire n4395;
   wire n4396;
   wire n4397;
   wire n4398;
   wire n4399;
   wire n4400;
   wire n4401;
   wire n4402;
   wire n4403;
   wire n4404;
   wire n4405;
   wire n4406;
   wire n4407;
   wire n4408;
   wire n4409;
   wire n4410;
   wire n4411;
   wire n4412;
   wire n4413;
   wire n4414;
   wire n4415;
   wire n4416;
   wire n4417;
   wire n4418;
   wire n4419;
   wire n4420;
   wire n4421;
   wire n4422;
   wire n4423;
   wire n4424;
   wire n4425;
   wire n4426;
   wire n4427;
   wire n4428;
   wire n4429;
   wire n4430;
   wire n4431;
   wire n4432;
   wire n4433;
   wire n4434;
   wire n4435;
   wire n4436;
   wire n4437;
   wire n4438;
   wire n4439;
   wire n4440;
   wire n4441;
   wire n4442;
   wire n4443;
   wire n4444;
   wire n4445;
   wire n4446;
   wire n4447;
   wire n4448;
   wire n4449;
   wire n4450;
   wire n4451;
   wire n4452;
   wire n4453;
   wire n4454;
   wire n4455;
   wire n4456;
   wire n4457;
   wire n4458;
   wire n4459;
   wire n4460;
   wire n4461;
   wire n4462;
   wire n4463;
   wire n4464;
   wire n4465;
   wire n4466;
   wire n4467;
   wire n4468;
   wire n4469;
   wire n4470;
   wire n4471;
   wire n4472;
   wire n4473;
   wire n4474;
   wire n4475;
   wire n4476;
   wire n4477;
   wire n4478;
   wire n4479;
   wire n4480;
   wire n4481;
   wire n4482;
   wire n4483;
   wire n4484;
   wire n4485;
   wire n4486;
   wire n4487;
   wire n4488;
   wire n4489;
   wire n4490;
   wire n4491;
   wire n4492;
   wire n4493;
   wire n4494;
   wire n4495;
   wire n4496;
   wire n4497;
   wire n4498;
   wire n4499;
   wire n4500;
   wire n4501;
   wire n4502;
   wire n4503;
   wire n4504;
   wire n4505;
   wire n4506;
   wire n4507;
   wire n4508;
   wire n4509;
   wire n4510;
   wire n4511;
   wire n4512;
   wire n4513;
   wire n4514;
   wire n4515;
   wire n4516;
   wire n4517;
   wire n4518;
   wire n4519;
   wire n4520;
   wire n4521;
   wire n4522;
   wire n4523;
   wire n4524;
   wire n4525;
   wire n4526;
   wire n4527;
   wire n4528;
   wire n4529;
   wire n4530;
   wire n4531;
   wire n4532;
   wire n4533;
   wire n4534;
   wire n4535;
   wire n4536;
   wire n4537;
   wire n4538;
   wire n4539;
   wire n4540;
   wire n4541;
   wire n4542;
   wire n4543;
   wire n4544;
   wire n4545;
   wire n4546;
   wire n4547;
   wire n4548;
   wire n4549;
   wire n4550;
   wire n4551;
   wire n4552;
   wire n4553;
   wire n4554;
   wire n4555;
   wire n4556;
   wire n4557;
   wire n4558;
   wire n4559;
   wire n4560;
   wire n4561;
   wire n4562;
   wire n4563;
   wire n4564;
   wire n4565;
   wire n4566;
   wire n4567;
   wire n4568;
   wire n4569;
   wire n4570;
   wire n4571;
   wire n4572;
   wire n4573;
   wire n4574;
   wire n4575;
   wire n4576;
   wire n4577;
   wire n4578;
   wire n4579;
   wire n4580;
   wire n4581;
   wire n4582;
   wire n4583;
   wire n4584;
   wire n4585;
   wire n4586;
   wire n4587;
   wire n4588;
   wire n4589;
   wire n4590;
   wire n4591;
   wire n4592;
   wire n4593;
   wire n4594;
   wire n4595;
   wire n4596;
   wire n4597;
   wire n4598;
   wire n4599;
   wire n4600;
   wire n4601;
   wire n4602;
   wire n4603;
   wire n4604;
   wire n4605;
   wire n4606;
   wire n4607;
   wire n4608;
   wire n4609;
   wire n4610;
   wire n4611;
   wire n4612;
   wire n4613;
   wire n4614;
   wire n4615;
   wire n4616;
   wire n4617;
   wire n4618;
   wire n4619;
   wire n4620;
   wire n4621;
   wire n4622;
   wire n4623;
   wire n4624;
   wire n4625;
   wire n4626;
   wire n4627;
   wire n4628;
   wire n4629;
   wire n4630;
   wire n4631;
   wire n4632;
   wire n4633;
   wire n4634;
   wire n4635;
   wire n4636;
   wire n4637;
   wire n4638;
   wire n4639;
   wire n4640;
   wire n4641;
   wire n4642;
   wire n4643;
   wire n4644;
   wire n4645;
   wire n4646;
   wire n4647;
   wire n4648;
   wire n4649;
   wire n4650;
   wire n4651;
   wire n4652;
   wire n4653;
   wire n4654;
   wire n4655;
   wire n4656;
   wire n4657;
   wire n4658;
   wire n4659;
   wire n4660;
   wire n4661;
   wire n4662;
   wire n4663;
   wire n4664;
   wire n4665;
   wire n4666;
   wire n4667;
   wire n4668;
   wire n4669;
   wire n4670;
   wire n4671;
   wire n4672;
   wire n4673;
   wire n4674;
   wire n4675;
   wire n4676;
   wire n4677;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n7;
   wire n24;
   wire n25;
   wire n26;
   wire n28;
   wire n29;
   wire n31;
   wire n32;
   wire n34;
   wire n35;
   wire n37;
   wire n38;
   wire n40;
   wire n41;
   wire n43;
   wire n44;
   wire n46;
   wire n47;
   wire n49;
   wire n50;
   wire n52;
   wire n53;
   wire n55;
   wire n56;
   wire n58;
   wire n59;
   wire n61;
   wire n62;
   wire n64;
   wire n65;
   wire n67;
   wire n68;
   wire n70;
   wire n73;
   wire n75;
   wire n76;
   wire n78;
   wire n80;
   wire n82;
   wire n84;
   wire n86;
   wire n88;
   wire n90;
   wire n92;
   wire n94;
   wire n96;
   wire n98;
   wire n100;
   wire n102;
   wire n104;
   wire n107;
   wire n109;
   wire n110;
   wire n112;
   wire n114;
   wire n116;
   wire n118;
   wire n120;
   wire n122;
   wire n124;
   wire n126;
   wire n128;
   wire n130;
   wire n132;
   wire n134;
   wire n136;
   wire n138;
   wire n141;
   wire n143;
   wire n144;
   wire n146;
   wire n148;
   wire n150;
   wire n152;
   wire n154;
   wire n156;
   wire n158;
   wire n160;
   wire n162;
   wire n164;
   wire n166;
   wire n168;
   wire n170;
   wire n172;
   wire n175;
   wire n177;
   wire n178;
   wire n180;
   wire n182;
   wire n184;
   wire n186;
   wire n188;
   wire n190;
   wire n192;
   wire n194;
   wire n196;
   wire n198;
   wire n200;
   wire n202;
   wire n204;
   wire n206;
   wire n209;
   wire n211;
   wire n212;
   wire n214;
   wire n216;
   wire n218;
   wire n220;
   wire n222;
   wire n224;
   wire n226;
   wire n228;
   wire n230;
   wire n232;
   wire n234;
   wire n236;
   wire n238;
   wire n240;
   wire n242;
   wire n244;
   wire n245;
   wire n247;
   wire n249;
   wire n251;
   wire n253;
   wire n255;
   wire n257;
   wire n259;
   wire n261;
   wire n263;
   wire n265;
   wire n267;
   wire n269;
   wire n271;
   wire n273;
   wire n275;
   wire n277;
   wire n278;
   wire n280;
   wire n282;
   wire n284;
   wire n286;
   wire n288;
   wire n290;
   wire n292;
   wire n294;
   wire n296;
   wire n298;
   wire n300;
   wire n302;
   wire n304;
   wire n306;
   wire n308;
   wire n310;
   wire n311;
   wire n313;
   wire n315;
   wire n317;
   wire n319;
   wire n321;
   wire n323;
   wire n325;
   wire n327;
   wire n329;
   wire n331;
   wire n333;
   wire n335;
   wire n337;
   wire n339;
   wire n342;
   wire n344;
   wire n345;
   wire n347;
   wire n349;
   wire n351;
   wire n353;
   wire n355;
   wire n357;
   wire n359;
   wire n361;
   wire n363;
   wire n365;
   wire n367;
   wire n369;
   wire n371;
   wire n373;
   wire n375;
   wire n377;
   wire n378;
   wire n380;
   wire n382;
   wire n384;
   wire n386;
   wire n388;
   wire n390;
   wire n392;
   wire n394;
   wire n396;
   wire n398;
   wire n400;
   wire n402;
   wire n404;
   wire n406;
   wire n408;
   wire n410;
   wire n411;
   wire n413;
   wire n415;
   wire n417;
   wire n419;
   wire n421;
   wire n423;
   wire n425;
   wire n427;
   wire n429;
   wire n431;
   wire n433;
   wire n435;
   wire n437;
   wire n439;
   wire n441;
   wire n443;
   wire n444;
   wire n446;
   wire n448;
   wire n450;
   wire n452;
   wire n454;
   wire n456;
   wire n458;
   wire n460;
   wire n462;
   wire n464;
   wire n466;
   wire n468;
   wire n470;
   wire n472;
   wire n475;
   wire n477;
   wire n478;
   wire n480;
   wire n482;
   wire n484;
   wire n486;
   wire n488;
   wire n490;
   wire n492;
   wire n494;
   wire n496;
   wire n498;
   wire n500;
   wire n502;
   wire n504;
   wire n506;
   wire n508;
   wire n510;
   wire n511;
   wire n513;
   wire n515;
   wire n517;
   wire n519;
   wire n521;
   wire n523;
   wire n525;
   wire n527;
   wire n529;
   wire n531;
   wire n533;
   wire n535;
   wire n537;
   wire n539;
   wire n541;
   wire n543;
   wire n546;
   wire n549;
   wire n552;
   wire n555;
   wire n558;
   wire n560;
   wire n562;
   wire n564;
   wire n567;
   wire n569;
   wire n571;
   wire n573;
   wire n576;
   wire n578;
   wire n580;
   wire n4678;
   wire n4679;
   wire n4680;
   wire n4681;
   wire n4682;
   wire n4683;
   wire n4684;
   wire n4685;
   wire n4686;
   wire n4687;
   wire n4688;
   wire n4689;
   wire n4690;
   wire n4691;
   wire n4692;
   wire n4693;
   wire n4694;
   wire n4695;
   wire n4696;
   wire n4697;
   wire n4698;
   wire n4699;
   wire n4700;
   wire n4701;
   wire n4702;
   wire n4703;
   wire n4704;
   wire n4705;
   wire n4706;
   wire n4707;
   wire n4708;
   wire n4709;
   wire n4710;
   wire n4711;
   wire n4712;
   wire n4713;
   wire n4714;
   wire n4715;
   wire n4716;
   wire n4717;
   wire n4718;
   wire n4719;
   wire n4720;
   wire n4721;
   wire n4722;
   wire n4723;
   wire n4724;
   wire n4725;
   wire n4726;
   wire n4727;
   wire n4728;
   wire n4729;
   wire n4730;
   wire n4731;
   wire n4732;
   wire n4733;
   wire n4734;
   wire n4735;
   wire n4736;
   wire n4737;
   wire n4738;
   wire n4739;
   wire n4740;
   wire n4741;
   wire n4742;
   wire n4743;
   wire n4744;
   wire n4745;
   wire n4746;
   wire n4747;
   wire n4748;
   wire n4749;
   wire n4750;
   wire n4751;
   wire n4752;
   wire n4753;
   wire n4754;
   wire n4755;
   wire n4756;
   wire n4757;
   wire n4758;
   wire n4759;
   wire n4760;
   wire n4761;
   wire n4762;
   wire n4763;
   wire n4764;
   wire n4765;
   wire n4766;
   wire n4767;
   wire n4768;
   wire n4769;
   wire n4770;
   wire n4771;
   wire n4772;
   wire n4773;
   wire n4774;
   wire n4775;
   wire n4776;
   wire n4777;
   wire n4778;
   wire n4779;
   wire n4780;
   wire n4781;
   wire n4782;
   wire n4783;
   wire n4784;
   wire n4785;
   wire n4786;
   wire n4787;
   wire n4788;
   wire n4789;
   wire n4790;
   wire n4791;
   wire n4792;
   wire n4793;
   wire n4794;
   wire n4795;
   wire n4796;
   wire n4797;
   wire n4798;
   wire n4799;
   wire n4800;
   wire n4801;
   wire n4802;
   wire n4803;
   wire n4804;
   wire n4805;
   wire n4806;
   wire n4807;
   wire n4808;
   wire n4809;
   wire n4810;
   wire n4811;
   wire n4812;
   wire n4813;
   wire n4814;
   wire n4815;
   wire n4816;
   wire n4817;
   wire n4818;
   wire n4819;
   wire n4820;
   wire n4821;
   wire n4822;
   wire n4823;
   wire n4824;
   wire n4825;
   wire n4826;
   wire n4827;
   wire n4828;
   wire n4829;
   wire n4830;
   wire n4831;
   wire n4832;
   wire n4833;
   wire n4834;
   wire n4835;
   wire n4836;
   wire n4837;
   wire n4838;
   wire n4839;
   wire n4840;
   wire n4841;
   wire n4842;
   wire n4843;
   wire n4844;
   wire n4845;
   wire n4846;
   wire n4847;
   wire n4848;
   wire n4849;
   wire n4850;
   wire n4851;
   wire n4852;
   wire n4853;
   wire n4854;
   wire n4855;
   wire n4856;
   wire n4857;
   wire n4858;
   wire n4859;
   wire n4860;
   wire n4861;
   wire n4862;
   wire n4863;
   wire n4864;
   wire n4865;
   wire n4866;
   wire n4867;
   wire n4868;
   wire n4869;
   wire n4870;
   wire n4871;
   wire n4872;
   wire n4873;
   wire n4874;
   wire n4875;
   wire n4876;
   wire n4877;
   wire n4878;
   wire n4879;
   wire n4880;
   wire n4881;
   wire n4882;
   wire n4883;
   wire n4884;
   wire n4885;
   wire n4886;
   wire n4887;
   wire n4888;
   wire n4889;
   wire n4890;
   wire n4891;
   wire n4892;
   wire n4893;
   wire n4894;
   wire n4895;
   wire n4896;
   wire n4897;
   wire n4898;
   wire n4899;
   wire n4900;
   wire n4901;
   wire n4902;
   wire n4903;
   wire n4904;
   wire n4905;
   wire n4906;
   wire n4907;
   wire n4908;
   wire n4909;
   wire n4910;
   wire n4911;
   wire n4912;
   wire n4913;
   wire n4914;
   wire n4915;
   wire n4916;
   wire n4917;
   wire n4918;
   wire n4919;
   wire n4920;
   wire n4921;
   wire n4922;
   wire n4923;
   wire n4924;
   wire n4925;
   wire n4926;
   wire n4927;
   wire n4928;
   wire n4929;
   wire n4930;
   wire n4931;
   wire n4932;
   wire n4933;
   wire n4934;
   wire n4935;
   wire n4936;
   wire n4937;
   wire n4938;
   wire n4939;
   wire n4940;
   wire n4941;
   wire n4942;
   wire n4943;
   wire n4944;
   wire n4945;
   wire n4946;
   wire n4947;
   wire n4948;
   wire n4949;
   wire n4950;
   wire n4951;
   wire n4952;
   wire n4953;
   wire n4954;
   wire n4955;
   wire n4956;
   wire n4957;
   wire n4958;
   wire n4959;
   wire n4960;
   wire n4961;
   wire n4962;
   wire n4963;
   wire n4964;
   wire n4965;
   wire n4966;
   wire n4967;
   wire n4968;
   wire n4969;
   wire n4970;
   wire n4971;
   wire n4972;
   wire n4973;
   wire n4974;
   wire n4975;
   wire n4976;
   wire n4977;
   wire n4978;
   wire n4979;
   wire n4980;
   wire n4981;
   wire n4982;
   wire n4983;
   wire n4984;
   wire n4985;
   wire n4986;
   wire n4987;
   wire n4988;
   wire n4989;
   wire n4990;
   wire n4991;
   wire n4992;
   wire n4993;
   wire n4994;
   wire n4995;
   wire n4996;
   wire n4997;
   wire n4998;
   wire n4999;
   wire n5000;
   wire n5001;
   wire n5002;
   wire n5003;
   wire n5004;
   wire n5005;
   wire n5006;
   wire n5007;
   wire n5008;
   wire n5009;
   wire n5010;
   wire n5011;
   wire n5012;
   wire n5013;
   wire n5014;
   wire n5015;
   wire n5016;
   wire n5017;
   wire n5018;
   wire n5019;
   wire n5020;
   wire n5021;
   wire n5022;
   wire n5023;
   wire n5024;
   wire n5025;
   wire n5026;
   wire n5027;
   wire n5028;
   wire n5029;
   wire n5030;
   wire n5031;
   wire n5032;
   wire n5033;
   wire n5034;
   wire n5035;
   wire n5036;
   wire n5037;
   wire n5038;
   wire n5039;
   wire n5040;
   wire n5041;
   wire n5042;
   wire n5043;
   wire n5044;
   wire n5045;
   wire n5046;
   wire n5047;
   wire n5048;
   wire n5049;
   wire n5050;
   wire n5051;
   wire n5052;
   wire n5053;
   wire n5054;
   wire n5055;
   wire n5056;
   wire n5057;
   wire n5058;
   wire n5059;
   wire n5060;
   wire n5061;
   wire n5062;
   wire n5063;
   wire n5064;
   wire n5065;
   wire n5066;
   wire n5067;
   wire n5068;
   wire n5069;
   wire n5070;
   wire n5071;
   wire n5072;
   wire n5073;
   wire n5074;
   wire n5075;
   wire n5076;
   wire n5077;
   wire n5078;
   wire n5079;
   wire n5080;
   wire n5081;
   wire n5082;
   wire n5083;
   wire n5084;
   wire n5085;
   wire n5086;
   wire n5087;
   wire n5088;
   wire n5089;
   wire n5090;
   wire n5091;
   wire n5092;
   wire n5093;
   wire n5094;
   wire n5095;
   wire n5096;
   wire n5097;
   wire n5098;
   wire n5099;
   wire n5100;
   wire n5101;
   wire n5102;
   wire n5103;
   wire n5104;
   wire n5105;
   wire n5106;
   wire n5107;
   wire n5108;
   wire n5109;
   wire n5110;
   wire n5111;
   wire n5112;
   wire n5113;
   wire n5114;
   wire n5115;
   wire n5116;
   wire n5117;
   wire n5118;
   wire n5119;
   wire n5120;
   wire n5121;
   wire n5122;
   wire n5123;
   wire n5124;
   wire n5125;
   wire n5126;
   wire n5127;
   wire n5128;
   wire n5129;
   wire n5130;
   wire n5131;
   wire n5132;
   wire n5133;
   wire n5134;
   wire n5135;
   wire n5136;
   wire n5137;
   wire n5138;
   wire n5139;
   wire n5140;
   wire n5141;
   wire n5142;
   wire n5143;
   wire n5144;
   wire n5145;
   wire n5146;
   wire n5147;
   wire n5148;
   wire n5149;
   wire n5150;
   wire n5151;
   wire n5152;
   wire n5153;
   wire n5154;
   wire n5155;
   wire n5156;
   wire n5157;
   wire n5158;
   wire n5159;
   wire n5160;
   wire n5161;
   wire n5162;
   wire n5163;
   wire n5164;
   wire n5165;
   wire n5166;
   wire n5167;
   wire n5168;
   wire n5169;
   wire n5170;
   wire n5171;
   wire n5172;
   wire n5173;
   wire n5174;
   wire n5175;
   wire n5176;
   wire n5177;
   wire n5178;
   wire n5179;
   wire n5180;
   wire n5181;
   wire n5182;
   wire n5183;
   wire n5184;
   wire n5185;
   wire n5186;
   wire n5187;
   wire n5188;
   wire n5189;
   wire n5190;
   wire n5191;
   wire n5192;
   wire n5193;
   wire n5194;
   wire n5195;
   wire n5196;
   wire n5197;
   wire n5198;
   wire n5199;
   wire n5200;
   wire n5201;
   wire n5202;
   wire n5203;
   wire n5204;
   wire n5205;
   wire n5206;
   wire n5207;
   wire n5208;
   wire n5209;
   wire n5210;
   wire n5211;
   wire n5212;
   wire n5213;
   wire n5214;
   wire n5215;
   wire n5216;
   wire n5217;
   wire n5218;
   wire n5219;
   wire n5220;
   wire n5221;
   wire n5222;
   wire n5223;
   wire n5224;
   wire n5225;
   wire n5226;
   wire n5227;
   wire n5228;
   wire n5229;
   wire n5230;
   wire n5231;
   wire n5232;
   wire n5233;
   wire n5234;
   wire n5235;
   wire n5236;
   wire n5237;
   wire n5238;
   wire n5239;
   wire n5240;
   wire n5241;
   wire n5242;
   wire n5243;
   wire n5244;
   wire n5245;
   wire n5246;
   wire n5247;
   wire n5248;
   wire n5249;
   wire n5250;
   wire n5251;
   wire n5252;
   wire n5253;
   wire n5254;
   wire n5255;
   wire n5256;
   wire n5257;
   wire n5258;
   wire n5259;
   wire n5260;
   wire n5261;
   wire n5262;
   wire n5263;
   wire n5264;
   wire n5265;
   wire n5266;
   wire n5267;
   wire n5268;
   wire n5269;
   wire n5270;
   wire n5271;
   wire n5272;
   wire n5273;
   wire n5274;
   wire n5275;
   wire n5276;
   wire n5277;
   wire n5278;
   wire n5279;
   wire n5280;
   wire n5281;
   wire n5282;
   wire n5283;
   wire n5284;
   wire n5285;
   wire n5286;
   wire n5287;
   wire n5288;
   wire n5289;
   wire n5290;
   wire n5291;
   wire n5292;
   wire n5293;
   wire n5294;
   wire n5295;
   wire n5296;
   wire n5297;
   wire n5298;
   wire n5299;
   wire n5300;
   wire n5301;
   wire n5302;
   wire n5303;
   wire n5304;
   wire n5305;
   wire n5306;
   wire n5307;
   wire n5308;
   wire n5309;
   wire n5310;
   wire n5311;
   wire n5312;
   wire n5313;
   wire n5314;
   wire n5315;
   wire n5316;
   wire n5317;
   wire n5318;
   wire n5319;
   wire n5320;
   wire n5321;
   wire n5322;
   wire n5323;
   wire n5324;
   wire n5325;
   wire n5326;
   wire n5327;
   wire n5328;
   wire n5329;
   wire n5330;
   wire n5331;
   wire n5332;
   wire n5333;
   wire n5334;
   wire n5335;
   wire n5336;
   wire n5337;
   wire n5338;
   wire n5339;
   wire n5340;
   wire n5341;
   wire n5342;
   wire n5343;
   wire n5344;
   wire n5345;
   wire n5346;
   wire n5347;
   wire n5348;
   wire n5349;
   wire n5350;
   wire n5351;
   wire n5352;
   wire n5353;
   wire n5354;
   wire n5355;
   wire n5356;
   wire n5357;
   wire n5358;
   wire n5359;
   wire n5360;
   wire n5361;
   wire n5362;
   wire n5363;
   wire n5364;
   wire n5365;
   wire n5366;
   wire n5367;
   wire n5368;
   wire n5369;
   wire n5370;
   wire n5371;
   wire n5372;
   wire n5373;
   wire n5374;
   wire n5375;
   wire n5376;
   wire n5377;
   wire n5378;
   wire n5379;
   wire n5380;
   wire n5381;
   wire n5382;
   wire n5383;
   wire n5384;
   wire n5385;
   wire n5386;
   wire n5387;
   wire n5388;
   wire n5389;
   wire n5390;
   wire n5391;
   wire n5392;
   wire n5393;
   wire n5394;
   wire n5395;
   wire n5396;
   wire n5397;
   wire n5398;
   wire n5399;
   wire n5400;
   wire n5401;
   wire n5402;
   wire n5403;
   wire n5404;
   wire n5405;
   wire n5406;
   wire n5407;
   wire n5408;
   wire n5409;
   wire n5410;
   wire n5411;
   wire n5412;
   wire n5413;
   wire n5414;
   wire n5415;
   wire n5416;
   wire n5417;
   wire n5418;
   wire n5419;
   wire n5420;
   wire n5421;
   wire n5422;
   wire n5423;
   wire n5424;
   wire n5425;
   wire n5426;
   wire n5427;
   wire n5428;
   wire n5429;
   wire n5430;
   wire n5431;
   wire n5432;
   wire n5433;
   wire n5434;
   wire n5435;
   wire n5436;
   wire n5437;
   wire n5438;
   wire n5439;
   wire n5440;
   wire n5441;
   wire n5442;
   wire n5443;
   wire n5444;
   wire n5445;
   wire n5446;
   wire n5447;
   wire n5448;
   wire n5449;
   wire n5450;
   wire n5451;
   wire n5452;
   wire n5453;
   wire n5454;
   wire n5455;
   wire n5456;
   wire n5457;
   wire n5458;
   wire n5459;
   wire n5460;
   wire n5461;
   wire n5462;
   wire n5463;
   wire n5464;
   wire n5465;
   wire n5466;
   wire n5467;
   wire n5468;
   wire n5469;
   wire n5470;
   wire n5471;
   wire n5472;
   wire n5473;
   wire n5474;
   wire n5475;
   wire n5476;
   wire n5477;
   wire n5478;
   wire n5479;
   wire n5480;
   wire n5481;
   wire n5482;
   wire n5483;
   wire n5484;
   wire n5485;
   wire n5486;
   wire n5487;
   wire n5488;
   wire n5489;
   wire n5490;
   wire n5491;
   wire n5492;
   wire n5493;
   wire n5494;
   wire n5495;
   wire n5496;
   wire n5497;
   wire n5498;
   wire n5499;
   wire n5500;
   wire n5501;
   wire n5502;
   wire n5503;
   wire n5504;
   wire n5505;
   wire n5506;
   wire n5507;
   wire n5508;
   wire n5509;
   wire n5510;
   wire n5511;
   wire n5512;
   wire n5513;
   wire n5514;
   wire n5515;
   wire n5516;
   wire n5517;
   wire n5518;
   wire n5519;
   wire n5520;
   wire n5521;
   wire n5522;
   wire n5523;
   wire n5524;
   wire n5525;
   wire n5526;
   wire n5527;
   wire n5528;
   wire n5529;
   wire n5530;
   wire n5531;
   wire n5532;
   wire n5533;
   wire n5534;
   wire n5535;
   wire n5536;
   wire n5537;
   wire n5538;
   wire n5539;
   wire n5540;
   wire n5541;
   wire n5542;
   wire n5543;
   wire n5544;
   wire n5545;
   wire n5546;
   wire n5547;
   wire n5548;
   wire n5549;
   wire n5550;
   wire n5551;
   wire n5552;
   wire n5553;
   wire n5554;
   wire n5555;
   wire n5556;
   wire n5557;
   wire n5558;
   wire n5559;
   wire n5560;
   wire n5561;
   wire n5562;
   wire n5563;
   wire n5564;
   wire n5565;
   wire n5566;
   wire n5567;
   wire n5568;
   wire n5569;
   wire n5570;
   wire n5571;
   wire n5572;
   wire n5573;
   wire n5574;
   wire n5575;
   wire n5576;
   wire n5577;
   wire n5578;
   wire n5579;
   wire n5580;
   wire n5581;
   wire n5582;
   wire n5583;
   wire n5584;
   wire n5585;
   wire n5586;
   wire n5587;
   wire n5588;
   wire n5589;
   wire n5590;
   wire n5591;
   wire n5592;
   wire n5593;
   wire n5594;
   wire n5595;
   wire n5596;
   wire n5597;
   wire n5598;
   wire n5599;
   wire n5600;
   wire n5601;
   wire n5602;
   wire n5603;
   wire n5604;
   wire n5605;
   wire n5606;
   wire n5607;
   wire n5608;
   wire n5609;
   wire n5610;
   wire n5611;
   wire n5612;
   wire n5613;
   wire n5614;
   wire n5615;
   wire n5616;
   wire n5617;
   wire n5618;
   wire n5619;
   wire n5620;
   wire n5621;
   wire n5622;
   wire n5623;
   wire n5624;
   wire n5625;
   wire n5626;
   wire n5627;
   wire n5628;
   wire n5629;
   wire n5630;
   wire n5631;
   wire n5632;
   wire n5633;
   wire n5634;
   wire n5635;
   wire n5636;
   wire n5637;
   wire n5638;
   wire n5639;
   wire n5640;
   wire n5641;
   wire n5642;
   wire n5643;
   wire n5644;
   wire n5645;
   wire n5646;
   wire n5647;
   wire n5648;
   wire n5649;
   wire n5650;
   wire n5651;
   wire n5652;
   wire n5653;
   wire n5654;
   wire n5655;
   wire n5656;
   wire n5657;
   wire n5658;
   wire n5659;
   wire n5660;
   wire n5661;
   wire n5662;
   wire n5663;
   wire n5664;
   wire n5665;
   wire n5666;
   wire n5667;
   wire n5668;
   wire n5669;
   wire n5670;
   wire n5671;
   wire n5672;
   wire n5673;
   wire n5674;
   wire n5675;
   wire n5676;
   wire n5677;
   wire n5678;
   wire n5679;
   wire n5680;
   wire n5681;
   wire n5682;
   wire n5683;
   wire n5684;
   wire n5685;
   wire n5686;
   wire n5687;
   wire n5688;
   wire n5689;
   wire n5690;
   wire n5691;
   wire n5692;
   wire n5693;
   wire n5694;
   wire n5695;
   wire n5696;
   wire n5697;
   wire n5698;
   wire n5699;
   wire n5700;
   wire n5701;
   wire n5702;
   wire n5703;
   wire n5704;
   wire n5705;
   wire n5706;
   wire n5707;
   wire n5708;
   wire n5709;
   wire n5710;
   wire n5711;
   wire n5712;
   wire n5713;
   wire n5714;
   wire n5715;
   wire n5716;
   wire n5717;
   wire n5718;
   wire n5719;
   wire n5720;
   wire n5721;
   wire n5722;
   wire n5723;
   wire n5724;
   wire n5725;
   wire n5726;
   wire n5727;
   wire n5728;
   wire n5729;
   wire n5730;
   wire n5731;
   wire n5732;
   wire n5733;
   wire n5734;
   wire n5735;
   wire n5736;
   wire n5737;
   wire n5738;
   wire n5739;
   wire n5740;
   wire n5741;
   wire n5742;
   wire n5743;
   wire n5744;
   wire n5745;
   wire n5746;
   wire n5747;
   wire n5748;
   wire n5749;
   wire n5750;
   wire n5751;
   wire n5752;
   wire n5753;
   wire n5754;
   wire n5755;
   wire n5756;
   wire n5757;
   wire n5758;
   wire n5759;
   wire n5760;
   wire n5761;
   wire n5762;
   wire n5763;
   wire n5764;
   wire n5765;
   wire n5766;
   wire n5767;
   wire n5768;
   wire n5769;
   wire n5770;
   wire n5771;
   wire n5772;
   wire n5773;
   wire n5774;
   wire n5775;
   wire n5776;
   wire n5777;
   wire n5778;
   wire n5779;
   wire n5780;
   wire n5781;
   wire n5782;
   wire n5783;
   wire n5784;
   wire n5785;
   wire n5786;
   wire n5787;
   wire n5788;
   wire n5789;
   wire n5790;
   wire n5791;
   wire n5792;
   wire n5793;
   wire n5794;
   wire n5795;
   wire n5796;
   wire n5797;
   wire n5798;
   wire n5799;
   wire n5800;
   wire n5801;
   wire n5802;
   wire n5803;
   wire n5804;
   wire n5805;
   wire n5806;
   wire n5807;
   wire n5808;
   wire n5809;
   wire n5810;
   wire n5811;
   wire n5812;
   wire n5813;
   wire n5814;
   wire n5815;
   wire n5816;
   wire n5817;
   wire n5818;
   wire n5819;
   wire n5820;
   wire n5821;
   wire n5822;
   wire n5823;
   wire n5824;
   wire n5825;
   wire n5826;
   wire n5827;
   wire n5828;
   wire n5829;
   wire n5830;
   wire n5831;
   wire n5832;
   wire n5833;
   wire n5834;
   wire n5835;
   wire n5836;
   wire n5837;
   wire n5838;
   wire n5839;
   wire n5840;
   wire n5841;
   wire n5842;
   wire n5843;
   wire n5844;
   wire n5845;
   wire n5846;
   wire n5847;
   wire n5848;
   wire n5849;
   wire n5850;
   wire n5851;
   wire n5852;
   wire n5853;
   wire n5854;
   wire n5855;
   wire n5856;
   wire n5857;
   wire n5858;
   wire n5859;
   wire n5860;
   wire n5861;
   wire n5862;
   wire n5863;
   wire n5864;
   wire n5865;
   wire n5866;
   wire n5867;
   wire n5868;
   wire n5869;
   wire n5870;
   wire n5871;
   wire n5872;
   wire n5873;
   wire n5874;
   wire n5875;
   wire n5876;
   wire n5877;
   wire n5878;
   wire n5879;
   wire n5880;
   wire n5881;
   wire n5882;
   wire n5883;
   wire n5884;
   wire n5885;
   wire n5886;
   wire n5887;
   wire n5888;
   wire n5889;
   wire n5890;
   wire n5891;
   wire n5892;
   wire n5893;
   wire n5894;
   wire n5895;
   wire n5896;
   wire n5897;
   wire n5898;
   wire n5899;
   wire n5900;
   wire n5901;
   wire n5902;
   wire n5903;
   wire n5904;
   wire n5905;
   wire n5906;
   wire n5907;
   wire n5908;
   wire n5909;
   wire n5910;
   wire n5911;
   wire n5912;
   wire n5913;
   wire n5914;
   wire n5915;
   wire n5916;
   wire n5917;
   wire n5918;
   wire n5919;
   wire n5920;
   wire n5921;
   wire n5922;
   wire n5923;
   wire n5924;
   wire n5925;
   wire n5926;
   wire n5927;
   wire n5928;
   wire n5929;
   wire n5930;
   wire n5931;
   wire n5932;
   wire n5933;
   wire n5934;
   wire n5935;
   wire n5936;
   wire n5937;
   wire n5938;
   wire n5939;
   wire n5940;
   wire n5941;
   wire n5942;
   wire n5943;
   wire n5944;
   wire n5945;
   wire n5946;
   wire n5947;
   wire n5948;
   wire n5949;
   wire n5950;
   wire n5951;
   wire n5952;
   wire n5953;
   wire n5954;
   wire n5955;
   wire n5956;
   wire n5957;
   wire n5958;
   wire n5959;
   wire n5960;
   wire n5961;
   wire n5962;
   wire n5963;
   wire n5964;
   wire n5965;
   wire n5966;
   wire n5967;
   wire n5968;
   wire n5969;
   wire n5970;
   wire n5971;
   wire n5972;
   wire n5973;
   wire n5974;
   wire n5975;
   wire n5976;
   wire n5977;
   wire n5978;
   wire n5979;
   wire n5980;
   wire n5981;
   wire n5982;
   wire n5983;
   wire n5984;
   wire n5985;
   wire n5986;
   wire n5987;
   wire n5988;
   wire n5989;
   wire n5990;
   wire n5991;
   wire n5992;
   wire n5993;
   wire n5994;
   wire n5995;
   wire n5996;
   wire n5997;
   wire n5998;
   wire n5999;
   wire n6000;
   wire n6001;
   wire n6002;
   wire n6003;
   wire n6004;
   wire n6005;
   wire n6006;
   wire n6007;
   wire n6008;
   wire n6009;
   wire n6010;
   wire n6011;
   wire n6012;
   wire n6013;
   wire n6014;
   wire n6015;
   wire n6016;
   wire n6038;
   wire n6136;
   wire n6459;
   wire n6469;
   wire n6470;
   wire n6471;
   wire n7439;
   wire n7440;
   wire n7441;
   wire n7442;
   wire n7443;
   wire n7444;
   wire n7445;

   assign N20 = mem_access_addr[2] ;
   assign N21 = mem_access_addr[3] ;
   assign N22 = mem_access_addr[4] ;
   assign N23 = mem_access_addr[5] ;
   assign N24 = mem_access_addr[6] ;
   assign N25 = mem_access_addr[7] ;
   assign N26 = mem_access_addr[8] ;
   assign N27 = mem_access_addr[9] ;

   BUFHHD FE_OFC94_mem_write (.O(FE_OFN94_mem_write), 
	.I(mem_write_en));
   BUFHHD FE_OFC93_mem_write (.O(FE_OFN93_mem_write), 
	.I(mem_write_en));
   BUFHHD FE_OFC92_mem_write (.O(FE_OFN92_mem_write), 
	.I(mem_write_en));
   BUFGHD FE_OFC91_n23 (.O(FE_OFN91_n23), 
	.I(FE_OFN89_n23));
   BUFGHD FE_OFC90_n23 (.O(FE_OFN90_n23), 
	.I(n23));
   BUFGHD FE_OFC89_n23 (.O(FE_OFN89_n23), 
	.I(n23));
   BUFGHD FE_OFC88_n22 (.O(FE_OFN88_n22), 
	.I(n22));
   BUFEHD FE_OFC87_n22 (.O(FE_OFN87_n22), 
	.I(FE_OFN86_n22));
   BUFGHD FE_OFC86_n22 (.O(FE_OFN86_n22), 
	.I(n22));
   BUFGHD FE_OFC85_n21 (.O(FE_OFN85_n21), 
	.I(n21));
   BUFEHD FE_OFC84_n21 (.O(FE_OFN84_n21), 
	.I(FE_OFN83_n21));
   BUFGHD FE_OFC83_n21 (.O(FE_OFN83_n21), 
	.I(n21));
   BUFGHD FE_OFC82_n20 (.O(FE_OFN82_n20), 
	.I(FE_OFN79_n20));
   BUFHHD FE_OFC81_n20 (.O(FE_OFN81_n20), 
	.I(FE_OFN79_n20));
   BUFEHD FE_OFC80_n20 (.O(FE_OFN80_n20), 
	.I(FE_OFN79_n20));
   BUFGHD FE_OFC79_n20 (.O(FE_OFN79_n20), 
	.I(n20));
   BUFGHD FE_OFC78_n19 (.O(FE_OFN78_n19), 
	.I(FE_OFN77_n19));
   BUFGHD FE_OFC77_n19 (.O(FE_OFN77_n19), 
	.I(FE_OFN76_n19));
   BUFGHD FE_OFC76_n19 (.O(FE_OFN76_n19), 
	.I(n19));
   BUFGHD FE_OFC75_n18 (.O(FE_OFN75_n18), 
	.I(FE_OFN74_n18));
   BUFGHD FE_OFC74_n18 (.O(FE_OFN74_n18), 
	.I(FE_OFN73_n18));
   BUFGHD FE_OFC73_n18 (.O(FE_OFN73_n18), 
	.I(n18));
   BUFGHD FE_OFC72_n17 (.O(FE_OFN72_n17), 
	.I(FE_OFN71_n17));
   BUFGHD FE_OFC71_n17 (.O(FE_OFN71_n17), 
	.I(FE_OFN70_n17));
   BUFGHD FE_OFC70_n17 (.O(FE_OFN70_n17), 
	.I(n17));
   BUFGHD FE_OFC69_n16 (.O(FE_OFN69_n16), 
	.I(FE_OFN67_n16));
   BUFGHD FE_OFC68_n16 (.O(FE_OFN68_n16), 
	.I(FE_OFN66_n16));
   BUFGHD FE_OFC67_n16 (.O(FE_OFN67_n16), 
	.I(FE_OFN66_n16));
   BUFGHD FE_OFC66_n16 (.O(FE_OFN66_n16), 
	.I(n16));
   BUFGHD FE_OFC65_n15 (.O(FE_OFN65_n15), 
	.I(FE_OFN64_n15));
   BUFGHD FE_OFC64_n15 (.O(FE_OFN64_n15), 
	.I(FE_OFN63_n15));
   BUFGHD FE_OFC63_n15 (.O(FE_OFN63_n15), 
	.I(n15));
   BUFGHD FE_OFC62_n14 (.O(FE_OFN62_n14), 
	.I(FE_OFN61_n14));
   BUFGHD FE_OFC61_n14 (.O(FE_OFN61_n14), 
	.I(n14));
   BUFEHD FE_OFC60_n14 (.O(FE_OFN60_n14), 
	.I(FE_OFN59_n14));
   BUFGHD FE_OFC59_n14 (.O(FE_OFN59_n14), 
	.I(n14));
   BUFGHD FE_OFC58_n13 (.O(FE_OFN58_n13), 
	.I(FE_OFN57_n13));
   BUFGHD FE_OFC57_n13 (.O(FE_OFN57_n13), 
	.I(FE_OFN56_n13));
   BUFGHD FE_OFC56_n13 (.O(FE_OFN56_n13), 
	.I(n13));
   BUFGHD FE_OFC55_n12 (.O(FE_OFN55_n12), 
	.I(FE_OFN53_n12));
   BUFGHD FE_OFC54_n12 (.O(FE_OFN54_n12), 
	.I(n12));
   BUFGHD FE_OFC53_n12 (.O(FE_OFN53_n12), 
	.I(n12));
   BUFGHD FE_OFC52_n11 (.O(FE_OFN52_n11), 
	.I(FE_OFN51_n11));
   BUFGHD FE_OFC51_n11 (.O(FE_OFN51_n11), 
	.I(FE_OFN50_n11));
   BUFGHD FE_OFC50_n11 (.O(FE_OFN50_n11), 
	.I(n11));
   BUFGHD FE_OFC49_n10 (.O(FE_OFN49_n10), 
	.I(FE_OFN47_n10));
   BUFGHD FE_OFC48_n10 (.O(FE_OFN48_n10), 
	.I(n10));
   BUFGHD FE_OFC47_n10 (.O(FE_OFN47_n10), 
	.I(n10));
   BUFGHD FE_OFC46_n9 (.O(FE_OFN46_n9), 
	.I(FE_OFN44_n9));
   BUFGHD FE_OFC45_n9 (.O(FE_OFN45_n9), 
	.I(n9));
   BUFGHD FE_OFC44_n9 (.O(FE_OFN44_n9), 
	.I(n9));
   BUFGHD FE_OFC43_n6 (.O(FE_OFN43_n6), 
	.I(FE_OFN41_n6));
   BUFHHD FE_OFC42_n6 (.O(FE_OFN42_n6), 
	.I(FE_OFN41_n6));
   BUFGHD FE_OFC41_n6 (.O(FE_OFN41_n6), 
	.I(n6));
   BUFGHD FE_OFC40_n6459 (.O(FE_OFN40_n6459), 
	.I(FE_OFN34_n6459));
   BUFGHD FE_OFC39_n6459 (.O(FE_OFN39_n6459), 
	.I(FE_OFN34_n6459));
   BUFHHD FE_OFC38_n6459 (.O(FE_OFN38_n6459), 
	.I(FE_OFN34_n6459));
   BUFGHD FE_OFC37_n6459 (.O(FE_OFN37_n6459), 
	.I(FE_OFN34_n6459));
   BUFHHD FE_OFC36_n6459 (.O(FE_OFN36_n6459), 
	.I(FE_OFN35_n6459));
   BUFHHD FE_OFC35_n6459 (.O(FE_OFN35_n6459), 
	.I(FE_OFN28_n6459));
   BUFHHD FE_OFC34_n6459 (.O(FE_OFN34_n6459), 
	.I(FE_OFN28_n6459));
   BUFHHD FE_OFC33_n6459 (.O(FE_OFN33_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC32_n6459 (.O(FE_OFN32_n6459), 
	.I(FE_OFN26_n6459));
   BUFHHD FE_OFC31_n6459 (.O(FE_OFN31_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC30_n6459 (.O(FE_OFN30_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC29_n6459 (.O(FE_OFN29_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC28_n6459 (.O(FE_OFN28_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC27_n6459 (.O(FE_OFN27_n6459), 
	.I(FE_OFN26_n6459));
   BUFHHD FE_OFC26_n6459 (.O(FE_OFN26_n6459), 
	.I(FE_OFN25_n6459));
   BUFGHD FE_OFC25_n6459 (.O(FE_OFN25_n6459), 
	.I(n6459));
   BUFHHD FE_OFC24_n6136 (.O(FE_OFN24_n6136), 
	.I(FE_OFN23_n6136));
   BUFHHD FE_OFC23_n6136 (.O(FE_OFN23_n6136), 
	.I(n6136));
   BUFHHD FE_OFC22_n6136 (.O(FE_OFN22_n6136), 
	.I(n6136));
   BUFGHD FE_OFC21_n7440 (.O(FE_OFN21_n7440), 
	.I(FE_OFN9_n7440));
   BUFHHD FE_OFC20_n7440 (.O(FE_OFN20_n7440), 
	.I(FE_OFN9_n7440));
   BUFJHD FE_OFC19_n7440 (.O(FE_OFN19_n7440), 
	.I(FE_OFN14_n7440));
   BUFHHD FE_OFC18_n7440 (.O(FE_OFN18_n7440), 
	.I(FE_OFN9_n7440));
   BUFIHD FE_OFC17_n7440 (.O(FE_OFN17_n7440), 
	.I(n7440));
   BUFIHD FE_OFC16_n7440 (.O(FE_OFN16_n7440), 
	.I(n7440));
   BUFHHD FE_OFC15_n7440 (.O(FE_OFN15_n7440), 
	.I(FE_OFN10_n7440));
   BUFHHD FE_OFC14_n7440 (.O(FE_OFN14_n7440), 
	.I(FE_OFN9_n7440));
   BUFJHD FE_OFC13_n7440 (.O(FE_OFN13_n7440), 
	.I(FE_OFN11_n7440));
   BUFHHD FE_OFC12_n7440 (.O(FE_OFN12_n7440), 
	.I(n7440));
   BUFHHD FE_OFC11_n7440 (.O(FE_OFN11_n7440), 
	.I(FE_OFN7_n7440));
   BUFJHD FE_OFC10_n7440 (.O(FE_OFN10_n7440), 
	.I(n7440));
   BUFGHD FE_OFC9_n7440 (.O(FE_OFN9_n7440), 
	.I(n7440));
   BUFJHD FE_OFC8_n7440 (.O(FE_OFN8_n7440), 
	.I(FE_OFN6_n7440));
   BUFIHD FE_OFC7_n7440 (.O(FE_OFN7_n7440), 
	.I(n7440));
   BUFIHD FE_OFC6_n7440 (.O(FE_OFN6_n7440), 
	.I(n7440));
   BUFHHD FE_OFC5_n7440 (.O(FE_OFN5_n7440), 
	.I(n7440));
   BUFGHD FE_OFC4_n7442 (.O(FE_OFN4_n7442), 
	.I(FE_OFN2_n7442));
   BUFGHD FE_OFC3_n7442 (.O(FE_OFN3_n7442), 
	.I(FE_OFN0_n7442));
   BUFJHD FE_OFC2_n7442 (.O(FE_OFN2_n7442), 
	.I(n7442));
   BUFGHD FE_OFC1_n7442 (.O(FE_OFN1_n7442), 
	.I(n7442));
   BUFGHD FE_OFC0_n7442 (.O(FE_OFN0_n7442), 
	.I(n7442));
   QDFFEHD \ram_reg[253][15]  (.Q(\ram[253][15] ), 
	.D(n4645), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[253][14]  (.Q(\ram[253][14] ), 
	.D(n4644), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[253][13]  (.Q(\ram[253][13] ), 
	.D(n4643), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[253][12]  (.Q(\ram[253][12] ), 
	.D(n4642), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[253][11]  (.Q(\ram[253][11] ), 
	.D(n4641), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[253][10]  (.Q(\ram[253][10] ), 
	.D(n4640), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][9]  (.Q(\ram[253][9] ), 
	.D(n4639), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][8]  (.Q(\ram[253][8] ), 
	.D(n4638), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][7]  (.Q(\ram[253][7] ), 
	.D(n4637), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[253][6]  (.Q(\ram[253][6] ), 
	.D(n4636), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[253][5]  (.Q(\ram[253][5] ), 
	.D(n4635), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[253][4]  (.Q(\ram[253][4] ), 
	.D(n4634), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[253][3]  (.Q(\ram[253][3] ), 
	.D(n4633), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][2]  (.Q(\ram[253][2] ), 
	.D(n4632), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[253][1]  (.Q(\ram[253][1] ), 
	.D(n4631), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[253][0]  (.Q(\ram[253][0] ), 
	.D(n4630), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[249][15]  (.Q(\ram[249][15] ), 
	.D(n4581), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][14]  (.Q(\ram[249][14] ), 
	.D(n4580), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[249][13]  (.Q(\ram[249][13] ), 
	.D(n4579), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[249][12]  (.Q(\ram[249][12] ), 
	.D(n4578), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][11]  (.Q(\ram[249][11] ), 
	.D(n4577), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][10]  (.Q(\ram[249][10] ), 
	.D(n4576), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][9]  (.Q(\ram[249][9] ), 
	.D(n4575), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][8]  (.Q(\ram[249][8] ), 
	.D(n4574), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[249][7]  (.Q(\ram[249][7] ), 
	.D(n4573), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][6]  (.Q(\ram[249][6] ), 
	.D(n4572), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][5]  (.Q(\ram[249][5] ), 
	.D(n4571), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][4]  (.Q(\ram[249][4] ), 
	.D(n4570), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][3]  (.Q(\ram[249][3] ), 
	.D(n4569), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[249][2]  (.Q(\ram[249][2] ), 
	.D(n4568), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][1]  (.Q(\ram[249][1] ), 
	.D(n4567), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[249][0]  (.Q(\ram[249][0] ), 
	.D(n4566), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[245][15]  (.Q(\ram[245][15] ), 
	.D(n4517), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][14]  (.Q(\ram[245][14] ), 
	.D(n4516), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][13]  (.Q(\ram[245][13] ), 
	.D(n4515), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][12]  (.Q(\ram[245][12] ), 
	.D(n4514), 
	.CK(clk));
   QDFFEHD \ram_reg[245][11]  (.Q(\ram[245][11] ), 
	.D(n4513), 
	.CK(clk));
   QDFFEHD \ram_reg[245][10]  (.Q(\ram[245][10] ), 
	.D(n4512), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][9]  (.Q(\ram[245][9] ), 
	.D(n4511), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[245][8]  (.Q(\ram[245][8] ), 
	.D(n4510), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[245][7]  (.Q(\ram[245][7] ), 
	.D(n4509), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][6]  (.Q(\ram[245][6] ), 
	.D(n4508), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][5]  (.Q(\ram[245][5] ), 
	.D(n4507), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][4]  (.Q(\ram[245][4] ), 
	.D(n4506), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][3]  (.Q(\ram[245][3] ), 
	.D(n4505), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[245][2]  (.Q(\ram[245][2] ), 
	.D(n4504), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][1]  (.Q(\ram[245][1] ), 
	.D(n4503), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][0]  (.Q(\ram[245][0] ), 
	.D(n4502), 
	.CK(clk));
   QDFFEHD \ram_reg[241][15]  (.Q(\ram[241][15] ), 
	.D(n4453), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[241][14]  (.Q(\ram[241][14] ), 
	.D(n4452), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][13]  (.Q(\ram[241][13] ), 
	.D(n4451), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][12]  (.Q(\ram[241][12] ), 
	.D(n4450), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][11]  (.Q(\ram[241][11] ), 
	.D(n4449), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][10]  (.Q(\ram[241][10] ), 
	.D(n4448), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][9]  (.Q(\ram[241][9] ), 
	.D(n4447), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][8]  (.Q(\ram[241][8] ), 
	.D(n4446), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][7]  (.Q(\ram[241][7] ), 
	.D(n4445), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][6]  (.Q(\ram[241][6] ), 
	.D(n4444), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][5]  (.Q(\ram[241][5] ), 
	.D(n4443), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][4]  (.Q(\ram[241][4] ), 
	.D(n4442), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][3]  (.Q(\ram[241][3] ), 
	.D(n4441), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][2]  (.Q(\ram[241][2] ), 
	.D(n4440), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][1]  (.Q(\ram[241][1] ), 
	.D(n4439), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][0]  (.Q(\ram[241][0] ), 
	.D(n4438), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[237][15]  (.Q(\ram[237][15] ), 
	.D(n4389), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][14]  (.Q(\ram[237][14] ), 
	.D(n4388), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][13]  (.Q(\ram[237][13] ), 
	.D(n4387), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][12]  (.Q(\ram[237][12] ), 
	.D(n4386), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][11]  (.Q(\ram[237][11] ), 
	.D(n4385), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][10]  (.Q(\ram[237][10] ), 
	.D(n4384), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][9]  (.Q(\ram[237][9] ), 
	.D(n4383), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][8]  (.Q(\ram[237][8] ), 
	.D(n4382), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][7]  (.Q(\ram[237][7] ), 
	.D(n4381), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][6]  (.Q(\ram[237][6] ), 
	.D(n4380), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][5]  (.Q(\ram[237][5] ), 
	.D(n4379), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[237][4]  (.Q(\ram[237][4] ), 
	.D(n4378), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][3]  (.Q(\ram[237][3] ), 
	.D(n4377), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][2]  (.Q(\ram[237][2] ), 
	.D(n4376), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][1]  (.Q(\ram[237][1] ), 
	.D(n4375), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][0]  (.Q(\ram[237][0] ), 
	.D(n4374), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[233][15]  (.Q(\ram[233][15] ), 
	.D(n4325), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[233][14]  (.Q(\ram[233][14] ), 
	.D(n4324), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[233][13]  (.Q(\ram[233][13] ), 
	.D(n4323), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[233][12]  (.Q(\ram[233][12] ), 
	.D(n4322), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[233][11]  (.Q(\ram[233][11] ), 
	.D(n4321), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[233][10]  (.Q(\ram[233][10] ), 
	.D(n4320), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][9]  (.Q(\ram[233][9] ), 
	.D(n4319), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][8]  (.Q(\ram[233][8] ), 
	.D(n4318), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][7]  (.Q(\ram[233][7] ), 
	.D(n4317), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[233][6]  (.Q(\ram[233][6] ), 
	.D(n4316), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][5]  (.Q(\ram[233][5] ), 
	.D(n4315), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[233][4]  (.Q(\ram[233][4] ), 
	.D(n4314), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][3]  (.Q(\ram[233][3] ), 
	.D(n4313), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[233][2]  (.Q(\ram[233][2] ), 
	.D(n4312), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][1]  (.Q(\ram[233][1] ), 
	.D(n4311), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[233][0]  (.Q(\ram[233][0] ), 
	.D(n4310), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[229][15]  (.Q(\ram[229][15] ), 
	.D(n4261), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][14]  (.Q(\ram[229][14] ), 
	.D(n4260), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[229][13]  (.Q(\ram[229][13] ), 
	.D(n4259), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[229][12]  (.Q(\ram[229][12] ), 
	.D(n4258), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[229][11]  (.Q(\ram[229][11] ), 
	.D(n4257), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][10]  (.Q(\ram[229][10] ), 
	.D(n4256), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][9]  (.Q(\ram[229][9] ), 
	.D(n4255), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[229][8]  (.Q(\ram[229][8] ), 
	.D(n4254), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][7]  (.Q(\ram[229][7] ), 
	.D(n4253), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][6]  (.Q(\ram[229][6] ), 
	.D(n4252), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[229][5]  (.Q(\ram[229][5] ), 
	.D(n4251), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[229][4]  (.Q(\ram[229][4] ), 
	.D(n4250), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[229][3]  (.Q(\ram[229][3] ), 
	.D(n4249), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[229][2]  (.Q(\ram[229][2] ), 
	.D(n4248), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[229][1]  (.Q(\ram[229][1] ), 
	.D(n4247), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[229][0]  (.Q(\ram[229][0] ), 
	.D(n4246), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[225][15]  (.Q(\ram[225][15] ), 
	.D(n4197), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[225][14]  (.Q(\ram[225][14] ), 
	.D(n4196), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][13]  (.Q(\ram[225][13] ), 
	.D(n4195), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[225][12]  (.Q(\ram[225][12] ), 
	.D(n4194), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][11]  (.Q(\ram[225][11] ), 
	.D(n4193), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[225][10]  (.Q(\ram[225][10] ), 
	.D(n4192), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[225][9]  (.Q(\ram[225][9] ), 
	.D(n4191), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[225][8]  (.Q(\ram[225][8] ), 
	.D(n4190), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[225][7]  (.Q(\ram[225][7] ), 
	.D(n4189), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[225][6]  (.Q(\ram[225][6] ), 
	.D(n4188), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][5]  (.Q(\ram[225][5] ), 
	.D(n4187), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[225][4]  (.Q(\ram[225][4] ), 
	.D(n4186), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[225][3]  (.Q(\ram[225][3] ), 
	.D(n4185), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][2]  (.Q(\ram[225][2] ), 
	.D(n4184), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[225][1]  (.Q(\ram[225][1] ), 
	.D(n4183), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][0]  (.Q(\ram[225][0] ), 
	.D(n4182), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[221][15]  (.Q(\ram[221][15] ), 
	.D(n4133), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][14]  (.Q(\ram[221][14] ), 
	.D(n4132), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][13]  (.Q(\ram[221][13] ), 
	.D(n4131), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][12]  (.Q(\ram[221][12] ), 
	.D(n4130), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][11]  (.Q(\ram[221][11] ), 
	.D(n4129), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][10]  (.Q(\ram[221][10] ), 
	.D(n4128), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[221][9]  (.Q(\ram[221][9] ), 
	.D(n4127), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][8]  (.Q(\ram[221][8] ), 
	.D(n4126), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][7]  (.Q(\ram[221][7] ), 
	.D(n4125), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[221][6]  (.Q(\ram[221][6] ), 
	.D(n4124), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[221][5]  (.Q(\ram[221][5] ), 
	.D(n4123), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][4]  (.Q(\ram[221][4] ), 
	.D(n4122), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][3]  (.Q(\ram[221][3] ), 
	.D(n4121), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[221][2]  (.Q(\ram[221][2] ), 
	.D(n4120), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][1]  (.Q(\ram[221][1] ), 
	.D(n4119), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[221][0]  (.Q(\ram[221][0] ), 
	.D(n4118), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[217][15]  (.Q(\ram[217][15] ), 
	.D(n4069), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][14]  (.Q(\ram[217][14] ), 
	.D(n4068), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][13]  (.Q(\ram[217][13] ), 
	.D(n4067), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][12]  (.Q(\ram[217][12] ), 
	.D(n4066), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][11]  (.Q(\ram[217][11] ), 
	.D(n4065), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[217][10]  (.Q(\ram[217][10] ), 
	.D(n4064), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][9]  (.Q(\ram[217][9] ), 
	.D(n4063), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][8]  (.Q(\ram[217][8] ), 
	.D(n4062), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][7]  (.Q(\ram[217][7] ), 
	.D(n4061), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][6]  (.Q(\ram[217][6] ), 
	.D(n4060), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][5]  (.Q(\ram[217][5] ), 
	.D(n4059), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][4]  (.Q(\ram[217][4] ), 
	.D(n4058), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[217][3]  (.Q(\ram[217][3] ), 
	.D(n4057), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[217][2]  (.Q(\ram[217][2] ), 
	.D(n4056), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[217][1]  (.Q(\ram[217][1] ), 
	.D(n4055), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[217][0]  (.Q(\ram[217][0] ), 
	.D(n4054), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[213][15]  (.Q(\ram[213][15] ), 
	.D(n4005), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[213][14]  (.Q(\ram[213][14] ), 
	.D(n4004), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][13]  (.Q(\ram[213][13] ), 
	.D(n4003), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[213][12]  (.Q(\ram[213][12] ), 
	.D(n4002), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[213][11]  (.Q(\ram[213][11] ), 
	.D(n4001), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][10]  (.Q(\ram[213][10] ), 
	.D(n4000), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][9]  (.Q(\ram[213][9] ), 
	.D(n3999), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[213][8]  (.Q(\ram[213][8] ), 
	.D(n3998), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[213][7]  (.Q(\ram[213][7] ), 
	.D(n3997), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][6]  (.Q(\ram[213][6] ), 
	.D(n3996), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][5]  (.Q(\ram[213][5] ), 
	.D(n3995), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[213][4]  (.Q(\ram[213][4] ), 
	.D(n3994), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][3]  (.Q(\ram[213][3] ), 
	.D(n3993), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[213][2]  (.Q(\ram[213][2] ), 
	.D(n3992), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][1]  (.Q(\ram[213][1] ), 
	.D(n3991), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[213][0]  (.Q(\ram[213][0] ), 
	.D(n3990), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[209][15]  (.Q(\ram[209][15] ), 
	.D(n3941), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[209][14]  (.Q(\ram[209][14] ), 
	.D(n3940), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[209][13]  (.Q(\ram[209][13] ), 
	.D(n3939), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][12]  (.Q(\ram[209][12] ), 
	.D(n3938), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][11]  (.Q(\ram[209][11] ), 
	.D(n3937), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][10]  (.Q(\ram[209][10] ), 
	.D(n3936), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][9]  (.Q(\ram[209][9] ), 
	.D(n3935), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][8]  (.Q(\ram[209][8] ), 
	.D(n3934), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][7]  (.Q(\ram[209][7] ), 
	.D(n3933), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][6]  (.Q(\ram[209][6] ), 
	.D(n3932), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[209][5]  (.Q(\ram[209][5] ), 
	.D(n3931), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][4]  (.Q(\ram[209][4] ), 
	.D(n3930), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[209][3]  (.Q(\ram[209][3] ), 
	.D(n3929), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[209][2]  (.Q(\ram[209][2] ), 
	.D(n3928), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[209][1]  (.Q(\ram[209][1] ), 
	.D(n3927), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[209][0]  (.Q(\ram[209][0] ), 
	.D(n3926), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[205][15]  (.Q(\ram[205][15] ), 
	.D(n3877), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][14]  (.Q(\ram[205][14] ), 
	.D(n3876), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][13]  (.Q(\ram[205][13] ), 
	.D(n3875), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[205][12]  (.Q(\ram[205][12] ), 
	.D(n3874), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][11]  (.Q(\ram[205][11] ), 
	.D(n3873), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][10]  (.Q(\ram[205][10] ), 
	.D(n3872), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][9]  (.Q(\ram[205][9] ), 
	.D(n3871), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][8]  (.Q(\ram[205][8] ), 
	.D(n3870), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[205][7]  (.Q(\ram[205][7] ), 
	.D(n3869), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][6]  (.Q(\ram[205][6] ), 
	.D(n3868), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][5]  (.Q(\ram[205][5] ), 
	.D(n3867), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][4]  (.Q(\ram[205][4] ), 
	.D(n3866), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][3]  (.Q(\ram[205][3] ), 
	.D(n3865), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][2]  (.Q(\ram[205][2] ), 
	.D(n3864), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][1]  (.Q(\ram[205][1] ), 
	.D(n3863), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][0]  (.Q(\ram[205][0] ), 
	.D(n3862), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[201][15]  (.Q(\ram[201][15] ), 
	.D(n3813), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][14]  (.Q(\ram[201][14] ), 
	.D(n3812), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][13]  (.Q(\ram[201][13] ), 
	.D(n3811), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[201][12]  (.Q(\ram[201][12] ), 
	.D(n3810), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][11]  (.Q(\ram[201][11] ), 
	.D(n3809), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][10]  (.Q(\ram[201][10] ), 
	.D(n3808), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][9]  (.Q(\ram[201][9] ), 
	.D(n3807), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[201][8]  (.Q(\ram[201][8] ), 
	.D(n3806), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[201][7]  (.Q(\ram[201][7] ), 
	.D(n3805), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][6]  (.Q(\ram[201][6] ), 
	.D(n3804), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[201][5]  (.Q(\ram[201][5] ), 
	.D(n3803), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[201][4]  (.Q(\ram[201][4] ), 
	.D(n3802), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[201][3]  (.Q(\ram[201][3] ), 
	.D(n3801), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[201][2]  (.Q(\ram[201][2] ), 
	.D(n3800), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][1]  (.Q(\ram[201][1] ), 
	.D(n3799), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][0]  (.Q(\ram[201][0] ), 
	.D(n3798), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[197][15]  (.Q(\ram[197][15] ), 
	.D(n3749), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][14]  (.Q(\ram[197][14] ), 
	.D(n3748), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][13]  (.Q(\ram[197][13] ), 
	.D(n3747), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[197][12]  (.Q(\ram[197][12] ), 
	.D(n3746), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[197][11]  (.Q(\ram[197][11] ), 
	.D(n3745), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][10]  (.Q(\ram[197][10] ), 
	.D(n3744), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][9]  (.Q(\ram[197][9] ), 
	.D(n3743), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[197][8]  (.Q(\ram[197][8] ), 
	.D(n3742), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][7]  (.Q(\ram[197][7] ), 
	.D(n3741), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][6]  (.Q(\ram[197][6] ), 
	.D(n3740), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][5]  (.Q(\ram[197][5] ), 
	.D(n3739), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][4]  (.Q(\ram[197][4] ), 
	.D(n3738), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][3]  (.Q(\ram[197][3] ), 
	.D(n3737), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[197][2]  (.Q(\ram[197][2] ), 
	.D(n3736), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][1]  (.Q(\ram[197][1] ), 
	.D(n3735), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][0]  (.Q(\ram[197][0] ), 
	.D(n3734), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[193][15]  (.Q(\ram[193][15] ), 
	.D(n3685), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][14]  (.Q(\ram[193][14] ), 
	.D(n3684), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][13]  (.Q(\ram[193][13] ), 
	.D(n3683), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[193][12]  (.Q(\ram[193][12] ), 
	.D(n3682), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][11]  (.Q(\ram[193][11] ), 
	.D(n3681), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][10]  (.Q(\ram[193][10] ), 
	.D(n3680), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[193][9]  (.Q(\ram[193][9] ), 
	.D(n3679), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][8]  (.Q(\ram[193][8] ), 
	.D(n3678), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[193][7]  (.Q(\ram[193][7] ), 
	.D(n3677), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[193][6]  (.Q(\ram[193][6] ), 
	.D(n3676), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][5]  (.Q(\ram[193][5] ), 
	.D(n3675), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][4]  (.Q(\ram[193][4] ), 
	.D(n3674), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][3]  (.Q(\ram[193][3] ), 
	.D(n3673), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][2]  (.Q(\ram[193][2] ), 
	.D(n3672), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][1]  (.Q(\ram[193][1] ), 
	.D(n3671), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[193][0]  (.Q(\ram[193][0] ), 
	.D(n3670), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[189][15]  (.Q(\ram[189][15] ), 
	.D(n3621), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][14]  (.Q(\ram[189][14] ), 
	.D(n3620), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[189][13]  (.Q(\ram[189][13] ), 
	.D(n3619), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[189][12]  (.Q(\ram[189][12] ), 
	.D(n3618), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[189][11]  (.Q(\ram[189][11] ), 
	.D(n3617), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[189][10]  (.Q(\ram[189][10] ), 
	.D(n3616), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[189][9]  (.Q(\ram[189][9] ), 
	.D(n3615), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[189][8]  (.Q(\ram[189][8] ), 
	.D(n3614), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][7]  (.Q(\ram[189][7] ), 
	.D(n3613), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][6]  (.Q(\ram[189][6] ), 
	.D(n3612), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[189][5]  (.Q(\ram[189][5] ), 
	.D(n3611), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[189][4]  (.Q(\ram[189][4] ), 
	.D(n3610), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][3]  (.Q(\ram[189][3] ), 
	.D(n3609), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[189][2]  (.Q(\ram[189][2] ), 
	.D(n3608), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[189][1]  (.Q(\ram[189][1] ), 
	.D(n3607), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][0]  (.Q(\ram[189][0] ), 
	.D(n3606), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[185][15]  (.Q(\ram[185][15] ), 
	.D(n3557), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][14]  (.Q(\ram[185][14] ), 
	.D(n3556), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][13]  (.Q(\ram[185][13] ), 
	.D(n3555), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][12]  (.Q(\ram[185][12] ), 
	.D(n3554), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[185][11]  (.Q(\ram[185][11] ), 
	.D(n3553), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][10]  (.Q(\ram[185][10] ), 
	.D(n3552), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[185][9]  (.Q(\ram[185][9] ), 
	.D(n3551), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[185][8]  (.Q(\ram[185][8] ), 
	.D(n3550), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][7]  (.Q(\ram[185][7] ), 
	.D(n3549), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][6]  (.Q(\ram[185][6] ), 
	.D(n3548), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][5]  (.Q(\ram[185][5] ), 
	.D(n3547), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][4]  (.Q(\ram[185][4] ), 
	.D(n3546), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[185][3]  (.Q(\ram[185][3] ), 
	.D(n3545), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][2]  (.Q(\ram[185][2] ), 
	.D(n3544), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][1]  (.Q(\ram[185][1] ), 
	.D(n3543), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][0]  (.Q(\ram[185][0] ), 
	.D(n3542), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[181][15]  (.Q(\ram[181][15] ), 
	.D(n3493), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[181][14]  (.Q(\ram[181][14] ), 
	.D(n3492), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[181][13]  (.Q(\ram[181][13] ), 
	.D(n3491), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[181][12]  (.Q(\ram[181][12] ), 
	.D(n3490), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[181][11]  (.Q(\ram[181][11] ), 
	.D(n3489), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[181][10]  (.Q(\ram[181][10] ), 
	.D(n3488), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][9]  (.Q(\ram[181][9] ), 
	.D(n3487), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][8]  (.Q(\ram[181][8] ), 
	.D(n3486), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][7]  (.Q(\ram[181][7] ), 
	.D(n3485), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[181][6]  (.Q(\ram[181][6] ), 
	.D(n3484), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][5]  (.Q(\ram[181][5] ), 
	.D(n3483), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[181][4]  (.Q(\ram[181][4] ), 
	.D(n3482), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[181][3]  (.Q(\ram[181][3] ), 
	.D(n3481), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[181][2]  (.Q(\ram[181][2] ), 
	.D(n3480), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[181][1]  (.Q(\ram[181][1] ), 
	.D(n3479), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[181][0]  (.Q(\ram[181][0] ), 
	.D(n3478), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[177][15]  (.Q(\ram[177][15] ), 
	.D(n3429), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[177][14]  (.Q(\ram[177][14] ), 
	.D(n3428), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][13]  (.Q(\ram[177][13] ), 
	.D(n3427), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[177][12]  (.Q(\ram[177][12] ), 
	.D(n3426), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[177][11]  (.Q(\ram[177][11] ), 
	.D(n3425), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[177][10]  (.Q(\ram[177][10] ), 
	.D(n3424), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[177][9]  (.Q(\ram[177][9] ), 
	.D(n3423), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][8]  (.Q(\ram[177][8] ), 
	.D(n3422), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[177][7]  (.Q(\ram[177][7] ), 
	.D(n3421), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][6]  (.Q(\ram[177][6] ), 
	.D(n3420), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[177][5]  (.Q(\ram[177][5] ), 
	.D(n3419), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[177][4]  (.Q(\ram[177][4] ), 
	.D(n3418), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][3]  (.Q(\ram[177][3] ), 
	.D(n3417), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[177][2]  (.Q(\ram[177][2] ), 
	.D(n3416), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][1]  (.Q(\ram[177][1] ), 
	.D(n3415), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][0]  (.Q(\ram[177][0] ), 
	.D(n3414), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[173][15]  (.Q(\ram[173][15] ), 
	.D(n3365), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][14]  (.Q(\ram[173][14] ), 
	.D(n3364), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][13]  (.Q(\ram[173][13] ), 
	.D(n3363), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[173][12]  (.Q(\ram[173][12] ), 
	.D(n3362), 
	.CK(clk));
   QDFFEHD \ram_reg[173][11]  (.Q(\ram[173][11] ), 
	.D(n3361), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[173][10]  (.Q(\ram[173][10] ), 
	.D(n3360), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[173][9]  (.Q(\ram[173][9] ), 
	.D(n3359), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][8]  (.Q(\ram[173][8] ), 
	.D(n3358), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[173][7]  (.Q(\ram[173][7] ), 
	.D(n3357), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][6]  (.Q(\ram[173][6] ), 
	.D(n3356), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][5]  (.Q(\ram[173][5] ), 
	.D(n3355), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][4]  (.Q(\ram[173][4] ), 
	.D(n3354), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][3]  (.Q(\ram[173][3] ), 
	.D(n3353), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][2]  (.Q(\ram[173][2] ), 
	.D(n3352), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][1]  (.Q(\ram[173][1] ), 
	.D(n3351), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][0]  (.Q(\ram[173][0] ), 
	.D(n3350), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[169][15]  (.Q(\ram[169][15] ), 
	.D(n3301), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][14]  (.Q(\ram[169][14] ), 
	.D(n3300), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][13]  (.Q(\ram[169][13] ), 
	.D(n3299), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][12]  (.Q(\ram[169][12] ), 
	.D(n3298), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][11]  (.Q(\ram[169][11] ), 
	.D(n3297), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][10]  (.Q(\ram[169][10] ), 
	.D(n3296), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][9]  (.Q(\ram[169][9] ), 
	.D(n3295), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][8]  (.Q(\ram[169][8] ), 
	.D(n3294), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[169][7]  (.Q(\ram[169][7] ), 
	.D(n3293), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][6]  (.Q(\ram[169][6] ), 
	.D(n3292), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][5]  (.Q(\ram[169][5] ), 
	.D(n3291), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][4]  (.Q(\ram[169][4] ), 
	.D(n3290), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][3]  (.Q(\ram[169][3] ), 
	.D(n3289), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][2]  (.Q(\ram[169][2] ), 
	.D(n3288), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][1]  (.Q(\ram[169][1] ), 
	.D(n3287), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[169][0]  (.Q(\ram[169][0] ), 
	.D(n3286), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[165][15]  (.Q(\ram[165][15] ), 
	.D(n3237), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[165][14]  (.Q(\ram[165][14] ), 
	.D(n3236), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[165][13]  (.Q(\ram[165][13] ), 
	.D(n3235), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[165][12]  (.Q(\ram[165][12] ), 
	.D(n3234), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[165][11]  (.Q(\ram[165][11] ), 
	.D(n3233), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][10]  (.Q(\ram[165][10] ), 
	.D(n3232), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][9]  (.Q(\ram[165][9] ), 
	.D(n3231), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][8]  (.Q(\ram[165][8] ), 
	.D(n3230), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][7]  (.Q(\ram[165][7] ), 
	.D(n3229), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][6]  (.Q(\ram[165][6] ), 
	.D(n3228), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][5]  (.Q(\ram[165][5] ), 
	.D(n3227), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][4]  (.Q(\ram[165][4] ), 
	.D(n3226), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][3]  (.Q(\ram[165][3] ), 
	.D(n3225), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][2]  (.Q(\ram[165][2] ), 
	.D(n3224), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[165][1]  (.Q(\ram[165][1] ), 
	.D(n3223), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][0]  (.Q(\ram[165][0] ), 
	.D(n3222), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[161][15]  (.Q(\ram[161][15] ), 
	.D(n3173), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][14]  (.Q(\ram[161][14] ), 
	.D(n3172), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][13]  (.Q(\ram[161][13] ), 
	.D(n3171), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][12]  (.Q(\ram[161][12] ), 
	.D(n3170), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[161][11]  (.Q(\ram[161][11] ), 
	.D(n3169), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[161][10]  (.Q(\ram[161][10] ), 
	.D(n3168), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[161][9]  (.Q(\ram[161][9] ), 
	.D(n3167), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[161][8]  (.Q(\ram[161][8] ), 
	.D(n3166), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[161][7]  (.Q(\ram[161][7] ), 
	.D(n3165), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][6]  (.Q(\ram[161][6] ), 
	.D(n3164), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][5]  (.Q(\ram[161][5] ), 
	.D(n3163), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][4]  (.Q(\ram[161][4] ), 
	.D(n3162), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][3]  (.Q(\ram[161][3] ), 
	.D(n3161), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][2]  (.Q(\ram[161][2] ), 
	.D(n3160), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[161][1]  (.Q(\ram[161][1] ), 
	.D(n3159), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][0]  (.Q(\ram[161][0] ), 
	.D(n3158), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[157][15]  (.Q(\ram[157][15] ), 
	.D(n3109), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[157][14]  (.Q(\ram[157][14] ), 
	.D(n3108), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][13]  (.Q(\ram[157][13] ), 
	.D(n3107), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][12]  (.Q(\ram[157][12] ), 
	.D(n3106), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][11]  (.Q(\ram[157][11] ), 
	.D(n3105), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][10]  (.Q(\ram[157][10] ), 
	.D(n3104), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][9]  (.Q(\ram[157][9] ), 
	.D(n3103), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[157][8]  (.Q(\ram[157][8] ), 
	.D(n3102), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[157][7]  (.Q(\ram[157][7] ), 
	.D(n3101), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[157][6]  (.Q(\ram[157][6] ), 
	.D(n3100), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[157][5]  (.Q(\ram[157][5] ), 
	.D(n3099), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[157][4]  (.Q(\ram[157][4] ), 
	.D(n3098), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[157][3]  (.Q(\ram[157][3] ), 
	.D(n3097), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[157][2]  (.Q(\ram[157][2] ), 
	.D(n3096), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[157][1]  (.Q(\ram[157][1] ), 
	.D(n3095), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[157][0]  (.Q(\ram[157][0] ), 
	.D(n3094), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[153][15]  (.Q(\ram[153][15] ), 
	.D(n3045), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[153][14]  (.Q(\ram[153][14] ), 
	.D(n3044), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][13]  (.Q(\ram[153][13] ), 
	.D(n3043), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][12]  (.Q(\ram[153][12] ), 
	.D(n3042), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[153][11]  (.Q(\ram[153][11] ), 
	.D(n3041), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][10]  (.Q(\ram[153][10] ), 
	.D(n3040), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][9]  (.Q(\ram[153][9] ), 
	.D(n3039), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[153][8]  (.Q(\ram[153][8] ), 
	.D(n3038), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[153][7]  (.Q(\ram[153][7] ), 
	.D(n3037), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][6]  (.Q(\ram[153][6] ), 
	.D(n3036), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[153][5]  (.Q(\ram[153][5] ), 
	.D(n3035), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[153][4]  (.Q(\ram[153][4] ), 
	.D(n3034), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[153][3]  (.Q(\ram[153][3] ), 
	.D(n3033), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][2]  (.Q(\ram[153][2] ), 
	.D(n3032), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][1]  (.Q(\ram[153][1] ), 
	.D(n3031), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][0]  (.Q(\ram[153][0] ), 
	.D(n3030), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[149][15]  (.Q(\ram[149][15] ), 
	.D(n2981), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][14]  (.Q(\ram[149][14] ), 
	.D(n2980), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][13]  (.Q(\ram[149][13] ), 
	.D(n2979), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][12]  (.Q(\ram[149][12] ), 
	.D(n2978), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][11]  (.Q(\ram[149][11] ), 
	.D(n2977), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][10]  (.Q(\ram[149][10] ), 
	.D(n2976), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[149][9]  (.Q(\ram[149][9] ), 
	.D(n2975), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[149][8]  (.Q(\ram[149][8] ), 
	.D(n2974), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[149][7]  (.Q(\ram[149][7] ), 
	.D(n2973), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][6]  (.Q(\ram[149][6] ), 
	.D(n2972), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][5]  (.Q(\ram[149][5] ), 
	.D(n2971), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][4]  (.Q(\ram[149][4] ), 
	.D(n2970), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][3]  (.Q(\ram[149][3] ), 
	.D(n2969), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][2]  (.Q(\ram[149][2] ), 
	.D(n2968), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[149][1]  (.Q(\ram[149][1] ), 
	.D(n2967), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][0]  (.Q(\ram[149][0] ), 
	.D(n2966), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[145][15]  (.Q(\ram[145][15] ), 
	.D(n2917), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[145][14]  (.Q(\ram[145][14] ), 
	.D(n2916), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][13]  (.Q(\ram[145][13] ), 
	.D(n2915), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[145][12]  (.Q(\ram[145][12] ), 
	.D(n2914), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][11]  (.Q(\ram[145][11] ), 
	.D(n2913), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[145][10]  (.Q(\ram[145][10] ), 
	.D(n2912), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[145][9]  (.Q(\ram[145][9] ), 
	.D(n2911), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][8]  (.Q(\ram[145][8] ), 
	.D(n2910), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][7]  (.Q(\ram[145][7] ), 
	.D(n2909), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][6]  (.Q(\ram[145][6] ), 
	.D(n2908), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][5]  (.Q(\ram[145][5] ), 
	.D(n2907), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][4]  (.Q(\ram[145][4] ), 
	.D(n2906), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][3]  (.Q(\ram[145][3] ), 
	.D(n2905), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][2]  (.Q(\ram[145][2] ), 
	.D(n2904), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[145][1]  (.Q(\ram[145][1] ), 
	.D(n2903), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][0]  (.Q(\ram[145][0] ), 
	.D(n2902), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[141][15]  (.Q(\ram[141][15] ), 
	.D(n2853), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[141][14]  (.Q(\ram[141][14] ), 
	.D(n2852), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][13]  (.Q(\ram[141][13] ), 
	.D(n2851), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][12]  (.Q(\ram[141][12] ), 
	.D(n2850), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[141][11]  (.Q(\ram[141][11] ), 
	.D(n2849), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[141][10]  (.Q(\ram[141][10] ), 
	.D(n2848), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[141][9]  (.Q(\ram[141][9] ), 
	.D(n2847), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][8]  (.Q(\ram[141][8] ), 
	.D(n2846), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][7]  (.Q(\ram[141][7] ), 
	.D(n2845), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][6]  (.Q(\ram[141][6] ), 
	.D(n2844), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[141][5]  (.Q(\ram[141][5] ), 
	.D(n2843), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[141][4]  (.Q(\ram[141][4] ), 
	.D(n2842), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][3]  (.Q(\ram[141][3] ), 
	.D(n2841), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[141][2]  (.Q(\ram[141][2] ), 
	.D(n2840), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][1]  (.Q(\ram[141][1] ), 
	.D(n2839), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][0]  (.Q(\ram[141][0] ), 
	.D(n2838), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[137][15]  (.Q(\ram[137][15] ), 
	.D(n2789), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][14]  (.Q(\ram[137][14] ), 
	.D(n2788), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][13]  (.Q(\ram[137][13] ), 
	.D(n2787), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[137][12]  (.Q(\ram[137][12] ), 
	.D(n2786), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][11]  (.Q(\ram[137][11] ), 
	.D(n2785), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[137][10]  (.Q(\ram[137][10] ), 
	.D(n2784), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[137][9]  (.Q(\ram[137][9] ), 
	.D(n2783), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][8]  (.Q(\ram[137][8] ), 
	.D(n2782), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[137][7]  (.Q(\ram[137][7] ), 
	.D(n2781), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][6]  (.Q(\ram[137][6] ), 
	.D(n2780), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[137][5]  (.Q(\ram[137][5] ), 
	.D(n2779), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][4]  (.Q(\ram[137][4] ), 
	.D(n2778), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][3]  (.Q(\ram[137][3] ), 
	.D(n2777), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][2]  (.Q(\ram[137][2] ), 
	.D(n2776), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[137][1]  (.Q(\ram[137][1] ), 
	.D(n2775), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][0]  (.Q(\ram[137][0] ), 
	.D(n2774), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[133][15]  (.Q(\ram[133][15] ), 
	.D(n2725), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][14]  (.Q(\ram[133][14] ), 
	.D(n2724), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][13]  (.Q(\ram[133][13] ), 
	.D(n2723), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][12]  (.Q(\ram[133][12] ), 
	.D(n2722), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][11]  (.Q(\ram[133][11] ), 
	.D(n2721), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[133][10]  (.Q(\ram[133][10] ), 
	.D(n2720), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[133][9]  (.Q(\ram[133][9] ), 
	.D(n2719), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[133][8]  (.Q(\ram[133][8] ), 
	.D(n2718), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[133][7]  (.Q(\ram[133][7] ), 
	.D(n2717), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][6]  (.Q(\ram[133][6] ), 
	.D(n2716), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][5]  (.Q(\ram[133][5] ), 
	.D(n2715), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][4]  (.Q(\ram[133][4] ), 
	.D(n2714), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[133][3]  (.Q(\ram[133][3] ), 
	.D(n2713), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][2]  (.Q(\ram[133][2] ), 
	.D(n2712), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[133][1]  (.Q(\ram[133][1] ), 
	.D(n2711), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][0]  (.Q(\ram[133][0] ), 
	.D(n2710), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[129][15]  (.Q(\ram[129][15] ), 
	.D(n2661), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][14]  (.Q(\ram[129][14] ), 
	.D(n2660), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][13]  (.Q(\ram[129][13] ), 
	.D(n2659), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][12]  (.Q(\ram[129][12] ), 
	.D(n2658), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[129][11]  (.Q(\ram[129][11] ), 
	.D(n2657), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[129][10]  (.Q(\ram[129][10] ), 
	.D(n2656), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[129][9]  (.Q(\ram[129][9] ), 
	.D(n2655), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][8]  (.Q(\ram[129][8] ), 
	.D(n2654), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[129][7]  (.Q(\ram[129][7] ), 
	.D(n2653), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[129][6]  (.Q(\ram[129][6] ), 
	.D(n2652), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[129][5]  (.Q(\ram[129][5] ), 
	.D(n2651), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[129][4]  (.Q(\ram[129][4] ), 
	.D(n2650), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[129][3]  (.Q(\ram[129][3] ), 
	.D(n2649), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[129][2]  (.Q(\ram[129][2] ), 
	.D(n2648), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[129][1]  (.Q(\ram[129][1] ), 
	.D(n2647), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[129][0]  (.Q(\ram[129][0] ), 
	.D(n2646), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[125][15]  (.Q(\ram[125][15] ), 
	.D(n2597), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][14]  (.Q(\ram[125][14] ), 
	.D(n2596), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][13]  (.Q(\ram[125][13] ), 
	.D(n2595), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][12]  (.Q(\ram[125][12] ), 
	.D(n2594), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[125][11]  (.Q(\ram[125][11] ), 
	.D(n2593), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[125][10]  (.Q(\ram[125][10] ), 
	.D(n2592), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][9]  (.Q(\ram[125][9] ), 
	.D(n2591), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][8]  (.Q(\ram[125][8] ), 
	.D(n2590), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[125][7]  (.Q(\ram[125][7] ), 
	.D(n2589), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][6]  (.Q(\ram[125][6] ), 
	.D(n2588), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][5]  (.Q(\ram[125][5] ), 
	.D(n2587), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][4]  (.Q(\ram[125][4] ), 
	.D(n2586), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][3]  (.Q(\ram[125][3] ), 
	.D(n2585), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[125][2]  (.Q(\ram[125][2] ), 
	.D(n2584), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][1]  (.Q(\ram[125][1] ), 
	.D(n2583), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[125][0]  (.Q(\ram[125][0] ), 
	.D(n2582), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[121][15]  (.Q(\ram[121][15] ), 
	.D(n2533), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][14]  (.Q(\ram[121][14] ), 
	.D(n2532), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][13]  (.Q(\ram[121][13] ), 
	.D(n2531), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[121][12]  (.Q(\ram[121][12] ), 
	.D(n2530), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][11]  (.Q(\ram[121][11] ), 
	.D(n2529), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][10]  (.Q(\ram[121][10] ), 
	.D(n2528), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][9]  (.Q(\ram[121][9] ), 
	.D(n2527), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][8]  (.Q(\ram[121][8] ), 
	.D(n2526), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][7]  (.Q(\ram[121][7] ), 
	.D(n2525), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][6]  (.Q(\ram[121][6] ), 
	.D(n2524), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[121][5]  (.Q(\ram[121][5] ), 
	.D(n2523), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[121][4]  (.Q(\ram[121][4] ), 
	.D(n2522), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[121][3]  (.Q(\ram[121][3] ), 
	.D(n2521), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[121][2]  (.Q(\ram[121][2] ), 
	.D(n2520), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[121][1]  (.Q(\ram[121][1] ), 
	.D(n2519), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[121][0]  (.Q(\ram[121][0] ), 
	.D(n2518), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[117][15]  (.Q(\ram[117][15] ), 
	.D(n2469), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[117][14]  (.Q(\ram[117][14] ), 
	.D(n2468), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][13]  (.Q(\ram[117][13] ), 
	.D(n2467), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[117][12]  (.Q(\ram[117][12] ), 
	.D(n2466), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[117][11]  (.Q(\ram[117][11] ), 
	.D(n2465), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][10]  (.Q(\ram[117][10] ), 
	.D(n2464), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][9]  (.Q(\ram[117][9] ), 
	.D(n2463), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][8]  (.Q(\ram[117][8] ), 
	.D(n2462), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][7]  (.Q(\ram[117][7] ), 
	.D(n2461), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][6]  (.Q(\ram[117][6] ), 
	.D(n2460), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[117][5]  (.Q(\ram[117][5] ), 
	.D(n2459), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[117][4]  (.Q(\ram[117][4] ), 
	.D(n2458), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[117][3]  (.Q(\ram[117][3] ), 
	.D(n2457), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[117][2]  (.Q(\ram[117][2] ), 
	.D(n2456), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][1]  (.Q(\ram[117][1] ), 
	.D(n2455), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[117][0]  (.Q(\ram[117][0] ), 
	.D(n2454), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[113][15]  (.Q(\ram[113][15] ), 
	.D(n2405), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[113][14]  (.Q(\ram[113][14] ), 
	.D(n2404), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[113][13]  (.Q(\ram[113][13] ), 
	.D(n2403), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][12]  (.Q(\ram[113][12] ), 
	.D(n2402), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[113][11]  (.Q(\ram[113][11] ), 
	.D(n2401), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][10]  (.Q(\ram[113][10] ), 
	.D(n2400), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][9]  (.Q(\ram[113][9] ), 
	.D(n2399), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][8]  (.Q(\ram[113][8] ), 
	.D(n2398), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][7]  (.Q(\ram[113][7] ), 
	.D(n2397), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][6]  (.Q(\ram[113][6] ), 
	.D(n2396), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][5]  (.Q(\ram[113][5] ), 
	.D(n2395), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[113][4]  (.Q(\ram[113][4] ), 
	.D(n2394), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][3]  (.Q(\ram[113][3] ), 
	.D(n2393), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][2]  (.Q(\ram[113][2] ), 
	.D(n2392), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][1]  (.Q(\ram[113][1] ), 
	.D(n2391), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][0]  (.Q(\ram[113][0] ), 
	.D(n2390), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[109][15]  (.Q(\ram[109][15] ), 
	.D(n2341), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][14]  (.Q(\ram[109][14] ), 
	.D(n2340), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[109][13]  (.Q(\ram[109][13] ), 
	.D(n2339), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[109][12]  (.Q(\ram[109][12] ), 
	.D(n2338), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[109][11]  (.Q(\ram[109][11] ), 
	.D(n2337), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[109][10]  (.Q(\ram[109][10] ), 
	.D(n2336), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][9]  (.Q(\ram[109][9] ), 
	.D(n2335), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[109][8]  (.Q(\ram[109][8] ), 
	.D(n2334), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][7]  (.Q(\ram[109][7] ), 
	.D(n2333), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[109][6]  (.Q(\ram[109][6] ), 
	.D(n2332), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][5]  (.Q(\ram[109][5] ), 
	.D(n2331), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[109][4]  (.Q(\ram[109][4] ), 
	.D(n2330), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[109][3]  (.Q(\ram[109][3] ), 
	.D(n2329), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][2]  (.Q(\ram[109][2] ), 
	.D(n2328), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][1]  (.Q(\ram[109][1] ), 
	.D(n2327), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][0]  (.Q(\ram[109][0] ), 
	.D(n2326), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[105][15]  (.Q(\ram[105][15] ), 
	.D(n2277), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][14]  (.Q(\ram[105][14] ), 
	.D(n2276), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][13]  (.Q(\ram[105][13] ), 
	.D(n2275), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[105][12]  (.Q(\ram[105][12] ), 
	.D(n2274), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][11]  (.Q(\ram[105][11] ), 
	.D(n2273), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][10]  (.Q(\ram[105][10] ), 
	.D(n2272), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[105][9]  (.Q(\ram[105][9] ), 
	.D(n2271), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][8]  (.Q(\ram[105][8] ), 
	.D(n2270), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[105][7]  (.Q(\ram[105][7] ), 
	.D(n2269), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[105][6]  (.Q(\ram[105][6] ), 
	.D(n2268), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][5]  (.Q(\ram[105][5] ), 
	.D(n2267), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][4]  (.Q(\ram[105][4] ), 
	.D(n2266), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[105][3]  (.Q(\ram[105][3] ), 
	.D(n2265), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][2]  (.Q(\ram[105][2] ), 
	.D(n2264), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][1]  (.Q(\ram[105][1] ), 
	.D(n2263), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[105][0]  (.Q(\ram[105][0] ), 
	.D(n2262), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[101][15]  (.Q(\ram[101][15] ), 
	.D(n2213), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[101][14]  (.Q(\ram[101][14] ), 
	.D(n2212), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][13]  (.Q(\ram[101][13] ), 
	.D(n2211), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[101][12]  (.Q(\ram[101][12] ), 
	.D(n2210), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[101][11]  (.Q(\ram[101][11] ), 
	.D(n2209), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[101][10]  (.Q(\ram[101][10] ), 
	.D(n2208), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][9]  (.Q(\ram[101][9] ), 
	.D(n2207), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][8]  (.Q(\ram[101][8] ), 
	.D(n2206), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][7]  (.Q(\ram[101][7] ), 
	.D(n2205), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[101][6]  (.Q(\ram[101][6] ), 
	.D(n2204), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][5]  (.Q(\ram[101][5] ), 
	.D(n2203), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][4]  (.Q(\ram[101][4] ), 
	.D(n2202), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[101][3]  (.Q(\ram[101][3] ), 
	.D(n2201), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[101][2]  (.Q(\ram[101][2] ), 
	.D(n2200), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][1]  (.Q(\ram[101][1] ), 
	.D(n2199), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[101][0]  (.Q(\ram[101][0] ), 
	.D(n2198), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[97][15]  (.Q(\ram[97][15] ), 
	.D(n2149), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][14]  (.Q(\ram[97][14] ), 
	.D(n2148), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][13]  (.Q(\ram[97][13] ), 
	.D(n2147), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[97][12]  (.Q(\ram[97][12] ), 
	.D(n2146), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[97][11]  (.Q(\ram[97][11] ), 
	.D(n2145), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[97][10]  (.Q(\ram[97][10] ), 
	.D(n2144), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[97][9]  (.Q(\ram[97][9] ), 
	.D(n2143), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[97][8]  (.Q(\ram[97][8] ), 
	.D(n2142), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][7]  (.Q(\ram[97][7] ), 
	.D(n2141), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[97][6]  (.Q(\ram[97][6] ), 
	.D(n2140), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][5]  (.Q(\ram[97][5] ), 
	.D(n2139), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[97][4]  (.Q(\ram[97][4] ), 
	.D(n2138), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[97][3]  (.Q(\ram[97][3] ), 
	.D(n2137), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[97][2]  (.Q(\ram[97][2] ), 
	.D(n2136), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[97][1]  (.Q(\ram[97][1] ), 
	.D(n2135), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[97][0]  (.Q(\ram[97][0] ), 
	.D(n2134), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[93][15]  (.Q(\ram[93][15] ), 
	.D(n2085), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][14]  (.Q(\ram[93][14] ), 
	.D(n2084), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][13]  (.Q(\ram[93][13] ), 
	.D(n2083), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[93][12]  (.Q(\ram[93][12] ), 
	.D(n2082), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][11]  (.Q(\ram[93][11] ), 
	.D(n2081), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][10]  (.Q(\ram[93][10] ), 
	.D(n2080), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[93][9]  (.Q(\ram[93][9] ), 
	.D(n2079), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][8]  (.Q(\ram[93][8] ), 
	.D(n2078), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[93][7]  (.Q(\ram[93][7] ), 
	.D(n2077), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][6]  (.Q(\ram[93][6] ), 
	.D(n2076), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][5]  (.Q(\ram[93][5] ), 
	.D(n2075), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][4]  (.Q(\ram[93][4] ), 
	.D(n2074), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][3]  (.Q(\ram[93][3] ), 
	.D(n2073), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][2]  (.Q(\ram[93][2] ), 
	.D(n2072), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][1]  (.Q(\ram[93][1] ), 
	.D(n2071), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[93][0]  (.Q(\ram[93][0] ), 
	.D(n2070), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[89][15]  (.Q(\ram[89][15] ), 
	.D(n2021), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][14]  (.Q(\ram[89][14] ), 
	.D(n2020), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[89][13]  (.Q(\ram[89][13] ), 
	.D(n2019), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][12]  (.Q(\ram[89][12] ), 
	.D(n2018), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[89][11]  (.Q(\ram[89][11] ), 
	.D(n2017), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[89][10]  (.Q(\ram[89][10] ), 
	.D(n2016), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][9]  (.Q(\ram[89][9] ), 
	.D(n2015), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][8]  (.Q(\ram[89][8] ), 
	.D(n2014), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][7]  (.Q(\ram[89][7] ), 
	.D(n2013), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][6]  (.Q(\ram[89][6] ), 
	.D(n2012), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][5]  (.Q(\ram[89][5] ), 
	.D(n2011), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[89][4]  (.Q(\ram[89][4] ), 
	.D(n2010), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][3]  (.Q(\ram[89][3] ), 
	.D(n2009), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][2]  (.Q(\ram[89][2] ), 
	.D(n2008), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][1]  (.Q(\ram[89][1] ), 
	.D(n2007), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[89][0]  (.Q(\ram[89][0] ), 
	.D(n2006), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[85][15]  (.Q(\ram[85][15] ), 
	.D(n1957), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][14]  (.Q(\ram[85][14] ), 
	.D(n1956), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][13]  (.Q(\ram[85][13] ), 
	.D(n1955), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][12]  (.Q(\ram[85][12] ), 
	.D(n1954), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][11]  (.Q(\ram[85][11] ), 
	.D(n1953), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][10]  (.Q(\ram[85][10] ), 
	.D(n1952), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[85][9]  (.Q(\ram[85][9] ), 
	.D(n1951), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][8]  (.Q(\ram[85][8] ), 
	.D(n1950), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][7]  (.Q(\ram[85][7] ), 
	.D(n1949), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[85][6]  (.Q(\ram[85][6] ), 
	.D(n1948), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][5]  (.Q(\ram[85][5] ), 
	.D(n1947), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][4]  (.Q(\ram[85][4] ), 
	.D(n1946), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][3]  (.Q(\ram[85][3] ), 
	.D(n1945), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][2]  (.Q(\ram[85][2] ), 
	.D(n1944), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][1]  (.Q(\ram[85][1] ), 
	.D(n1943), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[85][0]  (.Q(\ram[85][0] ), 
	.D(n1942), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[81][15]  (.Q(\ram[81][15] ), 
	.D(n1893), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][14]  (.Q(\ram[81][14] ), 
	.D(n1892), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][13]  (.Q(\ram[81][13] ), 
	.D(n1891), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][12]  (.Q(\ram[81][12] ), 
	.D(n1890), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][11]  (.Q(\ram[81][11] ), 
	.D(n1889), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][10]  (.Q(\ram[81][10] ), 
	.D(n1888), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[81][9]  (.Q(\ram[81][9] ), 
	.D(n1887), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[81][8]  (.Q(\ram[81][8] ), 
	.D(n1886), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[81][7]  (.Q(\ram[81][7] ), 
	.D(n1885), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[81][6]  (.Q(\ram[81][6] ), 
	.D(n1884), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][5]  (.Q(\ram[81][5] ), 
	.D(n1883), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][4]  (.Q(\ram[81][4] ), 
	.D(n1882), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][3]  (.Q(\ram[81][3] ), 
	.D(n1881), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][2]  (.Q(\ram[81][2] ), 
	.D(n1880), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][1]  (.Q(\ram[81][1] ), 
	.D(n1879), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[81][0]  (.Q(\ram[81][0] ), 
	.D(n1878), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[77][15]  (.Q(\ram[77][15] ), 
	.D(n1829), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][14]  (.Q(\ram[77][14] ), 
	.D(n1828), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][13]  (.Q(\ram[77][13] ), 
	.D(n1827), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][12]  (.Q(\ram[77][12] ), 
	.D(n1826), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][11]  (.Q(\ram[77][11] ), 
	.D(n1825), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][10]  (.Q(\ram[77][10] ), 
	.D(n1824), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][9]  (.Q(\ram[77][9] ), 
	.D(n1823), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][8]  (.Q(\ram[77][8] ), 
	.D(n1822), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][7]  (.Q(\ram[77][7] ), 
	.D(n1821), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][6]  (.Q(\ram[77][6] ), 
	.D(n1820), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[77][5]  (.Q(\ram[77][5] ), 
	.D(n1819), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][4]  (.Q(\ram[77][4] ), 
	.D(n1818), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][3]  (.Q(\ram[77][3] ), 
	.D(n1817), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[77][2]  (.Q(\ram[77][2] ), 
	.D(n1816), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][1]  (.Q(\ram[77][1] ), 
	.D(n1815), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][0]  (.Q(\ram[77][0] ), 
	.D(n1814), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[73][15]  (.Q(\ram[73][15] ), 
	.D(n1765), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][14]  (.Q(\ram[73][14] ), 
	.D(n1764), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][13]  (.Q(\ram[73][13] ), 
	.D(n1763), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[73][12]  (.Q(\ram[73][12] ), 
	.D(n1762), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][11]  (.Q(\ram[73][11] ), 
	.D(n1761), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][10]  (.Q(\ram[73][10] ), 
	.D(n1760), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][9]  (.Q(\ram[73][9] ), 
	.D(n1759), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][8]  (.Q(\ram[73][8] ), 
	.D(n1758), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[73][7]  (.Q(\ram[73][7] ), 
	.D(n1757), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][6]  (.Q(\ram[73][6] ), 
	.D(n1756), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][5]  (.Q(\ram[73][5] ), 
	.D(n1755), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][4]  (.Q(\ram[73][4] ), 
	.D(n1754), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][3]  (.Q(\ram[73][3] ), 
	.D(n1753), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[73][2]  (.Q(\ram[73][2] ), 
	.D(n1752), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][1]  (.Q(\ram[73][1] ), 
	.D(n1751), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[73][0]  (.Q(\ram[73][0] ), 
	.D(n1750), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[69][15]  (.Q(\ram[69][15] ), 
	.D(n1701), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[69][14]  (.Q(\ram[69][14] ), 
	.D(n1700), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][13]  (.Q(\ram[69][13] ), 
	.D(n1699), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[69][12]  (.Q(\ram[69][12] ), 
	.D(n1698), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][11]  (.Q(\ram[69][11] ), 
	.D(n1697), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][10]  (.Q(\ram[69][10] ), 
	.D(n1696), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][9]  (.Q(\ram[69][9] ), 
	.D(n1695), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][8]  (.Q(\ram[69][8] ), 
	.D(n1694), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][7]  (.Q(\ram[69][7] ), 
	.D(n1693), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[69][6]  (.Q(\ram[69][6] ), 
	.D(n1692), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[69][5]  (.Q(\ram[69][5] ), 
	.D(n1691), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][4]  (.Q(\ram[69][4] ), 
	.D(n1690), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][3]  (.Q(\ram[69][3] ), 
	.D(n1689), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][2]  (.Q(\ram[69][2] ), 
	.D(n1688), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][1]  (.Q(\ram[69][1] ), 
	.D(n1687), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[69][0]  (.Q(\ram[69][0] ), 
	.D(n1686), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[65][15]  (.Q(\ram[65][15] ), 
	.D(n1637), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[65][14]  (.Q(\ram[65][14] ), 
	.D(n1636), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][13]  (.Q(\ram[65][13] ), 
	.D(n1635), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][12]  (.Q(\ram[65][12] ), 
	.D(n1634), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[65][11]  (.Q(\ram[65][11] ), 
	.D(n1633), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][10]  (.Q(\ram[65][10] ), 
	.D(n1632), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][9]  (.Q(\ram[65][9] ), 
	.D(n1631), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][8]  (.Q(\ram[65][8] ), 
	.D(n1630), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][7]  (.Q(\ram[65][7] ), 
	.D(n1629), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[65][6]  (.Q(\ram[65][6] ), 
	.D(n1628), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[65][5]  (.Q(\ram[65][5] ), 
	.D(n1627), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[65][4]  (.Q(\ram[65][4] ), 
	.D(n1626), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][3]  (.Q(\ram[65][3] ), 
	.D(n1625), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][2]  (.Q(\ram[65][2] ), 
	.D(n1624), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[65][1]  (.Q(\ram[65][1] ), 
	.D(n1623), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][0]  (.Q(\ram[65][0] ), 
	.D(n1622), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[61][15]  (.Q(\ram[61][15] ), 
	.D(n1573), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][14]  (.Q(\ram[61][14] ), 
	.D(n1572), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[61][13]  (.Q(\ram[61][13] ), 
	.D(n1571), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[61][12]  (.Q(\ram[61][12] ), 
	.D(n1570), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][11]  (.Q(\ram[61][11] ), 
	.D(n1569), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][10]  (.Q(\ram[61][10] ), 
	.D(n1568), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][9]  (.Q(\ram[61][9] ), 
	.D(n1567), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[61][8]  (.Q(\ram[61][8] ), 
	.D(n1566), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][7]  (.Q(\ram[61][7] ), 
	.D(n1565), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][6]  (.Q(\ram[61][6] ), 
	.D(n1564), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][5]  (.Q(\ram[61][5] ), 
	.D(n1563), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][4]  (.Q(\ram[61][4] ), 
	.D(n1562), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][3]  (.Q(\ram[61][3] ), 
	.D(n1561), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][2]  (.Q(\ram[61][2] ), 
	.D(n1560), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][1]  (.Q(\ram[61][1] ), 
	.D(n1559), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[61][0]  (.Q(\ram[61][0] ), 
	.D(n1558), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[57][15]  (.Q(\ram[57][15] ), 
	.D(n1509), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[57][14]  (.Q(\ram[57][14] ), 
	.D(n1508), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[57][13]  (.Q(\ram[57][13] ), 
	.D(n1507), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[57][12]  (.Q(\ram[57][12] ), 
	.D(n1506), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[57][11]  (.Q(\ram[57][11] ), 
	.D(n1505), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][10]  (.Q(\ram[57][10] ), 
	.D(n1504), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][9]  (.Q(\ram[57][9] ), 
	.D(n1503), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[57][8]  (.Q(\ram[57][8] ), 
	.D(n1502), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[57][7]  (.Q(\ram[57][7] ), 
	.D(n1501), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[57][6]  (.Q(\ram[57][6] ), 
	.D(n1500), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][5]  (.Q(\ram[57][5] ), 
	.D(n1499), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][4]  (.Q(\ram[57][4] ), 
	.D(n1498), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[57][3]  (.Q(\ram[57][3] ), 
	.D(n1497), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[57][2]  (.Q(\ram[57][2] ), 
	.D(n1496), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[57][1]  (.Q(\ram[57][1] ), 
	.D(n1495), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[57][0]  (.Q(\ram[57][0] ), 
	.D(n1494), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[53][15]  (.Q(\ram[53][15] ), 
	.D(n1445), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][14]  (.Q(\ram[53][14] ), 
	.D(n1444), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][13]  (.Q(\ram[53][13] ), 
	.D(n1443), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][12]  (.Q(\ram[53][12] ), 
	.D(n1442), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][11]  (.Q(\ram[53][11] ), 
	.D(n1441), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][10]  (.Q(\ram[53][10] ), 
	.D(n1440), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[53][9]  (.Q(\ram[53][9] ), 
	.D(n1439), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][8]  (.Q(\ram[53][8] ), 
	.D(n1438), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][7]  (.Q(\ram[53][7] ), 
	.D(n1437), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[53][6]  (.Q(\ram[53][6] ), 
	.D(n1436), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[53][5]  (.Q(\ram[53][5] ), 
	.D(n1435), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[53][4]  (.Q(\ram[53][4] ), 
	.D(n1434), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][3]  (.Q(\ram[53][3] ), 
	.D(n1433), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][2]  (.Q(\ram[53][2] ), 
	.D(n1432), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][1]  (.Q(\ram[53][1] ), 
	.D(n1431), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][0]  (.Q(\ram[53][0] ), 
	.D(n1430), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[49][15]  (.Q(\ram[49][15] ), 
	.D(n1381), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[49][14]  (.Q(\ram[49][14] ), 
	.D(n1380), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[49][13]  (.Q(\ram[49][13] ), 
	.D(n1379), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[49][12]  (.Q(\ram[49][12] ), 
	.D(n1378), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][11]  (.Q(\ram[49][11] ), 
	.D(n1377), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][10]  (.Q(\ram[49][10] ), 
	.D(n1376), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][9]  (.Q(\ram[49][9] ), 
	.D(n1375), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[49][8]  (.Q(\ram[49][8] ), 
	.D(n1374), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[49][7]  (.Q(\ram[49][7] ), 
	.D(n1373), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[49][6]  (.Q(\ram[49][6] ), 
	.D(n1372), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[49][5]  (.Q(\ram[49][5] ), 
	.D(n1371), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][4]  (.Q(\ram[49][4] ), 
	.D(n1370), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][3]  (.Q(\ram[49][3] ), 
	.D(n1369), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[49][2]  (.Q(\ram[49][2] ), 
	.D(n1368), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[49][1]  (.Q(\ram[49][1] ), 
	.D(n1367), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[49][0]  (.Q(\ram[49][0] ), 
	.D(n1366), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[45][15]  (.Q(\ram[45][15] ), 
	.D(n1317), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][14]  (.Q(\ram[45][14] ), 
	.D(n1316), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][13]  (.Q(\ram[45][13] ), 
	.D(n1315), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][12]  (.Q(\ram[45][12] ), 
	.D(n1314), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][11]  (.Q(\ram[45][11] ), 
	.D(n1313), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][10]  (.Q(\ram[45][10] ), 
	.D(n1312), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[45][9]  (.Q(\ram[45][9] ), 
	.D(n1311), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][8]  (.Q(\ram[45][8] ), 
	.D(n1310), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[45][7]  (.Q(\ram[45][7] ), 
	.D(n1309), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][6]  (.Q(\ram[45][6] ), 
	.D(n1308), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][5]  (.Q(\ram[45][5] ), 
	.D(n1307), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][4]  (.Q(\ram[45][4] ), 
	.D(n1306), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][3]  (.Q(\ram[45][3] ), 
	.D(n1305), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][2]  (.Q(\ram[45][2] ), 
	.D(n1304), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[45][1]  (.Q(\ram[45][1] ), 
	.D(n1303), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][0]  (.Q(\ram[45][0] ), 
	.D(n1302), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[41][15]  (.Q(\ram[41][15] ), 
	.D(n1253), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][14]  (.Q(\ram[41][14] ), 
	.D(n1252), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][13]  (.Q(\ram[41][13] ), 
	.D(n1251), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[41][12]  (.Q(\ram[41][12] ), 
	.D(n1250), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[41][11]  (.Q(\ram[41][11] ), 
	.D(n1249), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[41][10]  (.Q(\ram[41][10] ), 
	.D(n1248), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][9]  (.Q(\ram[41][9] ), 
	.D(n1247), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][8]  (.Q(\ram[41][8] ), 
	.D(n1246), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][7]  (.Q(\ram[41][7] ), 
	.D(n1245), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][6]  (.Q(\ram[41][6] ), 
	.D(n1244), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[41][5]  (.Q(\ram[41][5] ), 
	.D(n1243), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[41][4]  (.Q(\ram[41][4] ), 
	.D(n1242), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][3]  (.Q(\ram[41][3] ), 
	.D(n1241), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[41][2]  (.Q(\ram[41][2] ), 
	.D(n1240), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][1]  (.Q(\ram[41][1] ), 
	.D(n1239), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[41][0]  (.Q(\ram[41][0] ), 
	.D(n1238), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[37][15]  (.Q(\ram[37][15] ), 
	.D(n1189), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][14]  (.Q(\ram[37][14] ), 
	.D(n1188), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][13]  (.Q(\ram[37][13] ), 
	.D(n1187), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][12]  (.Q(\ram[37][12] ), 
	.D(n1186), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[37][11]  (.Q(\ram[37][11] ), 
	.D(n1185), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[37][10]  (.Q(\ram[37][10] ), 
	.D(n1184), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[37][9]  (.Q(\ram[37][9] ), 
	.D(n1183), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[37][8]  (.Q(\ram[37][8] ), 
	.D(n1182), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][7]  (.Q(\ram[37][7] ), 
	.D(n1181), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[37][6]  (.Q(\ram[37][6] ), 
	.D(n1180), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[37][5]  (.Q(\ram[37][5] ), 
	.D(n1179), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[37][4]  (.Q(\ram[37][4] ), 
	.D(n1178), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[37][3]  (.Q(\ram[37][3] ), 
	.D(n1177), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[37][2]  (.Q(\ram[37][2] ), 
	.D(n1176), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][1]  (.Q(\ram[37][1] ), 
	.D(n1175), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[37][0]  (.Q(\ram[37][0] ), 
	.D(n1174), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[33][15]  (.Q(\ram[33][15] ), 
	.D(n1125), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[33][14]  (.Q(\ram[33][14] ), 
	.D(n1124), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][13]  (.Q(\ram[33][13] ), 
	.D(n1123), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[33][12]  (.Q(\ram[33][12] ), 
	.D(n1122), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][11]  (.Q(\ram[33][11] ), 
	.D(n1121), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][10]  (.Q(\ram[33][10] ), 
	.D(n1120), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[33][9]  (.Q(\ram[33][9] ), 
	.D(n1119), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[33][8]  (.Q(\ram[33][8] ), 
	.D(n1118), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][7]  (.Q(\ram[33][7] ), 
	.D(n1117), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[33][6]  (.Q(\ram[33][6] ), 
	.D(n1116), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][5]  (.Q(\ram[33][5] ), 
	.D(n1115), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][4]  (.Q(\ram[33][4] ), 
	.D(n1114), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][3]  (.Q(\ram[33][3] ), 
	.D(n1113), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][2]  (.Q(\ram[33][2] ), 
	.D(n1112), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][1]  (.Q(\ram[33][1] ), 
	.D(n1111), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[33][0]  (.Q(\ram[33][0] ), 
	.D(n1110), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[29][15]  (.Q(\ram[29][15] ), 
	.D(n1061), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[29][14]  (.Q(\ram[29][14] ), 
	.D(n1060), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][13]  (.Q(\ram[29][13] ), 
	.D(n1059), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[29][12]  (.Q(\ram[29][12] ), 
	.D(n1058), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[29][11]  (.Q(\ram[29][11] ), 
	.D(n1057), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][10]  (.Q(\ram[29][10] ), 
	.D(n1056), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[29][9]  (.Q(\ram[29][9] ), 
	.D(n1055), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][8]  (.Q(\ram[29][8] ), 
	.D(n1054), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][7]  (.Q(\ram[29][7] ), 
	.D(n1053), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][6]  (.Q(\ram[29][6] ), 
	.D(n1052), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][5]  (.Q(\ram[29][5] ), 
	.D(n1051), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][4]  (.Q(\ram[29][4] ), 
	.D(n1050), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[29][3]  (.Q(\ram[29][3] ), 
	.D(n1049), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][2]  (.Q(\ram[29][2] ), 
	.D(n1048), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[29][1]  (.Q(\ram[29][1] ), 
	.D(n1047), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][0]  (.Q(\ram[29][0] ), 
	.D(n1046), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][15]  (.Q(\ram[25][15] ), 
	.D(n997), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[25][14]  (.Q(\ram[25][14] ), 
	.D(n996), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][13]  (.Q(\ram[25][13] ), 
	.D(n995), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[25][12]  (.Q(\ram[25][12] ), 
	.D(n994), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][11]  (.Q(\ram[25][11] ), 
	.D(n993), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[25][10]  (.Q(\ram[25][10] ), 
	.D(n992), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][9]  (.Q(\ram[25][9] ), 
	.D(n991), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[25][8]  (.Q(\ram[25][8] ), 
	.D(n990), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[25][7]  (.Q(\ram[25][7] ), 
	.D(n989), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][6]  (.Q(\ram[25][6] ), 
	.D(n988), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[25][5]  (.Q(\ram[25][5] ), 
	.D(n987), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[25][4]  (.Q(\ram[25][4] ), 
	.D(n986), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][3]  (.Q(\ram[25][3] ), 
	.D(n985), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[25][2]  (.Q(\ram[25][2] ), 
	.D(n984), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][1]  (.Q(\ram[25][1] ), 
	.D(n983), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][0]  (.Q(\ram[25][0] ), 
	.D(n982), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[21][15]  (.Q(\ram[21][15] ), 
	.D(n933), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[21][14]  (.Q(\ram[21][14] ), 
	.D(n932), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][13]  (.Q(\ram[21][13] ), 
	.D(n931), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[21][12]  (.Q(\ram[21][12] ), 
	.D(n930), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[21][11]  (.Q(\ram[21][11] ), 
	.D(n929), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][10]  (.Q(\ram[21][10] ), 
	.D(n928), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[21][9]  (.Q(\ram[21][9] ), 
	.D(n927), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][8]  (.Q(\ram[21][8] ), 
	.D(n926), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[21][7]  (.Q(\ram[21][7] ), 
	.D(n925), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][6]  (.Q(\ram[21][6] ), 
	.D(n924), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[21][5]  (.Q(\ram[21][5] ), 
	.D(n923), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[21][4]  (.Q(\ram[21][4] ), 
	.D(n922), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[21][3]  (.Q(\ram[21][3] ), 
	.D(n921), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][2]  (.Q(\ram[21][2] ), 
	.D(n920), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[21][1]  (.Q(\ram[21][1] ), 
	.D(n919), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[21][0]  (.Q(\ram[21][0] ), 
	.D(n918), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[17][15]  (.Q(\ram[17][15] ), 
	.D(n869), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[17][14]  (.Q(\ram[17][14] ), 
	.D(n868), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][13]  (.Q(\ram[17][13] ), 
	.D(n867), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][12]  (.Q(\ram[17][12] ), 
	.D(n866), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][11]  (.Q(\ram[17][11] ), 
	.D(n865), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][10]  (.Q(\ram[17][10] ), 
	.D(n864), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[17][9]  (.Q(\ram[17][9] ), 
	.D(n863), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][8]  (.Q(\ram[17][8] ), 
	.D(n862), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[17][7]  (.Q(\ram[17][7] ), 
	.D(n861), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][6]  (.Q(\ram[17][6] ), 
	.D(n860), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[17][5]  (.Q(\ram[17][5] ), 
	.D(n859), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[17][4]  (.Q(\ram[17][4] ), 
	.D(n858), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[17][3]  (.Q(\ram[17][3] ), 
	.D(n857), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][2]  (.Q(\ram[17][2] ), 
	.D(n856), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[17][1]  (.Q(\ram[17][1] ), 
	.D(n855), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][0]  (.Q(\ram[17][0] ), 
	.D(n854), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[13][15]  (.Q(\ram[13][15] ), 
	.D(n805), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[13][14]  (.Q(\ram[13][14] ), 
	.D(n804), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[13][13]  (.Q(\ram[13][13] ), 
	.D(n803), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][12]  (.Q(\ram[13][12] ), 
	.D(n802), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[13][11]  (.Q(\ram[13][11] ), 
	.D(n801), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][10]  (.Q(\ram[13][10] ), 
	.D(n800), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[13][9]  (.Q(\ram[13][9] ), 
	.D(n799), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[13][8]  (.Q(\ram[13][8] ), 
	.D(n798), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][7]  (.Q(\ram[13][7] ), 
	.D(n797), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[13][6]  (.Q(\ram[13][6] ), 
	.D(n796), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][5]  (.Q(\ram[13][5] ), 
	.D(n795), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][4]  (.Q(\ram[13][4] ), 
	.D(n794), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][3]  (.Q(\ram[13][3] ), 
	.D(n793), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][2]  (.Q(\ram[13][2] ), 
	.D(n792), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][1]  (.Q(\ram[13][1] ), 
	.D(n791), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[13][0]  (.Q(\ram[13][0] ), 
	.D(n790), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][15]  (.Q(\ram[9][15] ), 
	.D(n741), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][14]  (.Q(\ram[9][14] ), 
	.D(n740), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[9][13]  (.Q(\ram[9][13] ), 
	.D(n739), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[9][12]  (.Q(\ram[9][12] ), 
	.D(n738), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][11]  (.Q(\ram[9][11] ), 
	.D(n737), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][10]  (.Q(\ram[9][10] ), 
	.D(n736), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][9]  (.Q(\ram[9][9] ), 
	.D(n735), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][8]  (.Q(\ram[9][8] ), 
	.D(n734), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][7]  (.Q(\ram[9][7] ), 
	.D(n733), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][6]  (.Q(\ram[9][6] ), 
	.D(n732), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][5]  (.Q(\ram[9][5] ), 
	.D(n731), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][4]  (.Q(\ram[9][4] ), 
	.D(n730), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][3]  (.Q(\ram[9][3] ), 
	.D(n729), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][2]  (.Q(\ram[9][2] ), 
	.D(n728), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[9][1]  (.Q(\ram[9][1] ), 
	.D(n727), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][0]  (.Q(\ram[9][0] ), 
	.D(n726), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[5][15]  (.Q(\ram[5][15] ), 
	.D(n677), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][14]  (.Q(\ram[5][14] ), 
	.D(n676), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][13]  (.Q(\ram[5][13] ), 
	.D(n675), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[5][12]  (.Q(\ram[5][12] ), 
	.D(n674), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[5][11]  (.Q(\ram[5][11] ), 
	.D(n673), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[5][10]  (.Q(\ram[5][10] ), 
	.D(n672), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][9]  (.Q(\ram[5][9] ), 
	.D(n671), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[5][8]  (.Q(\ram[5][8] ), 
	.D(n670), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][7]  (.Q(\ram[5][7] ), 
	.D(n669), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][6]  (.Q(\ram[5][6] ), 
	.D(n668), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][5]  (.Q(\ram[5][5] ), 
	.D(n667), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[5][4]  (.Q(\ram[5][4] ), 
	.D(n666), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][3]  (.Q(\ram[5][3] ), 
	.D(n665), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[5][2]  (.Q(\ram[5][2] ), 
	.D(n664), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[5][1]  (.Q(\ram[5][1] ), 
	.D(n663), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][0]  (.Q(\ram[5][0] ), 
	.D(n662), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[1][15]  (.Q(\ram[1][15] ), 
	.D(n613), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[1][14]  (.Q(\ram[1][14] ), 
	.D(n612), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[1][13]  (.Q(\ram[1][13] ), 
	.D(n611), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[1][12]  (.Q(\ram[1][12] ), 
	.D(n610), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[1][11]  (.Q(\ram[1][11] ), 
	.D(n609), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[1][10]  (.Q(\ram[1][10] ), 
	.D(n608), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[1][9]  (.Q(\ram[1][9] ), 
	.D(n607), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[1][8]  (.Q(\ram[1][8] ), 
	.D(n606), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[1][7]  (.Q(\ram[1][7] ), 
	.D(n605), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[1][6]  (.Q(\ram[1][6] ), 
	.D(n604), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[1][5]  (.Q(\ram[1][5] ), 
	.D(n603), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[1][4]  (.Q(\ram[1][4] ), 
	.D(n602), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[1][3]  (.Q(\ram[1][3] ), 
	.D(n601), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[1][2]  (.Q(\ram[1][2] ), 
	.D(n600), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[1][1]  (.Q(\ram[1][1] ), 
	.D(n599), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[1][0]  (.Q(\ram[1][0] ), 
	.D(n598), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[254][15]  (.Q(\ram[254][15] ), 
	.D(n4661), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[254][14]  (.Q(\ram[254][14] ), 
	.D(n4660), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[254][13]  (.Q(\ram[254][13] ), 
	.D(n4659), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[254][12]  (.Q(\ram[254][12] ), 
	.D(n4658), 
	.CK(clk));
   QDFFEHD \ram_reg[254][11]  (.Q(\ram[254][11] ), 
	.D(n4657), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][10]  (.Q(\ram[254][10] ), 
	.D(n4656), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[254][9]  (.Q(\ram[254][9] ), 
	.D(n4655), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][8]  (.Q(\ram[254][8] ), 
	.D(n4654), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][7]  (.Q(\ram[254][7] ), 
	.D(n4653), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[254][6]  (.Q(\ram[254][6] ), 
	.D(n4652), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][5]  (.Q(\ram[254][5] ), 
	.D(n4651), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[254][4]  (.Q(\ram[254][4] ), 
	.D(n4650), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[254][3]  (.Q(\ram[254][3] ), 
	.D(n4649), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[254][2]  (.Q(\ram[254][2] ), 
	.D(n4648), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[254][1]  (.Q(\ram[254][1] ), 
	.D(n4647), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[254][0]  (.Q(\ram[254][0] ), 
	.D(n4646), 
	.CK(clk));
   QDFFEHD \ram_reg[250][15]  (.Q(\ram[250][15] ), 
	.D(n4597), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][14]  (.Q(\ram[250][14] ), 
	.D(n4596), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][13]  (.Q(\ram[250][13] ), 
	.D(n4595), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[250][12]  (.Q(\ram[250][12] ), 
	.D(n4594), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][11]  (.Q(\ram[250][11] ), 
	.D(n4593), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][10]  (.Q(\ram[250][10] ), 
	.D(n4592), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][9]  (.Q(\ram[250][9] ), 
	.D(n4591), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[250][8]  (.Q(\ram[250][8] ), 
	.D(n4590), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[250][7]  (.Q(\ram[250][7] ), 
	.D(n4589), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][6]  (.Q(\ram[250][6] ), 
	.D(n4588), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[250][5]  (.Q(\ram[250][5] ), 
	.D(n4587), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][4]  (.Q(\ram[250][4] ), 
	.D(n4586), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][3]  (.Q(\ram[250][3] ), 
	.D(n4585), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[250][2]  (.Q(\ram[250][2] ), 
	.D(n4584), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][1]  (.Q(\ram[250][1] ), 
	.D(n4583), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[250][0]  (.Q(\ram[250][0] ), 
	.D(n4582), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[246][15]  (.Q(\ram[246][15] ), 
	.D(n4533), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[246][14]  (.Q(\ram[246][14] ), 
	.D(n4532), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[246][13]  (.Q(\ram[246][13] ), 
	.D(n4531), 
	.CK(clk));
   QDFFEHD \ram_reg[246][12]  (.Q(\ram[246][12] ), 
	.D(n4530), 
	.CK(clk));
   QDFFEHD \ram_reg[246][11]  (.Q(\ram[246][11] ), 
	.D(n4529), 
	.CK(clk));
   QDFFEHD \ram_reg[246][10]  (.Q(\ram[246][10] ), 
	.D(n4528), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][9]  (.Q(\ram[246][9] ), 
	.D(n4527), 
	.CK(clk));
   QDFFEHD \ram_reg[246][8]  (.Q(\ram[246][8] ), 
	.D(n4526), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][7]  (.Q(\ram[246][7] ), 
	.D(n4525), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[246][6]  (.Q(\ram[246][6] ), 
	.D(n4524), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[246][5]  (.Q(\ram[246][5] ), 
	.D(n4523), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][4]  (.Q(\ram[246][4] ), 
	.D(n4522), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[246][3]  (.Q(\ram[246][3] ), 
	.D(n4521), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[246][2]  (.Q(\ram[246][2] ), 
	.D(n4520), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[246][1]  (.Q(\ram[246][1] ), 
	.D(n4519), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][0]  (.Q(\ram[246][0] ), 
	.D(n4518), 
	.CK(clk));
   QDFFEHD \ram_reg[242][15]  (.Q(\ram[242][15] ), 
	.D(n4469), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[242][14]  (.Q(\ram[242][14] ), 
	.D(n4468), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][13]  (.Q(\ram[242][13] ), 
	.D(n4467), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][12]  (.Q(\ram[242][12] ), 
	.D(n4466), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][11]  (.Q(\ram[242][11] ), 
	.D(n4465), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][10]  (.Q(\ram[242][10] ), 
	.D(n4464), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][9]  (.Q(\ram[242][9] ), 
	.D(n4463), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][8]  (.Q(\ram[242][8] ), 
	.D(n4462), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][7]  (.Q(\ram[242][7] ), 
	.D(n4461), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][6]  (.Q(\ram[242][6] ), 
	.D(n4460), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][5]  (.Q(\ram[242][5] ), 
	.D(n4459), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][4]  (.Q(\ram[242][4] ), 
	.D(n4458), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][3]  (.Q(\ram[242][3] ), 
	.D(n4457), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][2]  (.Q(\ram[242][2] ), 
	.D(n4456), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][1]  (.Q(\ram[242][1] ), 
	.D(n4455), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][0]  (.Q(\ram[242][0] ), 
	.D(n4454), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[238][15]  (.Q(\ram[238][15] ), 
	.D(n4405), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][14]  (.Q(\ram[238][14] ), 
	.D(n4404), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][13]  (.Q(\ram[238][13] ), 
	.D(n4403), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][12]  (.Q(\ram[238][12] ), 
	.D(n4402), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][11]  (.Q(\ram[238][11] ), 
	.D(n4401), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][10]  (.Q(\ram[238][10] ), 
	.D(n4400), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[238][9]  (.Q(\ram[238][9] ), 
	.D(n4399), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[238][8]  (.Q(\ram[238][8] ), 
	.D(n4398), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][7]  (.Q(\ram[238][7] ), 
	.D(n4397), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[238][6]  (.Q(\ram[238][6] ), 
	.D(n4396), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][5]  (.Q(\ram[238][5] ), 
	.D(n4395), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[238][4]  (.Q(\ram[238][4] ), 
	.D(n4394), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][3]  (.Q(\ram[238][3] ), 
	.D(n4393), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[238][2]  (.Q(\ram[238][2] ), 
	.D(n4392), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][1]  (.Q(\ram[238][1] ), 
	.D(n4391), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[238][0]  (.Q(\ram[238][0] ), 
	.D(n4390), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[234][15]  (.Q(\ram[234][15] ), 
	.D(n4341), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[234][14]  (.Q(\ram[234][14] ), 
	.D(n4340), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[234][13]  (.Q(\ram[234][13] ), 
	.D(n4339), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[234][12]  (.Q(\ram[234][12] ), 
	.D(n4338), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[234][11]  (.Q(\ram[234][11] ), 
	.D(n4337), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][10]  (.Q(\ram[234][10] ), 
	.D(n4336), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][9]  (.Q(\ram[234][9] ), 
	.D(n4335), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][8]  (.Q(\ram[234][8] ), 
	.D(n4334), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][7]  (.Q(\ram[234][7] ), 
	.D(n4333), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][6]  (.Q(\ram[234][6] ), 
	.D(n4332), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[234][5]  (.Q(\ram[234][5] ), 
	.D(n4331), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[234][4]  (.Q(\ram[234][4] ), 
	.D(n4330), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[234][3]  (.Q(\ram[234][3] ), 
	.D(n4329), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[234][2]  (.Q(\ram[234][2] ), 
	.D(n4328), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][1]  (.Q(\ram[234][1] ), 
	.D(n4327), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[234][0]  (.Q(\ram[234][0] ), 
	.D(n4326), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[230][15]  (.Q(\ram[230][15] ), 
	.D(n4277), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[230][14]  (.Q(\ram[230][14] ), 
	.D(n4276), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[230][13]  (.Q(\ram[230][13] ), 
	.D(n4275), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[230][12]  (.Q(\ram[230][12] ), 
	.D(n4274), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[230][11]  (.Q(\ram[230][11] ), 
	.D(n4273), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][10]  (.Q(\ram[230][10] ), 
	.D(n4272), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][9]  (.Q(\ram[230][9] ), 
	.D(n4271), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][8]  (.Q(\ram[230][8] ), 
	.D(n4270), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][7]  (.Q(\ram[230][7] ), 
	.D(n4269), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][6]  (.Q(\ram[230][6] ), 
	.D(n4268), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[230][5]  (.Q(\ram[230][5] ), 
	.D(n4267), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[230][4]  (.Q(\ram[230][4] ), 
	.D(n4266), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][3]  (.Q(\ram[230][3] ), 
	.D(n4265), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[230][2]  (.Q(\ram[230][2] ), 
	.D(n4264), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[230][1]  (.Q(\ram[230][1] ), 
	.D(n4263), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[230][0]  (.Q(\ram[230][0] ), 
	.D(n4262), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[226][15]  (.Q(\ram[226][15] ), 
	.D(n4213), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][14]  (.Q(\ram[226][14] ), 
	.D(n4212), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][13]  (.Q(\ram[226][13] ), 
	.D(n4211), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[226][12]  (.Q(\ram[226][12] ), 
	.D(n4210), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[226][11]  (.Q(\ram[226][11] ), 
	.D(n4209), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][10]  (.Q(\ram[226][10] ), 
	.D(n4208), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[226][9]  (.Q(\ram[226][9] ), 
	.D(n4207), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][8]  (.Q(\ram[226][8] ), 
	.D(n4206), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][7]  (.Q(\ram[226][7] ), 
	.D(n4205), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[226][6]  (.Q(\ram[226][6] ), 
	.D(n4204), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[226][5]  (.Q(\ram[226][5] ), 
	.D(n4203), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][4]  (.Q(\ram[226][4] ), 
	.D(n4202), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][3]  (.Q(\ram[226][3] ), 
	.D(n4201), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][2]  (.Q(\ram[226][2] ), 
	.D(n4200), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[226][1]  (.Q(\ram[226][1] ), 
	.D(n4199), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][0]  (.Q(\ram[226][0] ), 
	.D(n4198), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[222][15]  (.Q(\ram[222][15] ), 
	.D(n4149), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[222][14]  (.Q(\ram[222][14] ), 
	.D(n4148), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[222][13]  (.Q(\ram[222][13] ), 
	.D(n4147), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][12]  (.Q(\ram[222][12] ), 
	.D(n4146), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][11]  (.Q(\ram[222][11] ), 
	.D(n4145), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[222][10]  (.Q(\ram[222][10] ), 
	.D(n4144), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[222][9]  (.Q(\ram[222][9] ), 
	.D(n4143), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][8]  (.Q(\ram[222][8] ), 
	.D(n4142), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][7]  (.Q(\ram[222][7] ), 
	.D(n4141), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][6]  (.Q(\ram[222][6] ), 
	.D(n4140), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][5]  (.Q(\ram[222][5] ), 
	.D(n4139), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][4]  (.Q(\ram[222][4] ), 
	.D(n4138), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[222][3]  (.Q(\ram[222][3] ), 
	.D(n4137), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][2]  (.Q(\ram[222][2] ), 
	.D(n4136), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[222][1]  (.Q(\ram[222][1] ), 
	.D(n4135), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][0]  (.Q(\ram[222][0] ), 
	.D(n4134), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[218][15]  (.Q(\ram[218][15] ), 
	.D(n4085), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][14]  (.Q(\ram[218][14] ), 
	.D(n4084), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][13]  (.Q(\ram[218][13] ), 
	.D(n4083), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][12]  (.Q(\ram[218][12] ), 
	.D(n4082), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[218][11]  (.Q(\ram[218][11] ), 
	.D(n4081), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][10]  (.Q(\ram[218][10] ), 
	.D(n4080), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][9]  (.Q(\ram[218][9] ), 
	.D(n4079), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[218][8]  (.Q(\ram[218][8] ), 
	.D(n4078), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[218][7]  (.Q(\ram[218][7] ), 
	.D(n4077), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][6]  (.Q(\ram[218][6] ), 
	.D(n4076), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][5]  (.Q(\ram[218][5] ), 
	.D(n4075), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][4]  (.Q(\ram[218][4] ), 
	.D(n4074), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[218][3]  (.Q(\ram[218][3] ), 
	.D(n4073), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[218][2]  (.Q(\ram[218][2] ), 
	.D(n4072), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][1]  (.Q(\ram[218][1] ), 
	.D(n4071), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][0]  (.Q(\ram[218][0] ), 
	.D(n4070), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[214][15]  (.Q(\ram[214][15] ), 
	.D(n4021), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][14]  (.Q(\ram[214][14] ), 
	.D(n4020), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][13]  (.Q(\ram[214][13] ), 
	.D(n4019), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][12]  (.Q(\ram[214][12] ), 
	.D(n4018), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][11]  (.Q(\ram[214][11] ), 
	.D(n4017), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][10]  (.Q(\ram[214][10] ), 
	.D(n4016), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][9]  (.Q(\ram[214][9] ), 
	.D(n4015), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][8]  (.Q(\ram[214][8] ), 
	.D(n4014), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][7]  (.Q(\ram[214][7] ), 
	.D(n4013), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][6]  (.Q(\ram[214][6] ), 
	.D(n4012), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][5]  (.Q(\ram[214][5] ), 
	.D(n4011), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][4]  (.Q(\ram[214][4] ), 
	.D(n4010), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[214][3]  (.Q(\ram[214][3] ), 
	.D(n4009), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][2]  (.Q(\ram[214][2] ), 
	.D(n4008), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][1]  (.Q(\ram[214][1] ), 
	.D(n4007), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][0]  (.Q(\ram[214][0] ), 
	.D(n4006), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[210][15]  (.Q(\ram[210][15] ), 
	.D(n3957), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[210][14]  (.Q(\ram[210][14] ), 
	.D(n3956), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[210][13]  (.Q(\ram[210][13] ), 
	.D(n3955), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][12]  (.Q(\ram[210][12] ), 
	.D(n3954), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][11]  (.Q(\ram[210][11] ), 
	.D(n3953), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][10]  (.Q(\ram[210][10] ), 
	.D(n3952), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][9]  (.Q(\ram[210][9] ), 
	.D(n3951), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][8]  (.Q(\ram[210][8] ), 
	.D(n3950), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][7]  (.Q(\ram[210][7] ), 
	.D(n3949), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][6]  (.Q(\ram[210][6] ), 
	.D(n3948), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][5]  (.Q(\ram[210][5] ), 
	.D(n3947), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][4]  (.Q(\ram[210][4] ), 
	.D(n3946), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[210][3]  (.Q(\ram[210][3] ), 
	.D(n3945), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[210][2]  (.Q(\ram[210][2] ), 
	.D(n3944), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][1]  (.Q(\ram[210][1] ), 
	.D(n3943), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[210][0]  (.Q(\ram[210][0] ), 
	.D(n3942), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[206][15]  (.Q(\ram[206][15] ), 
	.D(n3893), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][14]  (.Q(\ram[206][14] ), 
	.D(n3892), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[206][13]  (.Q(\ram[206][13] ), 
	.D(n3891), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[206][12]  (.Q(\ram[206][12] ), 
	.D(n3890), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[206][11]  (.Q(\ram[206][11] ), 
	.D(n3889), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][10]  (.Q(\ram[206][10] ), 
	.D(n3888), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[206][9]  (.Q(\ram[206][9] ), 
	.D(n3887), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[206][8]  (.Q(\ram[206][8] ), 
	.D(n3886), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[206][7]  (.Q(\ram[206][7] ), 
	.D(n3885), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[206][6]  (.Q(\ram[206][6] ), 
	.D(n3884), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[206][5]  (.Q(\ram[206][5] ), 
	.D(n3883), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[206][4]  (.Q(\ram[206][4] ), 
	.D(n3882), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][3]  (.Q(\ram[206][3] ), 
	.D(n3881), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[206][2]  (.Q(\ram[206][2] ), 
	.D(n3880), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][1]  (.Q(\ram[206][1] ), 
	.D(n3879), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[206][0]  (.Q(\ram[206][0] ), 
	.D(n3878), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[202][15]  (.Q(\ram[202][15] ), 
	.D(n3829), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][14]  (.Q(\ram[202][14] ), 
	.D(n3828), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][13]  (.Q(\ram[202][13] ), 
	.D(n3827), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[202][12]  (.Q(\ram[202][12] ), 
	.D(n3826), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][11]  (.Q(\ram[202][11] ), 
	.D(n3825), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][10]  (.Q(\ram[202][10] ), 
	.D(n3824), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][9]  (.Q(\ram[202][9] ), 
	.D(n3823), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][8]  (.Q(\ram[202][8] ), 
	.D(n3822), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[202][7]  (.Q(\ram[202][7] ), 
	.D(n3821), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][6]  (.Q(\ram[202][6] ), 
	.D(n3820), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[202][5]  (.Q(\ram[202][5] ), 
	.D(n3819), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[202][4]  (.Q(\ram[202][4] ), 
	.D(n3818), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][3]  (.Q(\ram[202][3] ), 
	.D(n3817), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][2]  (.Q(\ram[202][2] ), 
	.D(n3816), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][1]  (.Q(\ram[202][1] ), 
	.D(n3815), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][0]  (.Q(\ram[202][0] ), 
	.D(n3814), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[198][15]  (.Q(\ram[198][15] ), 
	.D(n3765), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][14]  (.Q(\ram[198][14] ), 
	.D(n3764), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][13]  (.Q(\ram[198][13] ), 
	.D(n3763), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][12]  (.Q(\ram[198][12] ), 
	.D(n3762), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][11]  (.Q(\ram[198][11] ), 
	.D(n3761), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][10]  (.Q(\ram[198][10] ), 
	.D(n3760), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][9]  (.Q(\ram[198][9] ), 
	.D(n3759), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[198][8]  (.Q(\ram[198][8] ), 
	.D(n3758), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][7]  (.Q(\ram[198][7] ), 
	.D(n3757), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][6]  (.Q(\ram[198][6] ), 
	.D(n3756), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][5]  (.Q(\ram[198][5] ), 
	.D(n3755), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][4]  (.Q(\ram[198][4] ), 
	.D(n3754), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][3]  (.Q(\ram[198][3] ), 
	.D(n3753), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[198][2]  (.Q(\ram[198][2] ), 
	.D(n3752), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][1]  (.Q(\ram[198][1] ), 
	.D(n3751), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][0]  (.Q(\ram[198][0] ), 
	.D(n3750), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[194][15]  (.Q(\ram[194][15] ), 
	.D(n3701), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][14]  (.Q(\ram[194][14] ), 
	.D(n3700), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][13]  (.Q(\ram[194][13] ), 
	.D(n3699), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[194][12]  (.Q(\ram[194][12] ), 
	.D(n3698), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][11]  (.Q(\ram[194][11] ), 
	.D(n3697), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][10]  (.Q(\ram[194][10] ), 
	.D(n3696), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[194][9]  (.Q(\ram[194][9] ), 
	.D(n3695), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][8]  (.Q(\ram[194][8] ), 
	.D(n3694), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[194][7]  (.Q(\ram[194][7] ), 
	.D(n3693), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][6]  (.Q(\ram[194][6] ), 
	.D(n3692), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][5]  (.Q(\ram[194][5] ), 
	.D(n3691), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][4]  (.Q(\ram[194][4] ), 
	.D(n3690), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][3]  (.Q(\ram[194][3] ), 
	.D(n3689), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[194][2]  (.Q(\ram[194][2] ), 
	.D(n3688), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][1]  (.Q(\ram[194][1] ), 
	.D(n3687), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][0]  (.Q(\ram[194][0] ), 
	.D(n3686), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[190][15]  (.Q(\ram[190][15] ), 
	.D(n3637), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][14]  (.Q(\ram[190][14] ), 
	.D(n3636), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][13]  (.Q(\ram[190][13] ), 
	.D(n3635), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[190][12]  (.Q(\ram[190][12] ), 
	.D(n3634), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[190][11]  (.Q(\ram[190][11] ), 
	.D(n3633), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][10]  (.Q(\ram[190][10] ), 
	.D(n3632), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][9]  (.Q(\ram[190][9] ), 
	.D(n3631), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][8]  (.Q(\ram[190][8] ), 
	.D(n3630), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][7]  (.Q(\ram[190][7] ), 
	.D(n3629), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][6]  (.Q(\ram[190][6] ), 
	.D(n3628), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[190][5]  (.Q(\ram[190][5] ), 
	.D(n3627), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[190][4]  (.Q(\ram[190][4] ), 
	.D(n3626), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][3]  (.Q(\ram[190][3] ), 
	.D(n3625), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[190][2]  (.Q(\ram[190][2] ), 
	.D(n3624), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][1]  (.Q(\ram[190][1] ), 
	.D(n3623), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][0]  (.Q(\ram[190][0] ), 
	.D(n3622), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[186][15]  (.Q(\ram[186][15] ), 
	.D(n3573), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][14]  (.Q(\ram[186][14] ), 
	.D(n3572), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][13]  (.Q(\ram[186][13] ), 
	.D(n3571), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][12]  (.Q(\ram[186][12] ), 
	.D(n3570), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[186][11]  (.Q(\ram[186][11] ), 
	.D(n3569), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][10]  (.Q(\ram[186][10] ), 
	.D(n3568), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[186][9]  (.Q(\ram[186][9] ), 
	.D(n3567), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[186][8]  (.Q(\ram[186][8] ), 
	.D(n3566), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[186][7]  (.Q(\ram[186][7] ), 
	.D(n3565), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][6]  (.Q(\ram[186][6] ), 
	.D(n3564), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][5]  (.Q(\ram[186][5] ), 
	.D(n3563), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][4]  (.Q(\ram[186][4] ), 
	.D(n3562), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[186][3]  (.Q(\ram[186][3] ), 
	.D(n3561), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][2]  (.Q(\ram[186][2] ), 
	.D(n3560), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][1]  (.Q(\ram[186][1] ), 
	.D(n3559), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][0]  (.Q(\ram[186][0] ), 
	.D(n3558), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[182][15]  (.Q(\ram[182][15] ), 
	.D(n3509), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[182][14]  (.Q(\ram[182][14] ), 
	.D(n3508), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[182][13]  (.Q(\ram[182][13] ), 
	.D(n3507), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[182][12]  (.Q(\ram[182][12] ), 
	.D(n3506), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[182][11]  (.Q(\ram[182][11] ), 
	.D(n3505), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[182][10]  (.Q(\ram[182][10] ), 
	.D(n3504), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[182][9]  (.Q(\ram[182][9] ), 
	.D(n3503), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[182][8]  (.Q(\ram[182][8] ), 
	.D(n3502), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[182][7]  (.Q(\ram[182][7] ), 
	.D(n3501), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[182][6]  (.Q(\ram[182][6] ), 
	.D(n3500), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[182][5]  (.Q(\ram[182][5] ), 
	.D(n3499), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[182][4]  (.Q(\ram[182][4] ), 
	.D(n3498), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[182][3]  (.Q(\ram[182][3] ), 
	.D(n3497), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[182][2]  (.Q(\ram[182][2] ), 
	.D(n3496), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[182][1]  (.Q(\ram[182][1] ), 
	.D(n3495), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[182][0]  (.Q(\ram[182][0] ), 
	.D(n3494), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[178][15]  (.Q(\ram[178][15] ), 
	.D(n3445), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][14]  (.Q(\ram[178][14] ), 
	.D(n3444), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][13]  (.Q(\ram[178][13] ), 
	.D(n3443), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][12]  (.Q(\ram[178][12] ), 
	.D(n3442), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][11]  (.Q(\ram[178][11] ), 
	.D(n3441), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][10]  (.Q(\ram[178][10] ), 
	.D(n3440), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[178][9]  (.Q(\ram[178][9] ), 
	.D(n3439), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][8]  (.Q(\ram[178][8] ), 
	.D(n3438), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][7]  (.Q(\ram[178][7] ), 
	.D(n3437), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][6]  (.Q(\ram[178][6] ), 
	.D(n3436), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][5]  (.Q(\ram[178][5] ), 
	.D(n3435), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][4]  (.Q(\ram[178][4] ), 
	.D(n3434), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][3]  (.Q(\ram[178][3] ), 
	.D(n3433), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][2]  (.Q(\ram[178][2] ), 
	.D(n3432), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][1]  (.Q(\ram[178][1] ), 
	.D(n3431), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][0]  (.Q(\ram[178][0] ), 
	.D(n3430), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[174][15]  (.Q(\ram[174][15] ), 
	.D(n3381), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][14]  (.Q(\ram[174][14] ), 
	.D(n3380), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][13]  (.Q(\ram[174][13] ), 
	.D(n3379), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[174][12]  (.Q(\ram[174][12] ), 
	.D(n3378), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[174][11]  (.Q(\ram[174][11] ), 
	.D(n3377), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[174][10]  (.Q(\ram[174][10] ), 
	.D(n3376), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[174][9]  (.Q(\ram[174][9] ), 
	.D(n3375), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][8]  (.Q(\ram[174][8] ), 
	.D(n3374), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][7]  (.Q(\ram[174][7] ), 
	.D(n3373), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][6]  (.Q(\ram[174][6] ), 
	.D(n3372), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[174][5]  (.Q(\ram[174][5] ), 
	.D(n3371), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][4]  (.Q(\ram[174][4] ), 
	.D(n3370), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][3]  (.Q(\ram[174][3] ), 
	.D(n3369), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][2]  (.Q(\ram[174][2] ), 
	.D(n3368), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][1]  (.Q(\ram[174][1] ), 
	.D(n3367), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][0]  (.Q(\ram[174][0] ), 
	.D(n3366), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[170][15]  (.Q(\ram[170][15] ), 
	.D(n3317), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][14]  (.Q(\ram[170][14] ), 
	.D(n3316), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][13]  (.Q(\ram[170][13] ), 
	.D(n3315), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][12]  (.Q(\ram[170][12] ), 
	.D(n3314), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][11]  (.Q(\ram[170][11] ), 
	.D(n3313), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][10]  (.Q(\ram[170][10] ), 
	.D(n3312), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][9]  (.Q(\ram[170][9] ), 
	.D(n3311), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][8]  (.Q(\ram[170][8] ), 
	.D(n3310), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][7]  (.Q(\ram[170][7] ), 
	.D(n3309), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][6]  (.Q(\ram[170][6] ), 
	.D(n3308), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][5]  (.Q(\ram[170][5] ), 
	.D(n3307), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][4]  (.Q(\ram[170][4] ), 
	.D(n3306), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][3]  (.Q(\ram[170][3] ), 
	.D(n3305), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][2]  (.Q(\ram[170][2] ), 
	.D(n3304), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][1]  (.Q(\ram[170][1] ), 
	.D(n3303), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][0]  (.Q(\ram[170][0] ), 
	.D(n3302), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[166][15]  (.Q(\ram[166][15] ), 
	.D(n3253), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[166][14]  (.Q(\ram[166][14] ), 
	.D(n3252), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][13]  (.Q(\ram[166][13] ), 
	.D(n3251), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[166][12]  (.Q(\ram[166][12] ), 
	.D(n3250), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][11]  (.Q(\ram[166][11] ), 
	.D(n3249), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][10]  (.Q(\ram[166][10] ), 
	.D(n3248), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[166][9]  (.Q(\ram[166][9] ), 
	.D(n3247), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][8]  (.Q(\ram[166][8] ), 
	.D(n3246), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][7]  (.Q(\ram[166][7] ), 
	.D(n3245), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[166][6]  (.Q(\ram[166][6] ), 
	.D(n3244), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][5]  (.Q(\ram[166][5] ), 
	.D(n3243), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][4]  (.Q(\ram[166][4] ), 
	.D(n3242), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[166][3]  (.Q(\ram[166][3] ), 
	.D(n3241), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][2]  (.Q(\ram[166][2] ), 
	.D(n3240), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][1]  (.Q(\ram[166][1] ), 
	.D(n3239), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][0]  (.Q(\ram[166][0] ), 
	.D(n3238), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][15]  (.Q(\ram[162][15] ), 
	.D(n3189), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][14]  (.Q(\ram[162][14] ), 
	.D(n3188), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][13]  (.Q(\ram[162][13] ), 
	.D(n3187), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][12]  (.Q(\ram[162][12] ), 
	.D(n3186), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][11]  (.Q(\ram[162][11] ), 
	.D(n3185), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][10]  (.Q(\ram[162][10] ), 
	.D(n3184), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][9]  (.Q(\ram[162][9] ), 
	.D(n3183), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][8]  (.Q(\ram[162][8] ), 
	.D(n3182), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[162][7]  (.Q(\ram[162][7] ), 
	.D(n3181), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][6]  (.Q(\ram[162][6] ), 
	.D(n3180), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][5]  (.Q(\ram[162][5] ), 
	.D(n3179), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][4]  (.Q(\ram[162][4] ), 
	.D(n3178), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][3]  (.Q(\ram[162][3] ), 
	.D(n3177), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[162][2]  (.Q(\ram[162][2] ), 
	.D(n3176), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][1]  (.Q(\ram[162][1] ), 
	.D(n3175), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][0]  (.Q(\ram[162][0] ), 
	.D(n3174), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[158][15]  (.Q(\ram[158][15] ), 
	.D(n3125), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][14]  (.Q(\ram[158][14] ), 
	.D(n3124), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][13]  (.Q(\ram[158][13] ), 
	.D(n3123), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][12]  (.Q(\ram[158][12] ), 
	.D(n3122), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[158][11]  (.Q(\ram[158][11] ), 
	.D(n3121), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][10]  (.Q(\ram[158][10] ), 
	.D(n3120), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[158][9]  (.Q(\ram[158][9] ), 
	.D(n3119), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][8]  (.Q(\ram[158][8] ), 
	.D(n3118), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[158][7]  (.Q(\ram[158][7] ), 
	.D(n3117), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[158][6]  (.Q(\ram[158][6] ), 
	.D(n3116), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[158][5]  (.Q(\ram[158][5] ), 
	.D(n3115), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[158][4]  (.Q(\ram[158][4] ), 
	.D(n3114), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[158][3]  (.Q(\ram[158][3] ), 
	.D(n3113), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[158][2]  (.Q(\ram[158][2] ), 
	.D(n3112), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[158][1]  (.Q(\ram[158][1] ), 
	.D(n3111), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[158][0]  (.Q(\ram[158][0] ), 
	.D(n3110), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[154][15]  (.Q(\ram[154][15] ), 
	.D(n3061), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[154][14]  (.Q(\ram[154][14] ), 
	.D(n3060), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[154][13]  (.Q(\ram[154][13] ), 
	.D(n3059), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[154][12]  (.Q(\ram[154][12] ), 
	.D(n3058), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[154][11]  (.Q(\ram[154][11] ), 
	.D(n3057), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[154][10]  (.Q(\ram[154][10] ), 
	.D(n3056), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[154][9]  (.Q(\ram[154][9] ), 
	.D(n3055), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[154][8]  (.Q(\ram[154][8] ), 
	.D(n3054), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[154][7]  (.Q(\ram[154][7] ), 
	.D(n3053), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][6]  (.Q(\ram[154][6] ), 
	.D(n3052), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][5]  (.Q(\ram[154][5] ), 
	.D(n3051), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][4]  (.Q(\ram[154][4] ), 
	.D(n3050), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[154][3]  (.Q(\ram[154][3] ), 
	.D(n3049), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][2]  (.Q(\ram[154][2] ), 
	.D(n3048), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[154][1]  (.Q(\ram[154][1] ), 
	.D(n3047), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][0]  (.Q(\ram[154][0] ), 
	.D(n3046), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[150][15]  (.Q(\ram[150][15] ), 
	.D(n2997), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][14]  (.Q(\ram[150][14] ), 
	.D(n2996), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][13]  (.Q(\ram[150][13] ), 
	.D(n2995), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][12]  (.Q(\ram[150][12] ), 
	.D(n2994), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][11]  (.Q(\ram[150][11] ), 
	.D(n2993), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][10]  (.Q(\ram[150][10] ), 
	.D(n2992), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[150][9]  (.Q(\ram[150][9] ), 
	.D(n2991), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][8]  (.Q(\ram[150][8] ), 
	.D(n2990), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[150][7]  (.Q(\ram[150][7] ), 
	.D(n2989), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][6]  (.Q(\ram[150][6] ), 
	.D(n2988), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[150][5]  (.Q(\ram[150][5] ), 
	.D(n2987), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][4]  (.Q(\ram[150][4] ), 
	.D(n2986), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[150][3]  (.Q(\ram[150][3] ), 
	.D(n2985), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][2]  (.Q(\ram[150][2] ), 
	.D(n2984), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[150][1]  (.Q(\ram[150][1] ), 
	.D(n2983), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][0]  (.Q(\ram[150][0] ), 
	.D(n2982), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[146][15]  (.Q(\ram[146][15] ), 
	.D(n2933), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[146][14]  (.Q(\ram[146][14] ), 
	.D(n2932), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[146][13]  (.Q(\ram[146][13] ), 
	.D(n2931), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[146][12]  (.Q(\ram[146][12] ), 
	.D(n2930), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[146][11]  (.Q(\ram[146][11] ), 
	.D(n2929), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[146][10]  (.Q(\ram[146][10] ), 
	.D(n2928), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[146][9]  (.Q(\ram[146][9] ), 
	.D(n2927), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[146][8]  (.Q(\ram[146][8] ), 
	.D(n2926), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[146][7]  (.Q(\ram[146][7] ), 
	.D(n2925), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[146][6]  (.Q(\ram[146][6] ), 
	.D(n2924), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][5]  (.Q(\ram[146][5] ), 
	.D(n2923), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][4]  (.Q(\ram[146][4] ), 
	.D(n2922), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[146][3]  (.Q(\ram[146][3] ), 
	.D(n2921), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][2]  (.Q(\ram[146][2] ), 
	.D(n2920), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[146][1]  (.Q(\ram[146][1] ), 
	.D(n2919), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][0]  (.Q(\ram[146][0] ), 
	.D(n2918), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[142][15]  (.Q(\ram[142][15] ), 
	.D(n2869), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[142][14]  (.Q(\ram[142][14] ), 
	.D(n2868), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[142][13]  (.Q(\ram[142][13] ), 
	.D(n2867), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[142][12]  (.Q(\ram[142][12] ), 
	.D(n2866), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[142][11]  (.Q(\ram[142][11] ), 
	.D(n2865), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[142][10]  (.Q(\ram[142][10] ), 
	.D(n2864), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[142][9]  (.Q(\ram[142][9] ), 
	.D(n2863), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[142][8]  (.Q(\ram[142][8] ), 
	.D(n2862), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[142][7]  (.Q(\ram[142][7] ), 
	.D(n2861), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[142][6]  (.Q(\ram[142][6] ), 
	.D(n2860), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[142][5]  (.Q(\ram[142][5] ), 
	.D(n2859), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[142][4]  (.Q(\ram[142][4] ), 
	.D(n2858), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[142][3]  (.Q(\ram[142][3] ), 
	.D(n2857), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[142][2]  (.Q(\ram[142][2] ), 
	.D(n2856), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[142][1]  (.Q(\ram[142][1] ), 
	.D(n2855), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[142][0]  (.Q(\ram[142][0] ), 
	.D(n2854), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[138][15]  (.Q(\ram[138][15] ), 
	.D(n2805), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][14]  (.Q(\ram[138][14] ), 
	.D(n2804), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][13]  (.Q(\ram[138][13] ), 
	.D(n2803), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[138][12]  (.Q(\ram[138][12] ), 
	.D(n2802), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][11]  (.Q(\ram[138][11] ), 
	.D(n2801), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][10]  (.Q(\ram[138][10] ), 
	.D(n2800), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][9]  (.Q(\ram[138][9] ), 
	.D(n2799), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][8]  (.Q(\ram[138][8] ), 
	.D(n2798), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[138][7]  (.Q(\ram[138][7] ), 
	.D(n2797), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][6]  (.Q(\ram[138][6] ), 
	.D(n2796), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][5]  (.Q(\ram[138][5] ), 
	.D(n2795), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][4]  (.Q(\ram[138][4] ), 
	.D(n2794), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][3]  (.Q(\ram[138][3] ), 
	.D(n2793), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][2]  (.Q(\ram[138][2] ), 
	.D(n2792), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][1]  (.Q(\ram[138][1] ), 
	.D(n2791), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][0]  (.Q(\ram[138][0] ), 
	.D(n2790), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[134][15]  (.Q(\ram[134][15] ), 
	.D(n2741), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[134][14]  (.Q(\ram[134][14] ), 
	.D(n2740), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[134][13]  (.Q(\ram[134][13] ), 
	.D(n2739), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[134][12]  (.Q(\ram[134][12] ), 
	.D(n2738), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][11]  (.Q(\ram[134][11] ), 
	.D(n2737), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[134][10]  (.Q(\ram[134][10] ), 
	.D(n2736), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][9]  (.Q(\ram[134][9] ), 
	.D(n2735), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[134][8]  (.Q(\ram[134][8] ), 
	.D(n2734), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[134][7]  (.Q(\ram[134][7] ), 
	.D(n2733), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][6]  (.Q(\ram[134][6] ), 
	.D(n2732), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][5]  (.Q(\ram[134][5] ), 
	.D(n2731), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][4]  (.Q(\ram[134][4] ), 
	.D(n2730), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[134][3]  (.Q(\ram[134][3] ), 
	.D(n2729), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][2]  (.Q(\ram[134][2] ), 
	.D(n2728), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][1]  (.Q(\ram[134][1] ), 
	.D(n2727), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][0]  (.Q(\ram[134][0] ), 
	.D(n2726), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[130][15]  (.Q(\ram[130][15] ), 
	.D(n2677), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][14]  (.Q(\ram[130][14] ), 
	.D(n2676), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][13]  (.Q(\ram[130][13] ), 
	.D(n2675), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][12]  (.Q(\ram[130][12] ), 
	.D(n2674), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][11]  (.Q(\ram[130][11] ), 
	.D(n2673), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[130][10]  (.Q(\ram[130][10] ), 
	.D(n2672), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[130][9]  (.Q(\ram[130][9] ), 
	.D(n2671), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][8]  (.Q(\ram[130][8] ), 
	.D(n2670), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[130][7]  (.Q(\ram[130][7] ), 
	.D(n2669), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[130][6]  (.Q(\ram[130][6] ), 
	.D(n2668), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[130][5]  (.Q(\ram[130][5] ), 
	.D(n2667), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[130][4]  (.Q(\ram[130][4] ), 
	.D(n2666), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[130][3]  (.Q(\ram[130][3] ), 
	.D(n2665), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[130][2]  (.Q(\ram[130][2] ), 
	.D(n2664), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[130][1]  (.Q(\ram[130][1] ), 
	.D(n2663), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[130][0]  (.Q(\ram[130][0] ), 
	.D(n2662), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[126][15]  (.Q(\ram[126][15] ), 
	.D(n2613), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][14]  (.Q(\ram[126][14] ), 
	.D(n2612), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][13]  (.Q(\ram[126][13] ), 
	.D(n2611), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][12]  (.Q(\ram[126][12] ), 
	.D(n2610), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][11]  (.Q(\ram[126][11] ), 
	.D(n2609), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][10]  (.Q(\ram[126][10] ), 
	.D(n2608), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][9]  (.Q(\ram[126][9] ), 
	.D(n2607), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][8]  (.Q(\ram[126][8] ), 
	.D(n2606), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][7]  (.Q(\ram[126][7] ), 
	.D(n2605), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[126][6]  (.Q(\ram[126][6] ), 
	.D(n2604), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[126][5]  (.Q(\ram[126][5] ), 
	.D(n2603), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[126][4]  (.Q(\ram[126][4] ), 
	.D(n2602), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[126][3]  (.Q(\ram[126][3] ), 
	.D(n2601), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[126][2]  (.Q(\ram[126][2] ), 
	.D(n2600), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][1]  (.Q(\ram[126][1] ), 
	.D(n2599), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][0]  (.Q(\ram[126][0] ), 
	.D(n2598), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[122][15]  (.Q(\ram[122][15] ), 
	.D(n2549), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][14]  (.Q(\ram[122][14] ), 
	.D(n2548), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][13]  (.Q(\ram[122][13] ), 
	.D(n2547), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[122][12]  (.Q(\ram[122][12] ), 
	.D(n2546), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][11]  (.Q(\ram[122][11] ), 
	.D(n2545), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][10]  (.Q(\ram[122][10] ), 
	.D(n2544), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][9]  (.Q(\ram[122][9] ), 
	.D(n2543), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][8]  (.Q(\ram[122][8] ), 
	.D(n2542), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][7]  (.Q(\ram[122][7] ), 
	.D(n2541), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][6]  (.Q(\ram[122][6] ), 
	.D(n2540), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[122][5]  (.Q(\ram[122][5] ), 
	.D(n2539), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[122][4]  (.Q(\ram[122][4] ), 
	.D(n2538), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[122][3]  (.Q(\ram[122][3] ), 
	.D(n2537), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[122][2]  (.Q(\ram[122][2] ), 
	.D(n2536), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][1]  (.Q(\ram[122][1] ), 
	.D(n2535), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][0]  (.Q(\ram[122][0] ), 
	.D(n2534), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[118][15]  (.Q(\ram[118][15] ), 
	.D(n2485), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[118][14]  (.Q(\ram[118][14] ), 
	.D(n2484), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][13]  (.Q(\ram[118][13] ), 
	.D(n2483), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[118][12]  (.Q(\ram[118][12] ), 
	.D(n2482), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[118][11]  (.Q(\ram[118][11] ), 
	.D(n2481), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[118][10]  (.Q(\ram[118][10] ), 
	.D(n2480), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[118][9]  (.Q(\ram[118][9] ), 
	.D(n2479), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][8]  (.Q(\ram[118][8] ), 
	.D(n2478), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][7]  (.Q(\ram[118][7] ), 
	.D(n2477), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][6]  (.Q(\ram[118][6] ), 
	.D(n2476), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][5]  (.Q(\ram[118][5] ), 
	.D(n2475), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[118][4]  (.Q(\ram[118][4] ), 
	.D(n2474), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][3]  (.Q(\ram[118][3] ), 
	.D(n2473), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][2]  (.Q(\ram[118][2] ), 
	.D(n2472), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][1]  (.Q(\ram[118][1] ), 
	.D(n2471), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][0]  (.Q(\ram[118][0] ), 
	.D(n2470), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[114][15]  (.Q(\ram[114][15] ), 
	.D(n2421), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[114][14]  (.Q(\ram[114][14] ), 
	.D(n2420), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[114][13]  (.Q(\ram[114][13] ), 
	.D(n2419), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[114][12]  (.Q(\ram[114][12] ), 
	.D(n2418), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][11]  (.Q(\ram[114][11] ), 
	.D(n2417), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][10]  (.Q(\ram[114][10] ), 
	.D(n2416), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[114][9]  (.Q(\ram[114][9] ), 
	.D(n2415), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[114][8]  (.Q(\ram[114][8] ), 
	.D(n2414), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][7]  (.Q(\ram[114][7] ), 
	.D(n2413), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[114][6]  (.Q(\ram[114][6] ), 
	.D(n2412), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[114][5]  (.Q(\ram[114][5] ), 
	.D(n2411), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[114][4]  (.Q(\ram[114][4] ), 
	.D(n2410), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[114][3]  (.Q(\ram[114][3] ), 
	.D(n2409), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[114][2]  (.Q(\ram[114][2] ), 
	.D(n2408), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][1]  (.Q(\ram[114][1] ), 
	.D(n2407), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[114][0]  (.Q(\ram[114][0] ), 
	.D(n2406), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[110][15]  (.Q(\ram[110][15] ), 
	.D(n2357), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[110][14]  (.Q(\ram[110][14] ), 
	.D(n2356), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[110][13]  (.Q(\ram[110][13] ), 
	.D(n2355), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[110][12]  (.Q(\ram[110][12] ), 
	.D(n2354), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[110][11]  (.Q(\ram[110][11] ), 
	.D(n2353), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[110][10]  (.Q(\ram[110][10] ), 
	.D(n2352), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[110][9]  (.Q(\ram[110][9] ), 
	.D(n2351), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[110][8]  (.Q(\ram[110][8] ), 
	.D(n2350), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][7]  (.Q(\ram[110][7] ), 
	.D(n2349), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[110][6]  (.Q(\ram[110][6] ), 
	.D(n2348), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][5]  (.Q(\ram[110][5] ), 
	.D(n2347), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[110][4]  (.Q(\ram[110][4] ), 
	.D(n2346), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][3]  (.Q(\ram[110][3] ), 
	.D(n2345), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[110][2]  (.Q(\ram[110][2] ), 
	.D(n2344), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][1]  (.Q(\ram[110][1] ), 
	.D(n2343), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][0]  (.Q(\ram[110][0] ), 
	.D(n2342), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[106][15]  (.Q(\ram[106][15] ), 
	.D(n2293), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][14]  (.Q(\ram[106][14] ), 
	.D(n2292), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[106][13]  (.Q(\ram[106][13] ), 
	.D(n2291), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[106][12]  (.Q(\ram[106][12] ), 
	.D(n2290), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][11]  (.Q(\ram[106][11] ), 
	.D(n2289), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[106][10]  (.Q(\ram[106][10] ), 
	.D(n2288), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[106][9]  (.Q(\ram[106][9] ), 
	.D(n2287), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[106][8]  (.Q(\ram[106][8] ), 
	.D(n2286), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][7]  (.Q(\ram[106][7] ), 
	.D(n2285), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[106][6]  (.Q(\ram[106][6] ), 
	.D(n2284), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][5]  (.Q(\ram[106][5] ), 
	.D(n2283), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[106][4]  (.Q(\ram[106][4] ), 
	.D(n2282), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[106][3]  (.Q(\ram[106][3] ), 
	.D(n2281), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[106][2]  (.Q(\ram[106][2] ), 
	.D(n2280), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][1]  (.Q(\ram[106][1] ), 
	.D(n2279), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][0]  (.Q(\ram[106][0] ), 
	.D(n2278), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[102][15]  (.Q(\ram[102][15] ), 
	.D(n2229), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][14]  (.Q(\ram[102][14] ), 
	.D(n2228), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][13]  (.Q(\ram[102][13] ), 
	.D(n2227), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[102][12]  (.Q(\ram[102][12] ), 
	.D(n2226), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][11]  (.Q(\ram[102][11] ), 
	.D(n2225), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[102][10]  (.Q(\ram[102][10] ), 
	.D(n2224), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][9]  (.Q(\ram[102][9] ), 
	.D(n2223), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][8]  (.Q(\ram[102][8] ), 
	.D(n2222), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][7]  (.Q(\ram[102][7] ), 
	.D(n2221), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[102][6]  (.Q(\ram[102][6] ), 
	.D(n2220), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][5]  (.Q(\ram[102][5] ), 
	.D(n2219), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][4]  (.Q(\ram[102][4] ), 
	.D(n2218), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][3]  (.Q(\ram[102][3] ), 
	.D(n2217), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[102][2]  (.Q(\ram[102][2] ), 
	.D(n2216), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][1]  (.Q(\ram[102][1] ), 
	.D(n2215), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[102][0]  (.Q(\ram[102][0] ), 
	.D(n2214), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[98][15]  (.Q(\ram[98][15] ), 
	.D(n2165), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][14]  (.Q(\ram[98][14] ), 
	.D(n2164), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][13]  (.Q(\ram[98][13] ), 
	.D(n2163), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[98][12]  (.Q(\ram[98][12] ), 
	.D(n2162), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][11]  (.Q(\ram[98][11] ), 
	.D(n2161), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[98][10]  (.Q(\ram[98][10] ), 
	.D(n2160), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[98][9]  (.Q(\ram[98][9] ), 
	.D(n2159), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][8]  (.Q(\ram[98][8] ), 
	.D(n2158), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][7]  (.Q(\ram[98][7] ), 
	.D(n2157), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[98][6]  (.Q(\ram[98][6] ), 
	.D(n2156), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][5]  (.Q(\ram[98][5] ), 
	.D(n2155), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][4]  (.Q(\ram[98][4] ), 
	.D(n2154), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[98][3]  (.Q(\ram[98][3] ), 
	.D(n2153), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[98][2]  (.Q(\ram[98][2] ), 
	.D(n2152), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[98][1]  (.Q(\ram[98][1] ), 
	.D(n2151), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[98][0]  (.Q(\ram[98][0] ), 
	.D(n2150), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[94][15]  (.Q(\ram[94][15] ), 
	.D(n2101), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][14]  (.Q(\ram[94][14] ), 
	.D(n2100), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][13]  (.Q(\ram[94][13] ), 
	.D(n2099), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][12]  (.Q(\ram[94][12] ), 
	.D(n2098), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][11]  (.Q(\ram[94][11] ), 
	.D(n2097), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][10]  (.Q(\ram[94][10] ), 
	.D(n2096), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][9]  (.Q(\ram[94][9] ), 
	.D(n2095), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][8]  (.Q(\ram[94][8] ), 
	.D(n2094), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][7]  (.Q(\ram[94][7] ), 
	.D(n2093), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][6]  (.Q(\ram[94][6] ), 
	.D(n2092), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][5]  (.Q(\ram[94][5] ), 
	.D(n2091), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[94][4]  (.Q(\ram[94][4] ), 
	.D(n2090), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][3]  (.Q(\ram[94][3] ), 
	.D(n2089), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][2]  (.Q(\ram[94][2] ), 
	.D(n2088), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][1]  (.Q(\ram[94][1] ), 
	.D(n2087), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][0]  (.Q(\ram[94][0] ), 
	.D(n2086), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[90][15]  (.Q(\ram[90][15] ), 
	.D(n2037), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][14]  (.Q(\ram[90][14] ), 
	.D(n2036), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[90][13]  (.Q(\ram[90][13] ), 
	.D(n2035), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][12]  (.Q(\ram[90][12] ), 
	.D(n2034), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[90][11]  (.Q(\ram[90][11] ), 
	.D(n2033), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[90][10]  (.Q(\ram[90][10] ), 
	.D(n2032), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][9]  (.Q(\ram[90][9] ), 
	.D(n2031), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][8]  (.Q(\ram[90][8] ), 
	.D(n2030), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][7]  (.Q(\ram[90][7] ), 
	.D(n2029), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][6]  (.Q(\ram[90][6] ), 
	.D(n2028), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][5]  (.Q(\ram[90][5] ), 
	.D(n2027), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[90][4]  (.Q(\ram[90][4] ), 
	.D(n2026), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][3]  (.Q(\ram[90][3] ), 
	.D(n2025), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][2]  (.Q(\ram[90][2] ), 
	.D(n2024), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][1]  (.Q(\ram[90][1] ), 
	.D(n2023), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][0]  (.Q(\ram[90][0] ), 
	.D(n2022), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[86][15]  (.Q(\ram[86][15] ), 
	.D(n1973), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][14]  (.Q(\ram[86][14] ), 
	.D(n1972), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][13]  (.Q(\ram[86][13] ), 
	.D(n1971), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][12]  (.Q(\ram[86][12] ), 
	.D(n1970), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[86][11]  (.Q(\ram[86][11] ), 
	.D(n1969), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][10]  (.Q(\ram[86][10] ), 
	.D(n1968), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[86][9]  (.Q(\ram[86][9] ), 
	.D(n1967), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][8]  (.Q(\ram[86][8] ), 
	.D(n1966), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][7]  (.Q(\ram[86][7] ), 
	.D(n1965), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][6]  (.Q(\ram[86][6] ), 
	.D(n1964), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][5]  (.Q(\ram[86][5] ), 
	.D(n1963), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][4]  (.Q(\ram[86][4] ), 
	.D(n1962), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][3]  (.Q(\ram[86][3] ), 
	.D(n1961), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][2]  (.Q(\ram[86][2] ), 
	.D(n1960), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][1]  (.Q(\ram[86][1] ), 
	.D(n1959), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[86][0]  (.Q(\ram[86][0] ), 
	.D(n1958), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[82][15]  (.Q(\ram[82][15] ), 
	.D(n1909), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][14]  (.Q(\ram[82][14] ), 
	.D(n1908), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][13]  (.Q(\ram[82][13] ), 
	.D(n1907), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][12]  (.Q(\ram[82][12] ), 
	.D(n1906), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][11]  (.Q(\ram[82][11] ), 
	.D(n1905), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[82][10]  (.Q(\ram[82][10] ), 
	.D(n1904), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[82][9]  (.Q(\ram[82][9] ), 
	.D(n1903), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[82][8]  (.Q(\ram[82][8] ), 
	.D(n1902), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][7]  (.Q(\ram[82][7] ), 
	.D(n1901), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[82][6]  (.Q(\ram[82][6] ), 
	.D(n1900), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][5]  (.Q(\ram[82][5] ), 
	.D(n1899), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][4]  (.Q(\ram[82][4] ), 
	.D(n1898), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][3]  (.Q(\ram[82][3] ), 
	.D(n1897), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[82][2]  (.Q(\ram[82][2] ), 
	.D(n1896), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][1]  (.Q(\ram[82][1] ), 
	.D(n1895), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[82][0]  (.Q(\ram[82][0] ), 
	.D(n1894), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[78][15]  (.Q(\ram[78][15] ), 
	.D(n1845), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][14]  (.Q(\ram[78][14] ), 
	.D(n1844), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[78][13]  (.Q(\ram[78][13] ), 
	.D(n1843), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][12]  (.Q(\ram[78][12] ), 
	.D(n1842), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][11]  (.Q(\ram[78][11] ), 
	.D(n1841), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][10]  (.Q(\ram[78][10] ), 
	.D(n1840), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][9]  (.Q(\ram[78][9] ), 
	.D(n1839), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[78][8]  (.Q(\ram[78][8] ), 
	.D(n1838), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[78][7]  (.Q(\ram[78][7] ), 
	.D(n1837), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][6]  (.Q(\ram[78][6] ), 
	.D(n1836), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][5]  (.Q(\ram[78][5] ), 
	.D(n1835), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][4]  (.Q(\ram[78][4] ), 
	.D(n1834), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][3]  (.Q(\ram[78][3] ), 
	.D(n1833), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[78][2]  (.Q(\ram[78][2] ), 
	.D(n1832), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[78][1]  (.Q(\ram[78][1] ), 
	.D(n1831), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[78][0]  (.Q(\ram[78][0] ), 
	.D(n1830), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[74][15]  (.Q(\ram[74][15] ), 
	.D(n1781), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][14]  (.Q(\ram[74][14] ), 
	.D(n1780), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][13]  (.Q(\ram[74][13] ), 
	.D(n1779), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[74][12]  (.Q(\ram[74][12] ), 
	.D(n1778), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][11]  (.Q(\ram[74][11] ), 
	.D(n1777), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][10]  (.Q(\ram[74][10] ), 
	.D(n1776), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][9]  (.Q(\ram[74][9] ), 
	.D(n1775), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[74][8]  (.Q(\ram[74][8] ), 
	.D(n1774), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[74][7]  (.Q(\ram[74][7] ), 
	.D(n1773), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][6]  (.Q(\ram[74][6] ), 
	.D(n1772), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][5]  (.Q(\ram[74][5] ), 
	.D(n1771), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][4]  (.Q(\ram[74][4] ), 
	.D(n1770), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][3]  (.Q(\ram[74][3] ), 
	.D(n1769), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[74][2]  (.Q(\ram[74][2] ), 
	.D(n1768), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][1]  (.Q(\ram[74][1] ), 
	.D(n1767), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[74][0]  (.Q(\ram[74][0] ), 
	.D(n1766), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[70][15]  (.Q(\ram[70][15] ), 
	.D(n1717), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][14]  (.Q(\ram[70][14] ), 
	.D(n1716), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][13]  (.Q(\ram[70][13] ), 
	.D(n1715), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][12]  (.Q(\ram[70][12] ), 
	.D(n1714), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][11]  (.Q(\ram[70][11] ), 
	.D(n1713), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][10]  (.Q(\ram[70][10] ), 
	.D(n1712), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][9]  (.Q(\ram[70][9] ), 
	.D(n1711), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][8]  (.Q(\ram[70][8] ), 
	.D(n1710), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][7]  (.Q(\ram[70][7] ), 
	.D(n1709), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][6]  (.Q(\ram[70][6] ), 
	.D(n1708), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][5]  (.Q(\ram[70][5] ), 
	.D(n1707), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][4]  (.Q(\ram[70][4] ), 
	.D(n1706), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][3]  (.Q(\ram[70][3] ), 
	.D(n1705), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[70][2]  (.Q(\ram[70][2] ), 
	.D(n1704), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][1]  (.Q(\ram[70][1] ), 
	.D(n1703), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[70][0]  (.Q(\ram[70][0] ), 
	.D(n1702), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[66][15]  (.Q(\ram[66][15] ), 
	.D(n1653), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][14]  (.Q(\ram[66][14] ), 
	.D(n1652), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][13]  (.Q(\ram[66][13] ), 
	.D(n1651), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[66][12]  (.Q(\ram[66][12] ), 
	.D(n1650), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[66][11]  (.Q(\ram[66][11] ), 
	.D(n1649), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][10]  (.Q(\ram[66][10] ), 
	.D(n1648), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[66][9]  (.Q(\ram[66][9] ), 
	.D(n1647), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[66][8]  (.Q(\ram[66][8] ), 
	.D(n1646), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][7]  (.Q(\ram[66][7] ), 
	.D(n1645), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][6]  (.Q(\ram[66][6] ), 
	.D(n1644), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][5]  (.Q(\ram[66][5] ), 
	.D(n1643), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][4]  (.Q(\ram[66][4] ), 
	.D(n1642), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][3]  (.Q(\ram[66][3] ), 
	.D(n1641), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][2]  (.Q(\ram[66][2] ), 
	.D(n1640), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][1]  (.Q(\ram[66][1] ), 
	.D(n1639), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][0]  (.Q(\ram[66][0] ), 
	.D(n1638), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[62][15]  (.Q(\ram[62][15] ), 
	.D(n1589), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][14]  (.Q(\ram[62][14] ), 
	.D(n1588), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][13]  (.Q(\ram[62][13] ), 
	.D(n1587), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][12]  (.Q(\ram[62][12] ), 
	.D(n1586), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[62][11]  (.Q(\ram[62][11] ), 
	.D(n1585), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][10]  (.Q(\ram[62][10] ), 
	.D(n1584), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][9]  (.Q(\ram[62][9] ), 
	.D(n1583), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[62][8]  (.Q(\ram[62][8] ), 
	.D(n1582), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][7]  (.Q(\ram[62][7] ), 
	.D(n1581), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][6]  (.Q(\ram[62][6] ), 
	.D(n1580), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][5]  (.Q(\ram[62][5] ), 
	.D(n1579), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][4]  (.Q(\ram[62][4] ), 
	.D(n1578), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[62][3]  (.Q(\ram[62][3] ), 
	.D(n1577), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][2]  (.Q(\ram[62][2] ), 
	.D(n1576), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[62][1]  (.Q(\ram[62][1] ), 
	.D(n1575), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[62][0]  (.Q(\ram[62][0] ), 
	.D(n1574), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[58][15]  (.Q(\ram[58][15] ), 
	.D(n1525), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[58][14]  (.Q(\ram[58][14] ), 
	.D(n1524), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[58][13]  (.Q(\ram[58][13] ), 
	.D(n1523), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[58][12]  (.Q(\ram[58][12] ), 
	.D(n1522), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][11]  (.Q(\ram[58][11] ), 
	.D(n1521), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][10]  (.Q(\ram[58][10] ), 
	.D(n1520), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[58][9]  (.Q(\ram[58][9] ), 
	.D(n1519), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][8]  (.Q(\ram[58][8] ), 
	.D(n1518), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[58][7]  (.Q(\ram[58][7] ), 
	.D(n1517), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][6]  (.Q(\ram[58][6] ), 
	.D(n1516), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][5]  (.Q(\ram[58][5] ), 
	.D(n1515), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[58][4]  (.Q(\ram[58][4] ), 
	.D(n1514), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][3]  (.Q(\ram[58][3] ), 
	.D(n1513), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][2]  (.Q(\ram[58][2] ), 
	.D(n1512), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][1]  (.Q(\ram[58][1] ), 
	.D(n1511), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][0]  (.Q(\ram[58][0] ), 
	.D(n1510), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[54][15]  (.Q(\ram[54][15] ), 
	.D(n1461), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][14]  (.Q(\ram[54][14] ), 
	.D(n1460), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[54][13]  (.Q(\ram[54][13] ), 
	.D(n1459), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[54][12]  (.Q(\ram[54][12] ), 
	.D(n1458), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][11]  (.Q(\ram[54][11] ), 
	.D(n1457), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][10]  (.Q(\ram[54][10] ), 
	.D(n1456), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][9]  (.Q(\ram[54][9] ), 
	.D(n1455), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][8]  (.Q(\ram[54][8] ), 
	.D(n1454), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][7]  (.Q(\ram[54][7] ), 
	.D(n1453), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][6]  (.Q(\ram[54][6] ), 
	.D(n1452), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][5]  (.Q(\ram[54][5] ), 
	.D(n1451), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][4]  (.Q(\ram[54][4] ), 
	.D(n1450), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][3]  (.Q(\ram[54][3] ), 
	.D(n1449), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][2]  (.Q(\ram[54][2] ), 
	.D(n1448), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][1]  (.Q(\ram[54][1] ), 
	.D(n1447), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][0]  (.Q(\ram[54][0] ), 
	.D(n1446), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[50][15]  (.Q(\ram[50][15] ), 
	.D(n1397), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[50][14]  (.Q(\ram[50][14] ), 
	.D(n1396), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[50][13]  (.Q(\ram[50][13] ), 
	.D(n1395), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[50][12]  (.Q(\ram[50][12] ), 
	.D(n1394), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][11]  (.Q(\ram[50][11] ), 
	.D(n1393), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][10]  (.Q(\ram[50][10] ), 
	.D(n1392), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][9]  (.Q(\ram[50][9] ), 
	.D(n1391), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[50][8]  (.Q(\ram[50][8] ), 
	.D(n1390), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[50][7]  (.Q(\ram[50][7] ), 
	.D(n1389), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[50][6]  (.Q(\ram[50][6] ), 
	.D(n1388), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[50][5]  (.Q(\ram[50][5] ), 
	.D(n1387), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][4]  (.Q(\ram[50][4] ), 
	.D(n1386), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][3]  (.Q(\ram[50][3] ), 
	.D(n1385), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[50][2]  (.Q(\ram[50][2] ), 
	.D(n1384), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[50][1]  (.Q(\ram[50][1] ), 
	.D(n1383), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[50][0]  (.Q(\ram[50][0] ), 
	.D(n1382), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[46][15]  (.Q(\ram[46][15] ), 
	.D(n1333), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[46][14]  (.Q(\ram[46][14] ), 
	.D(n1332), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][13]  (.Q(\ram[46][13] ), 
	.D(n1331), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[46][12]  (.Q(\ram[46][12] ), 
	.D(n1330), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[46][11]  (.Q(\ram[46][11] ), 
	.D(n1329), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][10]  (.Q(\ram[46][10] ), 
	.D(n1328), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[46][9]  (.Q(\ram[46][9] ), 
	.D(n1327), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[46][8]  (.Q(\ram[46][8] ), 
	.D(n1326), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[46][7]  (.Q(\ram[46][7] ), 
	.D(n1325), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[46][6]  (.Q(\ram[46][6] ), 
	.D(n1324), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][5]  (.Q(\ram[46][5] ), 
	.D(n1323), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][4]  (.Q(\ram[46][4] ), 
	.D(n1322), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][3]  (.Q(\ram[46][3] ), 
	.D(n1321), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][2]  (.Q(\ram[46][2] ), 
	.D(n1320), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][1]  (.Q(\ram[46][1] ), 
	.D(n1319), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][0]  (.Q(\ram[46][0] ), 
	.D(n1318), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[42][15]  (.Q(\ram[42][15] ), 
	.D(n1269), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[42][14]  (.Q(\ram[42][14] ), 
	.D(n1268), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][13]  (.Q(\ram[42][13] ), 
	.D(n1267), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][12]  (.Q(\ram[42][12] ), 
	.D(n1266), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[42][11]  (.Q(\ram[42][11] ), 
	.D(n1265), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][10]  (.Q(\ram[42][10] ), 
	.D(n1264), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[42][9]  (.Q(\ram[42][9] ), 
	.D(n1263), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[42][8]  (.Q(\ram[42][8] ), 
	.D(n1262), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][7]  (.Q(\ram[42][7] ), 
	.D(n1261), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[42][6]  (.Q(\ram[42][6] ), 
	.D(n1260), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][5]  (.Q(\ram[42][5] ), 
	.D(n1259), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][4]  (.Q(\ram[42][4] ), 
	.D(n1258), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][3]  (.Q(\ram[42][3] ), 
	.D(n1257), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][2]  (.Q(\ram[42][2] ), 
	.D(n1256), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][1]  (.Q(\ram[42][1] ), 
	.D(n1255), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[42][0]  (.Q(\ram[42][0] ), 
	.D(n1254), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[38][15]  (.Q(\ram[38][15] ), 
	.D(n1205), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][14]  (.Q(\ram[38][14] ), 
	.D(n1204), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][13]  (.Q(\ram[38][13] ), 
	.D(n1203), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][12]  (.Q(\ram[38][12] ), 
	.D(n1202), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[38][11]  (.Q(\ram[38][11] ), 
	.D(n1201), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[38][10]  (.Q(\ram[38][10] ), 
	.D(n1200), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[38][9]  (.Q(\ram[38][9] ), 
	.D(n1199), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][8]  (.Q(\ram[38][8] ), 
	.D(n1198), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][7]  (.Q(\ram[38][7] ), 
	.D(n1197), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[38][6]  (.Q(\ram[38][6] ), 
	.D(n1196), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[38][5]  (.Q(\ram[38][5] ), 
	.D(n1195), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[38][4]  (.Q(\ram[38][4] ), 
	.D(n1194), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[38][3]  (.Q(\ram[38][3] ), 
	.D(n1193), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[38][2]  (.Q(\ram[38][2] ), 
	.D(n1192), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[38][1]  (.Q(\ram[38][1] ), 
	.D(n1191), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[38][0]  (.Q(\ram[38][0] ), 
	.D(n1190), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[34][15]  (.Q(\ram[34][15] ), 
	.D(n1141), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][14]  (.Q(\ram[34][14] ), 
	.D(n1140), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][13]  (.Q(\ram[34][13] ), 
	.D(n1139), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][12]  (.Q(\ram[34][12] ), 
	.D(n1138), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[34][11]  (.Q(\ram[34][11] ), 
	.D(n1137), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][10]  (.Q(\ram[34][10] ), 
	.D(n1136), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[34][9]  (.Q(\ram[34][9] ), 
	.D(n1135), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][8]  (.Q(\ram[34][8] ), 
	.D(n1134), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[34][7]  (.Q(\ram[34][7] ), 
	.D(n1133), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][6]  (.Q(\ram[34][6] ), 
	.D(n1132), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][5]  (.Q(\ram[34][5] ), 
	.D(n1131), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][4]  (.Q(\ram[34][4] ), 
	.D(n1130), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[34][3]  (.Q(\ram[34][3] ), 
	.D(n1129), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][2]  (.Q(\ram[34][2] ), 
	.D(n1128), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[34][1]  (.Q(\ram[34][1] ), 
	.D(n1127), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[34][0]  (.Q(\ram[34][0] ), 
	.D(n1126), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[30][15]  (.Q(\ram[30][15] ), 
	.D(n1077), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[30][14]  (.Q(\ram[30][14] ), 
	.D(n1076), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][13]  (.Q(\ram[30][13] ), 
	.D(n1075), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[30][12]  (.Q(\ram[30][12] ), 
	.D(n1074), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[30][11]  (.Q(\ram[30][11] ), 
	.D(n1073), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][10]  (.Q(\ram[30][10] ), 
	.D(n1072), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[30][9]  (.Q(\ram[30][9] ), 
	.D(n1071), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][8]  (.Q(\ram[30][8] ), 
	.D(n1070), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][7]  (.Q(\ram[30][7] ), 
	.D(n1069), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][6]  (.Q(\ram[30][6] ), 
	.D(n1068), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][5]  (.Q(\ram[30][5] ), 
	.D(n1067), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][4]  (.Q(\ram[30][4] ), 
	.D(n1066), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[30][3]  (.Q(\ram[30][3] ), 
	.D(n1065), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][2]  (.Q(\ram[30][2] ), 
	.D(n1064), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[30][1]  (.Q(\ram[30][1] ), 
	.D(n1063), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][0]  (.Q(\ram[30][0] ), 
	.D(n1062), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[26][15]  (.Q(\ram[26][15] ), 
	.D(n1013), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][14]  (.Q(\ram[26][14] ), 
	.D(n1012), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][13]  (.Q(\ram[26][13] ), 
	.D(n1011), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][12]  (.Q(\ram[26][12] ), 
	.D(n1010), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][11]  (.Q(\ram[26][11] ), 
	.D(n1009), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][10]  (.Q(\ram[26][10] ), 
	.D(n1008), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][9]  (.Q(\ram[26][9] ), 
	.D(n1007), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][8]  (.Q(\ram[26][8] ), 
	.D(n1006), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][7]  (.Q(\ram[26][7] ), 
	.D(n1005), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][6]  (.Q(\ram[26][6] ), 
	.D(n1004), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][5]  (.Q(\ram[26][5] ), 
	.D(n1003), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][4]  (.Q(\ram[26][4] ), 
	.D(n1002), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][3]  (.Q(\ram[26][3] ), 
	.D(n1001), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][2]  (.Q(\ram[26][2] ), 
	.D(n1000), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[26][1]  (.Q(\ram[26][1] ), 
	.D(n999), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][0]  (.Q(\ram[26][0] ), 
	.D(n998), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[22][15]  (.Q(\ram[22][15] ), 
	.D(n949), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][14]  (.Q(\ram[22][14] ), 
	.D(n948), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][13]  (.Q(\ram[22][13] ), 
	.D(n947), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[22][12]  (.Q(\ram[22][12] ), 
	.D(n946), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[22][11]  (.Q(\ram[22][11] ), 
	.D(n945), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][10]  (.Q(\ram[22][10] ), 
	.D(n944), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[22][9]  (.Q(\ram[22][9] ), 
	.D(n943), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][8]  (.Q(\ram[22][8] ), 
	.D(n942), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][7]  (.Q(\ram[22][7] ), 
	.D(n941), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][6]  (.Q(\ram[22][6] ), 
	.D(n940), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[22][5]  (.Q(\ram[22][5] ), 
	.D(n939), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[22][4]  (.Q(\ram[22][4] ), 
	.D(n938), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][3]  (.Q(\ram[22][3] ), 
	.D(n937), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[22][2]  (.Q(\ram[22][2] ), 
	.D(n936), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[22][1]  (.Q(\ram[22][1] ), 
	.D(n935), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][0]  (.Q(\ram[22][0] ), 
	.D(n934), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[18][15]  (.Q(\ram[18][15] ), 
	.D(n885), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[18][14]  (.Q(\ram[18][14] ), 
	.D(n884), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][13]  (.Q(\ram[18][13] ), 
	.D(n883), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[18][12]  (.Q(\ram[18][12] ), 
	.D(n882), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][11]  (.Q(\ram[18][11] ), 
	.D(n881), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[18][10]  (.Q(\ram[18][10] ), 
	.D(n880), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][9]  (.Q(\ram[18][9] ), 
	.D(n879), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[18][8]  (.Q(\ram[18][8] ), 
	.D(n878), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][7]  (.Q(\ram[18][7] ), 
	.D(n877), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[18][6]  (.Q(\ram[18][6] ), 
	.D(n876), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][5]  (.Q(\ram[18][5] ), 
	.D(n875), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][4]  (.Q(\ram[18][4] ), 
	.D(n874), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][3]  (.Q(\ram[18][3] ), 
	.D(n873), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[18][2]  (.Q(\ram[18][2] ), 
	.D(n872), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][1]  (.Q(\ram[18][1] ), 
	.D(n871), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[18][0]  (.Q(\ram[18][0] ), 
	.D(n870), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[14][15]  (.Q(\ram[14][15] ), 
	.D(n821), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][14]  (.Q(\ram[14][14] ), 
	.D(n820), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][13]  (.Q(\ram[14][13] ), 
	.D(n819), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][12]  (.Q(\ram[14][12] ), 
	.D(n818), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[14][11]  (.Q(\ram[14][11] ), 
	.D(n817), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[14][10]  (.Q(\ram[14][10] ), 
	.D(n816), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[14][9]  (.Q(\ram[14][9] ), 
	.D(n815), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[14][8]  (.Q(\ram[14][8] ), 
	.D(n814), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][7]  (.Q(\ram[14][7] ), 
	.D(n813), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][6]  (.Q(\ram[14][6] ), 
	.D(n812), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][5]  (.Q(\ram[14][5] ), 
	.D(n811), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[14][4]  (.Q(\ram[14][4] ), 
	.D(n810), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][3]  (.Q(\ram[14][3] ), 
	.D(n809), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][2]  (.Q(\ram[14][2] ), 
	.D(n808), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][1]  (.Q(\ram[14][1] ), 
	.D(n807), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[14][0]  (.Q(\ram[14][0] ), 
	.D(n806), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[10][15]  (.Q(\ram[10][15] ), 
	.D(n757), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][14]  (.Q(\ram[10][14] ), 
	.D(n756), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[10][13]  (.Q(\ram[10][13] ), 
	.D(n755), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[10][12]  (.Q(\ram[10][12] ), 
	.D(n754), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[10][11]  (.Q(\ram[10][11] ), 
	.D(n753), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[10][10]  (.Q(\ram[10][10] ), 
	.D(n752), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][9]  (.Q(\ram[10][9] ), 
	.D(n751), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[10][8]  (.Q(\ram[10][8] ), 
	.D(n750), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][7]  (.Q(\ram[10][7] ), 
	.D(n749), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][6]  (.Q(\ram[10][6] ), 
	.D(n748), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][5]  (.Q(\ram[10][5] ), 
	.D(n747), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[10][4]  (.Q(\ram[10][4] ), 
	.D(n746), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[10][3]  (.Q(\ram[10][3] ), 
	.D(n745), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][2]  (.Q(\ram[10][2] ), 
	.D(n744), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[10][1]  (.Q(\ram[10][1] ), 
	.D(n743), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[10][0]  (.Q(\ram[10][0] ), 
	.D(n742), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[6][15]  (.Q(\ram[6][15] ), 
	.D(n693), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][14]  (.Q(\ram[6][14] ), 
	.D(n692), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][13]  (.Q(\ram[6][13] ), 
	.D(n691), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[6][12]  (.Q(\ram[6][12] ), 
	.D(n690), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[6][11]  (.Q(\ram[6][11] ), 
	.D(n689), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[6][10]  (.Q(\ram[6][10] ), 
	.D(n688), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][9]  (.Q(\ram[6][9] ), 
	.D(n687), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[6][8]  (.Q(\ram[6][8] ), 
	.D(n686), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][7]  (.Q(\ram[6][7] ), 
	.D(n685), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][6]  (.Q(\ram[6][6] ), 
	.D(n684), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][5]  (.Q(\ram[6][5] ), 
	.D(n683), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[6][4]  (.Q(\ram[6][4] ), 
	.D(n682), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][3]  (.Q(\ram[6][3] ), 
	.D(n681), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[6][2]  (.Q(\ram[6][2] ), 
	.D(n680), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][1]  (.Q(\ram[6][1] ), 
	.D(n679), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[6][0]  (.Q(\ram[6][0] ), 
	.D(n678), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[2][15]  (.Q(\ram[2][15] ), 
	.D(n629), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[2][14]  (.Q(\ram[2][14] ), 
	.D(n628), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][13]  (.Q(\ram[2][13] ), 
	.D(n627), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[2][12]  (.Q(\ram[2][12] ), 
	.D(n626), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][11]  (.Q(\ram[2][11] ), 
	.D(n625), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[2][10]  (.Q(\ram[2][10] ), 
	.D(n624), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[2][9]  (.Q(\ram[2][9] ), 
	.D(n623), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[2][8]  (.Q(\ram[2][8] ), 
	.D(n622), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[2][7]  (.Q(\ram[2][7] ), 
	.D(n621), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[2][6]  (.Q(\ram[2][6] ), 
	.D(n620), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[2][5]  (.Q(\ram[2][5] ), 
	.D(n619), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[2][4]  (.Q(\ram[2][4] ), 
	.D(n618), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][3]  (.Q(\ram[2][3] ), 
	.D(n617), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[2][2]  (.Q(\ram[2][2] ), 
	.D(n616), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][1]  (.Q(\ram[2][1] ), 
	.D(n615), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][0]  (.Q(\ram[2][0] ), 
	.D(n614), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[252][15]  (.Q(\ram[252][15] ), 
	.D(n4629), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[252][14]  (.Q(\ram[252][14] ), 
	.D(n4628), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[252][13]  (.Q(\ram[252][13] ), 
	.D(n4627), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][12]  (.Q(\ram[252][12] ), 
	.D(n4626), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[252][11]  (.Q(\ram[252][11] ), 
	.D(n4625), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[252][10]  (.Q(\ram[252][10] ), 
	.D(n4624), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][9]  (.Q(\ram[252][9] ), 
	.D(n4623), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][8]  (.Q(\ram[252][8] ), 
	.D(n4622), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][7]  (.Q(\ram[252][7] ), 
	.D(n4621), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[252][6]  (.Q(\ram[252][6] ), 
	.D(n4620), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[252][5]  (.Q(\ram[252][5] ), 
	.D(n4619), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[252][4]  (.Q(\ram[252][4] ), 
	.D(n4618), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[252][3]  (.Q(\ram[252][3] ), 
	.D(n4617), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[252][2]  (.Q(\ram[252][2] ), 
	.D(n4616), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[252][1]  (.Q(\ram[252][1] ), 
	.D(n4615), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[252][0]  (.Q(\ram[252][0] ), 
	.D(n4614), 
	.CK(clk));
   QDFFEHD \ram_reg[248][15]  (.Q(\ram[248][15] ), 
	.D(n4565), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][14]  (.Q(\ram[248][14] ), 
	.D(n4564), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][13]  (.Q(\ram[248][13] ), 
	.D(n4563), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][12]  (.Q(\ram[248][12] ), 
	.D(n4562), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[248][11]  (.Q(\ram[248][11] ), 
	.D(n4561), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][10]  (.Q(\ram[248][10] ), 
	.D(n4560), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][9]  (.Q(\ram[248][9] ), 
	.D(n4559), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][8]  (.Q(\ram[248][8] ), 
	.D(n4558), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][7]  (.Q(\ram[248][7] ), 
	.D(n4557), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][6]  (.Q(\ram[248][6] ), 
	.D(n4556), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][5]  (.Q(\ram[248][5] ), 
	.D(n4555), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[248][4]  (.Q(\ram[248][4] ), 
	.D(n4554), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[248][3]  (.Q(\ram[248][3] ), 
	.D(n4553), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[248][2]  (.Q(\ram[248][2] ), 
	.D(n4552), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][1]  (.Q(\ram[248][1] ), 
	.D(n4551), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[248][0]  (.Q(\ram[248][0] ), 
	.D(n4550), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][15]  (.Q(\ram[244][15] ), 
	.D(n4501), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][14]  (.Q(\ram[244][14] ), 
	.D(n4500), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[244][13]  (.Q(\ram[244][13] ), 
	.D(n4499), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][12]  (.Q(\ram[244][12] ), 
	.D(n4498), 
	.CK(clk));
   QDFFEHD \ram_reg[244][11]  (.Q(\ram[244][11] ), 
	.D(n4497), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][10]  (.Q(\ram[244][10] ), 
	.D(n4496), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][9]  (.Q(\ram[244][9] ), 
	.D(n4495), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[244][8]  (.Q(\ram[244][8] ), 
	.D(n4494), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[244][7]  (.Q(\ram[244][7] ), 
	.D(n4493), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[244][6]  (.Q(\ram[244][6] ), 
	.D(n4492), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][5]  (.Q(\ram[244][5] ), 
	.D(n4491), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][4]  (.Q(\ram[244][4] ), 
	.D(n4490), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][3]  (.Q(\ram[244][3] ), 
	.D(n4489), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[244][2]  (.Q(\ram[244][2] ), 
	.D(n4488), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][1]  (.Q(\ram[244][1] ), 
	.D(n4487), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][0]  (.Q(\ram[244][0] ), 
	.D(n4486), 
	.CK(clk));
   QDFFEHD \ram_reg[240][15]  (.Q(\ram[240][15] ), 
	.D(n4437), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[240][14]  (.Q(\ram[240][14] ), 
	.D(n4436), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][13]  (.Q(\ram[240][13] ), 
	.D(n4435), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][12]  (.Q(\ram[240][12] ), 
	.D(n4434), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[240][11]  (.Q(\ram[240][11] ), 
	.D(n4433), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[240][10]  (.Q(\ram[240][10] ), 
	.D(n4432), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][9]  (.Q(\ram[240][9] ), 
	.D(n4431), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[240][8]  (.Q(\ram[240][8] ), 
	.D(n4430), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][7]  (.Q(\ram[240][7] ), 
	.D(n4429), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[240][6]  (.Q(\ram[240][6] ), 
	.D(n4428), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][5]  (.Q(\ram[240][5] ), 
	.D(n4427), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][4]  (.Q(\ram[240][4] ), 
	.D(n4426), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][3]  (.Q(\ram[240][3] ), 
	.D(n4425), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][2]  (.Q(\ram[240][2] ), 
	.D(n4424), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][1]  (.Q(\ram[240][1] ), 
	.D(n4423), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][0]  (.Q(\ram[240][0] ), 
	.D(n4422), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[236][15]  (.Q(\ram[236][15] ), 
	.D(n4373), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][14]  (.Q(\ram[236][14] ), 
	.D(n4372), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[236][13]  (.Q(\ram[236][13] ), 
	.D(n4371), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][12]  (.Q(\ram[236][12] ), 
	.D(n4370), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[236][11]  (.Q(\ram[236][11] ), 
	.D(n4369), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[236][10]  (.Q(\ram[236][10] ), 
	.D(n4368), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[236][9]  (.Q(\ram[236][9] ), 
	.D(n4367), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[236][8]  (.Q(\ram[236][8] ), 
	.D(n4366), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[236][7]  (.Q(\ram[236][7] ), 
	.D(n4365), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[236][6]  (.Q(\ram[236][6] ), 
	.D(n4364), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[236][5]  (.Q(\ram[236][5] ), 
	.D(n4363), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][4]  (.Q(\ram[236][4] ), 
	.D(n4362), 
	.CK(clk_m__L3_N50));
   QDFFEHD \ram_reg[236][3]  (.Q(\ram[236][3] ), 
	.D(n4361), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[236][2]  (.Q(\ram[236][2] ), 
	.D(n4360), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][1]  (.Q(\ram[236][1] ), 
	.D(n4359), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[236][0]  (.Q(\ram[236][0] ), 
	.D(n4358), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[232][15]  (.Q(\ram[232][15] ), 
	.D(n4309), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[232][14]  (.Q(\ram[232][14] ), 
	.D(n4308), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[232][13]  (.Q(\ram[232][13] ), 
	.D(n4307), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[232][12]  (.Q(\ram[232][12] ), 
	.D(n4306), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][11]  (.Q(\ram[232][11] ), 
	.D(n4305), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[232][10]  (.Q(\ram[232][10] ), 
	.D(n4304), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][9]  (.Q(\ram[232][9] ), 
	.D(n4303), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][8]  (.Q(\ram[232][8] ), 
	.D(n4302), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][7]  (.Q(\ram[232][7] ), 
	.D(n4301), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][6]  (.Q(\ram[232][6] ), 
	.D(n4300), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][5]  (.Q(\ram[232][5] ), 
	.D(n4299), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[232][4]  (.Q(\ram[232][4] ), 
	.D(n4298), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[232][3]  (.Q(\ram[232][3] ), 
	.D(n4297), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[232][2]  (.Q(\ram[232][2] ), 
	.D(n4296), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[232][1]  (.Q(\ram[232][1] ), 
	.D(n4295), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[232][0]  (.Q(\ram[232][0] ), 
	.D(n4294), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[228][15]  (.Q(\ram[228][15] ), 
	.D(n4245), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[228][14]  (.Q(\ram[228][14] ), 
	.D(n4244), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[228][13]  (.Q(\ram[228][13] ), 
	.D(n4243), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[228][12]  (.Q(\ram[228][12] ), 
	.D(n4242), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[228][11]  (.Q(\ram[228][11] ), 
	.D(n4241), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][10]  (.Q(\ram[228][10] ), 
	.D(n4240), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][9]  (.Q(\ram[228][9] ), 
	.D(n4239), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][8]  (.Q(\ram[228][8] ), 
	.D(n4238), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][7]  (.Q(\ram[228][7] ), 
	.D(n4237), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[228][6]  (.Q(\ram[228][6] ), 
	.D(n4236), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[228][5]  (.Q(\ram[228][5] ), 
	.D(n4235), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[228][4]  (.Q(\ram[228][4] ), 
	.D(n4234), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[228][3]  (.Q(\ram[228][3] ), 
	.D(n4233), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[228][2]  (.Q(\ram[228][2] ), 
	.D(n4232), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[228][1]  (.Q(\ram[228][1] ), 
	.D(n4231), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[228][0]  (.Q(\ram[228][0] ), 
	.D(n4230), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][15]  (.Q(\ram[224][15] ), 
	.D(n4181), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][14]  (.Q(\ram[224][14] ), 
	.D(n4180), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][13]  (.Q(\ram[224][13] ), 
	.D(n4179), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][12]  (.Q(\ram[224][12] ), 
	.D(n4178), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][11]  (.Q(\ram[224][11] ), 
	.D(n4177), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][10]  (.Q(\ram[224][10] ), 
	.D(n4176), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[224][9]  (.Q(\ram[224][9] ), 
	.D(n4175), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][8]  (.Q(\ram[224][8] ), 
	.D(n4174), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][7]  (.Q(\ram[224][7] ), 
	.D(n4173), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[224][6]  (.Q(\ram[224][6] ), 
	.D(n4172), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[224][5]  (.Q(\ram[224][5] ), 
	.D(n4171), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][4]  (.Q(\ram[224][4] ), 
	.D(n4170), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][3]  (.Q(\ram[224][3] ), 
	.D(n4169), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[224][2]  (.Q(\ram[224][2] ), 
	.D(n4168), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][1]  (.Q(\ram[224][1] ), 
	.D(n4167), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[224][0]  (.Q(\ram[224][0] ), 
	.D(n4166), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[220][15]  (.Q(\ram[220][15] ), 
	.D(n4117), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][14]  (.Q(\ram[220][14] ), 
	.D(n4116), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][13]  (.Q(\ram[220][13] ), 
	.D(n4115), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][12]  (.Q(\ram[220][12] ), 
	.D(n4114), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][11]  (.Q(\ram[220][11] ), 
	.D(n4113), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][10]  (.Q(\ram[220][10] ), 
	.D(n4112), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][9]  (.Q(\ram[220][9] ), 
	.D(n4111), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][8]  (.Q(\ram[220][8] ), 
	.D(n4110), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][7]  (.Q(\ram[220][7] ), 
	.D(n4109), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][6]  (.Q(\ram[220][6] ), 
	.D(n4108), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[220][5]  (.Q(\ram[220][5] ), 
	.D(n4107), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[220][4]  (.Q(\ram[220][4] ), 
	.D(n4106), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][3]  (.Q(\ram[220][3] ), 
	.D(n4105), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[220][2]  (.Q(\ram[220][2] ), 
	.D(n4104), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][1]  (.Q(\ram[220][1] ), 
	.D(n4103), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][0]  (.Q(\ram[220][0] ), 
	.D(n4102), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[216][15]  (.Q(\ram[216][15] ), 
	.D(n4053), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][14]  (.Q(\ram[216][14] ), 
	.D(n4052), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][13]  (.Q(\ram[216][13] ), 
	.D(n4051), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][12]  (.Q(\ram[216][12] ), 
	.D(n4050), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][11]  (.Q(\ram[216][11] ), 
	.D(n4049), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[216][10]  (.Q(\ram[216][10] ), 
	.D(n4048), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][9]  (.Q(\ram[216][9] ), 
	.D(n4047), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[216][8]  (.Q(\ram[216][8] ), 
	.D(n4046), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][7]  (.Q(\ram[216][7] ), 
	.D(n4045), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][6]  (.Q(\ram[216][6] ), 
	.D(n4044), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][5]  (.Q(\ram[216][5] ), 
	.D(n4043), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[216][4]  (.Q(\ram[216][4] ), 
	.D(n4042), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[216][3]  (.Q(\ram[216][3] ), 
	.D(n4041), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][2]  (.Q(\ram[216][2] ), 
	.D(n4040), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][1]  (.Q(\ram[216][1] ), 
	.D(n4039), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][0]  (.Q(\ram[216][0] ), 
	.D(n4038), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[212][15]  (.Q(\ram[212][15] ), 
	.D(n3989), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[212][14]  (.Q(\ram[212][14] ), 
	.D(n3988), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][13]  (.Q(\ram[212][13] ), 
	.D(n3987), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][12]  (.Q(\ram[212][12] ), 
	.D(n3986), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][11]  (.Q(\ram[212][11] ), 
	.D(n3985), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][10]  (.Q(\ram[212][10] ), 
	.D(n3984), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][9]  (.Q(\ram[212][9] ), 
	.D(n3983), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][8]  (.Q(\ram[212][8] ), 
	.D(n3982), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][7]  (.Q(\ram[212][7] ), 
	.D(n3981), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][6]  (.Q(\ram[212][6] ), 
	.D(n3980), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][5]  (.Q(\ram[212][5] ), 
	.D(n3979), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][4]  (.Q(\ram[212][4] ), 
	.D(n3978), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[212][3]  (.Q(\ram[212][3] ), 
	.D(n3977), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][2]  (.Q(\ram[212][2] ), 
	.D(n3976), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][1]  (.Q(\ram[212][1] ), 
	.D(n3975), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][0]  (.Q(\ram[212][0] ), 
	.D(n3974), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[208][15]  (.Q(\ram[208][15] ), 
	.D(n3925), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[208][14]  (.Q(\ram[208][14] ), 
	.D(n3924), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[208][13]  (.Q(\ram[208][13] ), 
	.D(n3923), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][12]  (.Q(\ram[208][12] ), 
	.D(n3922), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][11]  (.Q(\ram[208][11] ), 
	.D(n3921), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[208][10]  (.Q(\ram[208][10] ), 
	.D(n3920), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[208][9]  (.Q(\ram[208][9] ), 
	.D(n3919), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][8]  (.Q(\ram[208][8] ), 
	.D(n3918), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][7]  (.Q(\ram[208][7] ), 
	.D(n3917), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[208][6]  (.Q(\ram[208][6] ), 
	.D(n3916), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][5]  (.Q(\ram[208][5] ), 
	.D(n3915), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][4]  (.Q(\ram[208][4] ), 
	.D(n3914), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[208][3]  (.Q(\ram[208][3] ), 
	.D(n3913), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[208][2]  (.Q(\ram[208][2] ), 
	.D(n3912), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[208][1]  (.Q(\ram[208][1] ), 
	.D(n3911), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[208][0]  (.Q(\ram[208][0] ), 
	.D(n3910), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[204][15]  (.Q(\ram[204][15] ), 
	.D(n3861), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][14]  (.Q(\ram[204][14] ), 
	.D(n3860), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][13]  (.Q(\ram[204][13] ), 
	.D(n3859), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[204][12]  (.Q(\ram[204][12] ), 
	.D(n3858), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][11]  (.Q(\ram[204][11] ), 
	.D(n3857), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][10]  (.Q(\ram[204][10] ), 
	.D(n3856), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][9]  (.Q(\ram[204][9] ), 
	.D(n3855), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][8]  (.Q(\ram[204][8] ), 
	.D(n3854), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][7]  (.Q(\ram[204][7] ), 
	.D(n3853), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][6]  (.Q(\ram[204][6] ), 
	.D(n3852), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[204][5]  (.Q(\ram[204][5] ), 
	.D(n3851), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][4]  (.Q(\ram[204][4] ), 
	.D(n3850), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][3]  (.Q(\ram[204][3] ), 
	.D(n3849), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][2]  (.Q(\ram[204][2] ), 
	.D(n3848), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][1]  (.Q(\ram[204][1] ), 
	.D(n3847), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][0]  (.Q(\ram[204][0] ), 
	.D(n3846), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[200][15]  (.Q(\ram[200][15] ), 
	.D(n3797), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[200][14]  (.Q(\ram[200][14] ), 
	.D(n3796), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][13]  (.Q(\ram[200][13] ), 
	.D(n3795), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][12]  (.Q(\ram[200][12] ), 
	.D(n3794), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[200][11]  (.Q(\ram[200][11] ), 
	.D(n3793), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][10]  (.Q(\ram[200][10] ), 
	.D(n3792), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[200][9]  (.Q(\ram[200][9] ), 
	.D(n3791), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][8]  (.Q(\ram[200][8] ), 
	.D(n3790), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][7]  (.Q(\ram[200][7] ), 
	.D(n3789), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][6]  (.Q(\ram[200][6] ), 
	.D(n3788), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][5]  (.Q(\ram[200][5] ), 
	.D(n3787), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][4]  (.Q(\ram[200][4] ), 
	.D(n3786), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][3]  (.Q(\ram[200][3] ), 
	.D(n3785), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][2]  (.Q(\ram[200][2] ), 
	.D(n3784), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][1]  (.Q(\ram[200][1] ), 
	.D(n3783), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][0]  (.Q(\ram[200][0] ), 
	.D(n3782), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[196][15]  (.Q(\ram[196][15] ), 
	.D(n3733), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[196][14]  (.Q(\ram[196][14] ), 
	.D(n3732), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][13]  (.Q(\ram[196][13] ), 
	.D(n3731), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[196][12]  (.Q(\ram[196][12] ), 
	.D(n3730), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[196][11]  (.Q(\ram[196][11] ), 
	.D(n3729), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][10]  (.Q(\ram[196][10] ), 
	.D(n3728), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][9]  (.Q(\ram[196][9] ), 
	.D(n3727), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[196][8]  (.Q(\ram[196][8] ), 
	.D(n3726), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][7]  (.Q(\ram[196][7] ), 
	.D(n3725), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][6]  (.Q(\ram[196][6] ), 
	.D(n3724), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][5]  (.Q(\ram[196][5] ), 
	.D(n3723), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][4]  (.Q(\ram[196][4] ), 
	.D(n3722), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][3]  (.Q(\ram[196][3] ), 
	.D(n3721), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[196][2]  (.Q(\ram[196][2] ), 
	.D(n3720), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][1]  (.Q(\ram[196][1] ), 
	.D(n3719), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][0]  (.Q(\ram[196][0] ), 
	.D(n3718), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[192][15]  (.Q(\ram[192][15] ), 
	.D(n3669), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][14]  (.Q(\ram[192][14] ), 
	.D(n3668), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][13]  (.Q(\ram[192][13] ), 
	.D(n3667), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][12]  (.Q(\ram[192][12] ), 
	.D(n3666), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][11]  (.Q(\ram[192][11] ), 
	.D(n3665), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][10]  (.Q(\ram[192][10] ), 
	.D(n3664), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][9]  (.Q(\ram[192][9] ), 
	.D(n3663), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][8]  (.Q(\ram[192][8] ), 
	.D(n3662), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][7]  (.Q(\ram[192][7] ), 
	.D(n3661), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][6]  (.Q(\ram[192][6] ), 
	.D(n3660), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][5]  (.Q(\ram[192][5] ), 
	.D(n3659), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][4]  (.Q(\ram[192][4] ), 
	.D(n3658), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][3]  (.Q(\ram[192][3] ), 
	.D(n3657), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[192][2]  (.Q(\ram[192][2] ), 
	.D(n3656), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][1]  (.Q(\ram[192][1] ), 
	.D(n3655), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][0]  (.Q(\ram[192][0] ), 
	.D(n3654), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[188][15]  (.Q(\ram[188][15] ), 
	.D(n3605), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][14]  (.Q(\ram[188][14] ), 
	.D(n3604), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][13]  (.Q(\ram[188][13] ), 
	.D(n3603), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][12]  (.Q(\ram[188][12] ), 
	.D(n3602), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][11]  (.Q(\ram[188][11] ), 
	.D(n3601), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[188][10]  (.Q(\ram[188][10] ), 
	.D(n3600), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][9]  (.Q(\ram[188][9] ), 
	.D(n3599), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[188][8]  (.Q(\ram[188][8] ), 
	.D(n3598), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][7]  (.Q(\ram[188][7] ), 
	.D(n3597), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][6]  (.Q(\ram[188][6] ), 
	.D(n3596), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][5]  (.Q(\ram[188][5] ), 
	.D(n3595), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][4]  (.Q(\ram[188][4] ), 
	.D(n3594), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][3]  (.Q(\ram[188][3] ), 
	.D(n3593), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[188][2]  (.Q(\ram[188][2] ), 
	.D(n3592), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][1]  (.Q(\ram[188][1] ), 
	.D(n3591), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][0]  (.Q(\ram[188][0] ), 
	.D(n3590), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][15]  (.Q(\ram[184][15] ), 
	.D(n3541), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][14]  (.Q(\ram[184][14] ), 
	.D(n3540), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][13]  (.Q(\ram[184][13] ), 
	.D(n3539), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[184][12]  (.Q(\ram[184][12] ), 
	.D(n3538), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[184][11]  (.Q(\ram[184][11] ), 
	.D(n3537), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][10]  (.Q(\ram[184][10] ), 
	.D(n3536), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][9]  (.Q(\ram[184][9] ), 
	.D(n3535), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][8]  (.Q(\ram[184][8] ), 
	.D(n3534), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][7]  (.Q(\ram[184][7] ), 
	.D(n3533), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[184][6]  (.Q(\ram[184][6] ), 
	.D(n3532), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[184][5]  (.Q(\ram[184][5] ), 
	.D(n3531), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[184][4]  (.Q(\ram[184][4] ), 
	.D(n3530), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][3]  (.Q(\ram[184][3] ), 
	.D(n3529), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[184][2]  (.Q(\ram[184][2] ), 
	.D(n3528), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][1]  (.Q(\ram[184][1] ), 
	.D(n3527), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][0]  (.Q(\ram[184][0] ), 
	.D(n3526), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[180][15]  (.Q(\ram[180][15] ), 
	.D(n3477), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[180][14]  (.Q(\ram[180][14] ), 
	.D(n3476), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[180][13]  (.Q(\ram[180][13] ), 
	.D(n3475), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[180][12]  (.Q(\ram[180][12] ), 
	.D(n3474), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][11]  (.Q(\ram[180][11] ), 
	.D(n3473), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[180][10]  (.Q(\ram[180][10] ), 
	.D(n3472), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][9]  (.Q(\ram[180][9] ), 
	.D(n3471), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][8]  (.Q(\ram[180][8] ), 
	.D(n3470), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][7]  (.Q(\ram[180][7] ), 
	.D(n3469), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][6]  (.Q(\ram[180][6] ), 
	.D(n3468), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][5]  (.Q(\ram[180][5] ), 
	.D(n3467), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][4]  (.Q(\ram[180][4] ), 
	.D(n3466), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][3]  (.Q(\ram[180][3] ), 
	.D(n3465), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[180][2]  (.Q(\ram[180][2] ), 
	.D(n3464), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[180][1]  (.Q(\ram[180][1] ), 
	.D(n3463), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][0]  (.Q(\ram[180][0] ), 
	.D(n3462), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[176][15]  (.Q(\ram[176][15] ), 
	.D(n3413), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[176][14]  (.Q(\ram[176][14] ), 
	.D(n3412), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][13]  (.Q(\ram[176][13] ), 
	.D(n3411), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[176][12]  (.Q(\ram[176][12] ), 
	.D(n3410), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[176][11]  (.Q(\ram[176][11] ), 
	.D(n3409), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[176][10]  (.Q(\ram[176][10] ), 
	.D(n3408), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[176][9]  (.Q(\ram[176][9] ), 
	.D(n3407), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][8]  (.Q(\ram[176][8] ), 
	.D(n3406), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[176][7]  (.Q(\ram[176][7] ), 
	.D(n3405), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][6]  (.Q(\ram[176][6] ), 
	.D(n3404), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][5]  (.Q(\ram[176][5] ), 
	.D(n3403), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][4]  (.Q(\ram[176][4] ), 
	.D(n3402), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][3]  (.Q(\ram[176][3] ), 
	.D(n3401), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][2]  (.Q(\ram[176][2] ), 
	.D(n3400), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][1]  (.Q(\ram[176][1] ), 
	.D(n3399), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][0]  (.Q(\ram[176][0] ), 
	.D(n3398), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[172][15]  (.Q(\ram[172][15] ), 
	.D(n3349), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[172][14]  (.Q(\ram[172][14] ), 
	.D(n3348), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][13]  (.Q(\ram[172][13] ), 
	.D(n3347), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[172][12]  (.Q(\ram[172][12] ), 
	.D(n3346), 
	.CK(clk));
   QDFFEHD \ram_reg[172][11]  (.Q(\ram[172][11] ), 
	.D(n3345), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[172][10]  (.Q(\ram[172][10] ), 
	.D(n3344), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[172][9]  (.Q(\ram[172][9] ), 
	.D(n3343), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][8]  (.Q(\ram[172][8] ), 
	.D(n3342), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[172][7]  (.Q(\ram[172][7] ), 
	.D(n3341), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[172][6]  (.Q(\ram[172][6] ), 
	.D(n3340), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][5]  (.Q(\ram[172][5] ), 
	.D(n3339), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[172][4]  (.Q(\ram[172][4] ), 
	.D(n3338), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[172][3]  (.Q(\ram[172][3] ), 
	.D(n3337), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][2]  (.Q(\ram[172][2] ), 
	.D(n3336), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[172][1]  (.Q(\ram[172][1] ), 
	.D(n3335), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[172][0]  (.Q(\ram[172][0] ), 
	.D(n3334), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][15]  (.Q(\ram[168][15] ), 
	.D(n3285), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][14]  (.Q(\ram[168][14] ), 
	.D(n3284), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][13]  (.Q(\ram[168][13] ), 
	.D(n3283), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][12]  (.Q(\ram[168][12] ), 
	.D(n3282), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][11]  (.Q(\ram[168][11] ), 
	.D(n3281), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[168][10]  (.Q(\ram[168][10] ), 
	.D(n3280), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[168][9]  (.Q(\ram[168][9] ), 
	.D(n3279), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][8]  (.Q(\ram[168][8] ), 
	.D(n3278), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[168][7]  (.Q(\ram[168][7] ), 
	.D(n3277), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[168][6]  (.Q(\ram[168][6] ), 
	.D(n3276), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][5]  (.Q(\ram[168][5] ), 
	.D(n3275), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][4]  (.Q(\ram[168][4] ), 
	.D(n3274), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][3]  (.Q(\ram[168][3] ), 
	.D(n3273), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[168][2]  (.Q(\ram[168][2] ), 
	.D(n3272), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[168][1]  (.Q(\ram[168][1] ), 
	.D(n3271), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[168][0]  (.Q(\ram[168][0] ), 
	.D(n3270), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[164][15]  (.Q(\ram[164][15] ), 
	.D(n3221), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[164][14]  (.Q(\ram[164][14] ), 
	.D(n3220), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][13]  (.Q(\ram[164][13] ), 
	.D(n3219), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[164][12]  (.Q(\ram[164][12] ), 
	.D(n3218), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][11]  (.Q(\ram[164][11] ), 
	.D(n3217), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[164][10]  (.Q(\ram[164][10] ), 
	.D(n3216), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[164][9]  (.Q(\ram[164][9] ), 
	.D(n3215), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][8]  (.Q(\ram[164][8] ), 
	.D(n3214), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][7]  (.Q(\ram[164][7] ), 
	.D(n3213), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[164][6]  (.Q(\ram[164][6] ), 
	.D(n3212), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][5]  (.Q(\ram[164][5] ), 
	.D(n3211), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][4]  (.Q(\ram[164][4] ), 
	.D(n3210), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[164][3]  (.Q(\ram[164][3] ), 
	.D(n3209), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][2]  (.Q(\ram[164][2] ), 
	.D(n3208), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][1]  (.Q(\ram[164][1] ), 
	.D(n3207), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][0]  (.Q(\ram[164][0] ), 
	.D(n3206), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][15]  (.Q(\ram[160][15] ), 
	.D(n3157), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][14]  (.Q(\ram[160][14] ), 
	.D(n3156), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][13]  (.Q(\ram[160][13] ), 
	.D(n3155), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][12]  (.Q(\ram[160][12] ), 
	.D(n3154), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][11]  (.Q(\ram[160][11] ), 
	.D(n3153), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][10]  (.Q(\ram[160][10] ), 
	.D(n3152), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][9]  (.Q(\ram[160][9] ), 
	.D(n3151), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][8]  (.Q(\ram[160][8] ), 
	.D(n3150), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[160][7]  (.Q(\ram[160][7] ), 
	.D(n3149), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][6]  (.Q(\ram[160][6] ), 
	.D(n3148), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][5]  (.Q(\ram[160][5] ), 
	.D(n3147), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[160][4]  (.Q(\ram[160][4] ), 
	.D(n3146), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[160][3]  (.Q(\ram[160][3] ), 
	.D(n3145), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][2]  (.Q(\ram[160][2] ), 
	.D(n3144), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][1]  (.Q(\ram[160][1] ), 
	.D(n3143), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][0]  (.Q(\ram[160][0] ), 
	.D(n3142), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[156][15]  (.Q(\ram[156][15] ), 
	.D(n3093), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][14]  (.Q(\ram[156][14] ), 
	.D(n3092), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][13]  (.Q(\ram[156][13] ), 
	.D(n3091), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][12]  (.Q(\ram[156][12] ), 
	.D(n3090), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][11]  (.Q(\ram[156][11] ), 
	.D(n3089), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][10]  (.Q(\ram[156][10] ), 
	.D(n3088), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[156][9]  (.Q(\ram[156][9] ), 
	.D(n3087), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[156][8]  (.Q(\ram[156][8] ), 
	.D(n3086), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[156][7]  (.Q(\ram[156][7] ), 
	.D(n3085), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[156][6]  (.Q(\ram[156][6] ), 
	.D(n3084), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[156][5]  (.Q(\ram[156][5] ), 
	.D(n3083), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[156][4]  (.Q(\ram[156][4] ), 
	.D(n3082), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[156][3]  (.Q(\ram[156][3] ), 
	.D(n3081), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[156][2]  (.Q(\ram[156][2] ), 
	.D(n3080), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[156][1]  (.Q(\ram[156][1] ), 
	.D(n3079), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[156][0]  (.Q(\ram[156][0] ), 
	.D(n3078), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[152][15]  (.Q(\ram[152][15] ), 
	.D(n3029), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[152][14]  (.Q(\ram[152][14] ), 
	.D(n3028), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[152][13]  (.Q(\ram[152][13] ), 
	.D(n3027), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[152][12]  (.Q(\ram[152][12] ), 
	.D(n3026), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[152][11]  (.Q(\ram[152][11] ), 
	.D(n3025), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[152][10]  (.Q(\ram[152][10] ), 
	.D(n3024), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[152][9]  (.Q(\ram[152][9] ), 
	.D(n3023), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[152][8]  (.Q(\ram[152][8] ), 
	.D(n3022), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[152][7]  (.Q(\ram[152][7] ), 
	.D(n3021), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][6]  (.Q(\ram[152][6] ), 
	.D(n3020), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[152][5]  (.Q(\ram[152][5] ), 
	.D(n3019), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[152][4]  (.Q(\ram[152][4] ), 
	.D(n3018), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[152][3]  (.Q(\ram[152][3] ), 
	.D(n3017), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][2]  (.Q(\ram[152][2] ), 
	.D(n3016), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][1]  (.Q(\ram[152][1] ), 
	.D(n3015), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][0]  (.Q(\ram[152][0] ), 
	.D(n3014), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[148][15]  (.Q(\ram[148][15] ), 
	.D(n2965), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][14]  (.Q(\ram[148][14] ), 
	.D(n2964), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][13]  (.Q(\ram[148][13] ), 
	.D(n2963), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][12]  (.Q(\ram[148][12] ), 
	.D(n2962), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][11]  (.Q(\ram[148][11] ), 
	.D(n2961), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][10]  (.Q(\ram[148][10] ), 
	.D(n2960), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[148][9]  (.Q(\ram[148][9] ), 
	.D(n2959), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[148][8]  (.Q(\ram[148][8] ), 
	.D(n2958), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[148][7]  (.Q(\ram[148][7] ), 
	.D(n2957), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[148][6]  (.Q(\ram[148][6] ), 
	.D(n2956), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[148][5]  (.Q(\ram[148][5] ), 
	.D(n2955), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[148][4]  (.Q(\ram[148][4] ), 
	.D(n2954), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[148][3]  (.Q(\ram[148][3] ), 
	.D(n2953), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[148][2]  (.Q(\ram[148][2] ), 
	.D(n2952), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[148][1]  (.Q(\ram[148][1] ), 
	.D(n2951), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[148][0]  (.Q(\ram[148][0] ), 
	.D(n2950), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[144][15]  (.Q(\ram[144][15] ), 
	.D(n2901), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[144][14]  (.Q(\ram[144][14] ), 
	.D(n2900), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][13]  (.Q(\ram[144][13] ), 
	.D(n2899), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[144][12]  (.Q(\ram[144][12] ), 
	.D(n2898), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[144][11]  (.Q(\ram[144][11] ), 
	.D(n2897), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][10]  (.Q(\ram[144][10] ), 
	.D(n2896), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[144][9]  (.Q(\ram[144][9] ), 
	.D(n2895), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][8]  (.Q(\ram[144][8] ), 
	.D(n2894), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][7]  (.Q(\ram[144][7] ), 
	.D(n2893), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][6]  (.Q(\ram[144][6] ), 
	.D(n2892), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][5]  (.Q(\ram[144][5] ), 
	.D(n2891), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][4]  (.Q(\ram[144][4] ), 
	.D(n2890), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][3]  (.Q(\ram[144][3] ), 
	.D(n2889), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][2]  (.Q(\ram[144][2] ), 
	.D(n2888), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[144][1]  (.Q(\ram[144][1] ), 
	.D(n2887), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[144][0]  (.Q(\ram[144][0] ), 
	.D(n2886), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[140][15]  (.Q(\ram[140][15] ), 
	.D(n2837), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][14]  (.Q(\ram[140][14] ), 
	.D(n2836), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][13]  (.Q(\ram[140][13] ), 
	.D(n2835), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][12]  (.Q(\ram[140][12] ), 
	.D(n2834), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[140][11]  (.Q(\ram[140][11] ), 
	.D(n2833), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[140][10]  (.Q(\ram[140][10] ), 
	.D(n2832), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[140][9]  (.Q(\ram[140][9] ), 
	.D(n2831), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[140][8]  (.Q(\ram[140][8] ), 
	.D(n2830), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][7]  (.Q(\ram[140][7] ), 
	.D(n2829), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[140][6]  (.Q(\ram[140][6] ), 
	.D(n2828), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[140][5]  (.Q(\ram[140][5] ), 
	.D(n2827), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[140][4]  (.Q(\ram[140][4] ), 
	.D(n2826), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[140][3]  (.Q(\ram[140][3] ), 
	.D(n2825), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[140][2]  (.Q(\ram[140][2] ), 
	.D(n2824), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[140][1]  (.Q(\ram[140][1] ), 
	.D(n2823), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[140][0]  (.Q(\ram[140][0] ), 
	.D(n2822), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[136][15]  (.Q(\ram[136][15] ), 
	.D(n2773), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][14]  (.Q(\ram[136][14] ), 
	.D(n2772), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][13]  (.Q(\ram[136][13] ), 
	.D(n2771), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[136][12]  (.Q(\ram[136][12] ), 
	.D(n2770), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][11]  (.Q(\ram[136][11] ), 
	.D(n2769), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][10]  (.Q(\ram[136][10] ), 
	.D(n2768), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[136][9]  (.Q(\ram[136][9] ), 
	.D(n2767), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][8]  (.Q(\ram[136][8] ), 
	.D(n2766), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][7]  (.Q(\ram[136][7] ), 
	.D(n2765), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[136][6]  (.Q(\ram[136][6] ), 
	.D(n2764), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[136][5]  (.Q(\ram[136][5] ), 
	.D(n2763), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[136][4]  (.Q(\ram[136][4] ), 
	.D(n2762), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[136][3]  (.Q(\ram[136][3] ), 
	.D(n2761), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[136][2]  (.Q(\ram[136][2] ), 
	.D(n2760), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[136][1]  (.Q(\ram[136][1] ), 
	.D(n2759), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[136][0]  (.Q(\ram[136][0] ), 
	.D(n2758), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[132][15]  (.Q(\ram[132][15] ), 
	.D(n2709), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[132][14]  (.Q(\ram[132][14] ), 
	.D(n2708), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[132][13]  (.Q(\ram[132][13] ), 
	.D(n2707), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[132][12]  (.Q(\ram[132][12] ), 
	.D(n2706), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[132][11]  (.Q(\ram[132][11] ), 
	.D(n2705), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[132][10]  (.Q(\ram[132][10] ), 
	.D(n2704), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[132][9]  (.Q(\ram[132][9] ), 
	.D(n2703), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[132][8]  (.Q(\ram[132][8] ), 
	.D(n2702), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[132][7]  (.Q(\ram[132][7] ), 
	.D(n2701), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[132][6]  (.Q(\ram[132][6] ), 
	.D(n2700), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[132][5]  (.Q(\ram[132][5] ), 
	.D(n2699), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[132][4]  (.Q(\ram[132][4] ), 
	.D(n2698), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[132][3]  (.Q(\ram[132][3] ), 
	.D(n2697), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[132][2]  (.Q(\ram[132][2] ), 
	.D(n2696), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[132][1]  (.Q(\ram[132][1] ), 
	.D(n2695), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[132][0]  (.Q(\ram[132][0] ), 
	.D(n2694), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[128][15]  (.Q(\ram[128][15] ), 
	.D(n2645), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][14]  (.Q(\ram[128][14] ), 
	.D(n2644), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][13]  (.Q(\ram[128][13] ), 
	.D(n2643), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][12]  (.Q(\ram[128][12] ), 
	.D(n2642), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[128][11]  (.Q(\ram[128][11] ), 
	.D(n2641), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[128][10]  (.Q(\ram[128][10] ), 
	.D(n2640), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[128][9]  (.Q(\ram[128][9] ), 
	.D(n2639), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][8]  (.Q(\ram[128][8] ), 
	.D(n2638), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[128][7]  (.Q(\ram[128][7] ), 
	.D(n2637), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[128][6]  (.Q(\ram[128][6] ), 
	.D(n2636), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][5]  (.Q(\ram[128][5] ), 
	.D(n2635), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][4]  (.Q(\ram[128][4] ), 
	.D(n2634), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][3]  (.Q(\ram[128][3] ), 
	.D(n2633), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][2]  (.Q(\ram[128][2] ), 
	.D(n2632), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[128][1]  (.Q(\ram[128][1] ), 
	.D(n2631), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][0]  (.Q(\ram[128][0] ), 
	.D(n2630), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[124][15]  (.Q(\ram[124][15] ), 
	.D(n2581), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[124][14]  (.Q(\ram[124][14] ), 
	.D(n2580), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[124][13]  (.Q(\ram[124][13] ), 
	.D(n2579), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[124][12]  (.Q(\ram[124][12] ), 
	.D(n2578), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[124][11]  (.Q(\ram[124][11] ), 
	.D(n2577), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[124][10]  (.Q(\ram[124][10] ), 
	.D(n2576), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[124][9]  (.Q(\ram[124][9] ), 
	.D(n2575), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[124][8]  (.Q(\ram[124][8] ), 
	.D(n2574), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[124][7]  (.Q(\ram[124][7] ), 
	.D(n2573), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[124][6]  (.Q(\ram[124][6] ), 
	.D(n2572), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][5]  (.Q(\ram[124][5] ), 
	.D(n2571), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][4]  (.Q(\ram[124][4] ), 
	.D(n2570), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][3]  (.Q(\ram[124][3] ), 
	.D(n2569), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[124][2]  (.Q(\ram[124][2] ), 
	.D(n2568), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][1]  (.Q(\ram[124][1] ), 
	.D(n2567), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[124][0]  (.Q(\ram[124][0] ), 
	.D(n2566), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[120][15]  (.Q(\ram[120][15] ), 
	.D(n2517), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[120][14]  (.Q(\ram[120][14] ), 
	.D(n2516), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[120][13]  (.Q(\ram[120][13] ), 
	.D(n2515), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[120][12]  (.Q(\ram[120][12] ), 
	.D(n2514), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[120][11]  (.Q(\ram[120][11] ), 
	.D(n2513), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[120][10]  (.Q(\ram[120][10] ), 
	.D(n2512), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][9]  (.Q(\ram[120][9] ), 
	.D(n2511), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][8]  (.Q(\ram[120][8] ), 
	.D(n2510), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][7]  (.Q(\ram[120][7] ), 
	.D(n2509), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][6]  (.Q(\ram[120][6] ), 
	.D(n2508), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[120][5]  (.Q(\ram[120][5] ), 
	.D(n2507), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[120][4]  (.Q(\ram[120][4] ), 
	.D(n2506), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[120][3]  (.Q(\ram[120][3] ), 
	.D(n2505), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[120][2]  (.Q(\ram[120][2] ), 
	.D(n2504), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[120][1]  (.Q(\ram[120][1] ), 
	.D(n2503), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[120][0]  (.Q(\ram[120][0] ), 
	.D(n2502), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[116][15]  (.Q(\ram[116][15] ), 
	.D(n2453), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][14]  (.Q(\ram[116][14] ), 
	.D(n2452), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][13]  (.Q(\ram[116][13] ), 
	.D(n2451), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[116][12]  (.Q(\ram[116][12] ), 
	.D(n2450), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[116][11]  (.Q(\ram[116][11] ), 
	.D(n2449), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][10]  (.Q(\ram[116][10] ), 
	.D(n2448), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[116][9]  (.Q(\ram[116][9] ), 
	.D(n2447), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][8]  (.Q(\ram[116][8] ), 
	.D(n2446), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][7]  (.Q(\ram[116][7] ), 
	.D(n2445), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][6]  (.Q(\ram[116][6] ), 
	.D(n2444), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][5]  (.Q(\ram[116][5] ), 
	.D(n2443), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[116][4]  (.Q(\ram[116][4] ), 
	.D(n2442), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][3]  (.Q(\ram[116][3] ), 
	.D(n2441), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][2]  (.Q(\ram[116][2] ), 
	.D(n2440), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][1]  (.Q(\ram[116][1] ), 
	.D(n2439), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][0]  (.Q(\ram[116][0] ), 
	.D(n2438), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[112][15]  (.Q(\ram[112][15] ), 
	.D(n2389), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][14]  (.Q(\ram[112][14] ), 
	.D(n2388), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[112][13]  (.Q(\ram[112][13] ), 
	.D(n2387), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[112][12]  (.Q(\ram[112][12] ), 
	.D(n2386), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][11]  (.Q(\ram[112][11] ), 
	.D(n2385), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][10]  (.Q(\ram[112][10] ), 
	.D(n2384), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][9]  (.Q(\ram[112][9] ), 
	.D(n2383), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][8]  (.Q(\ram[112][8] ), 
	.D(n2382), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][7]  (.Q(\ram[112][7] ), 
	.D(n2381), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][6]  (.Q(\ram[112][6] ), 
	.D(n2380), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][5]  (.Q(\ram[112][5] ), 
	.D(n2379), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][4]  (.Q(\ram[112][4] ), 
	.D(n2378), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][3]  (.Q(\ram[112][3] ), 
	.D(n2377), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][2]  (.Q(\ram[112][2] ), 
	.D(n2376), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][1]  (.Q(\ram[112][1] ), 
	.D(n2375), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][0]  (.Q(\ram[112][0] ), 
	.D(n2374), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[108][15]  (.Q(\ram[108][15] ), 
	.D(n2325), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[108][14]  (.Q(\ram[108][14] ), 
	.D(n2324), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[108][13]  (.Q(\ram[108][13] ), 
	.D(n2323), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[108][12]  (.Q(\ram[108][12] ), 
	.D(n2322), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][11]  (.Q(\ram[108][11] ), 
	.D(n2321), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][10]  (.Q(\ram[108][10] ), 
	.D(n2320), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[108][9]  (.Q(\ram[108][9] ), 
	.D(n2319), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[108][8]  (.Q(\ram[108][8] ), 
	.D(n2318), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][7]  (.Q(\ram[108][7] ), 
	.D(n2317), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[108][6]  (.Q(\ram[108][6] ), 
	.D(n2316), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][5]  (.Q(\ram[108][5] ), 
	.D(n2315), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][4]  (.Q(\ram[108][4] ), 
	.D(n2314), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[108][3]  (.Q(\ram[108][3] ), 
	.D(n2313), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][2]  (.Q(\ram[108][2] ), 
	.D(n2312), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][1]  (.Q(\ram[108][1] ), 
	.D(n2311), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][0]  (.Q(\ram[108][0] ), 
	.D(n2310), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[104][15]  (.Q(\ram[104][15] ), 
	.D(n2261), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][14]  (.Q(\ram[104][14] ), 
	.D(n2260), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][13]  (.Q(\ram[104][13] ), 
	.D(n2259), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][12]  (.Q(\ram[104][12] ), 
	.D(n2258), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][11]  (.Q(\ram[104][11] ), 
	.D(n2257), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][10]  (.Q(\ram[104][10] ), 
	.D(n2256), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][9]  (.Q(\ram[104][9] ), 
	.D(n2255), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][8]  (.Q(\ram[104][8] ), 
	.D(n2254), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[104][7]  (.Q(\ram[104][7] ), 
	.D(n2253), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[104][6]  (.Q(\ram[104][6] ), 
	.D(n2252), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][5]  (.Q(\ram[104][5] ), 
	.D(n2251), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][4]  (.Q(\ram[104][4] ), 
	.D(n2250), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][3]  (.Q(\ram[104][3] ), 
	.D(n2249), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][2]  (.Q(\ram[104][2] ), 
	.D(n2248), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][1]  (.Q(\ram[104][1] ), 
	.D(n2247), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[104][0]  (.Q(\ram[104][0] ), 
	.D(n2246), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[100][15]  (.Q(\ram[100][15] ), 
	.D(n2197), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][14]  (.Q(\ram[100][14] ), 
	.D(n2196), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][13]  (.Q(\ram[100][13] ), 
	.D(n2195), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][12]  (.Q(\ram[100][12] ), 
	.D(n2194), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][11]  (.Q(\ram[100][11] ), 
	.D(n2193), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][10]  (.Q(\ram[100][10] ), 
	.D(n2192), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][9]  (.Q(\ram[100][9] ), 
	.D(n2191), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][8]  (.Q(\ram[100][8] ), 
	.D(n2190), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[100][7]  (.Q(\ram[100][7] ), 
	.D(n2189), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[100][6]  (.Q(\ram[100][6] ), 
	.D(n2188), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][5]  (.Q(\ram[100][5] ), 
	.D(n2187), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][4]  (.Q(\ram[100][4] ), 
	.D(n2186), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][3]  (.Q(\ram[100][3] ), 
	.D(n2185), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][2]  (.Q(\ram[100][2] ), 
	.D(n2184), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][1]  (.Q(\ram[100][1] ), 
	.D(n2183), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[100][0]  (.Q(\ram[100][0] ), 
	.D(n2182), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[96][15]  (.Q(\ram[96][15] ), 
	.D(n2133), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][14]  (.Q(\ram[96][14] ), 
	.D(n2132), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][13]  (.Q(\ram[96][13] ), 
	.D(n2131), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[96][12]  (.Q(\ram[96][12] ), 
	.D(n2130), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[96][11]  (.Q(\ram[96][11] ), 
	.D(n2129), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[96][10]  (.Q(\ram[96][10] ), 
	.D(n2128), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][9]  (.Q(\ram[96][9] ), 
	.D(n2127), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][8]  (.Q(\ram[96][8] ), 
	.D(n2126), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[96][7]  (.Q(\ram[96][7] ), 
	.D(n2125), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][6]  (.Q(\ram[96][6] ), 
	.D(n2124), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][5]  (.Q(\ram[96][5] ), 
	.D(n2123), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[96][4]  (.Q(\ram[96][4] ), 
	.D(n2122), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[96][3]  (.Q(\ram[96][3] ), 
	.D(n2121), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[96][2]  (.Q(\ram[96][2] ), 
	.D(n2120), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[96][1]  (.Q(\ram[96][1] ), 
	.D(n2119), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[96][0]  (.Q(\ram[96][0] ), 
	.D(n2118), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[92][15]  (.Q(\ram[92][15] ), 
	.D(n2069), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[92][14]  (.Q(\ram[92][14] ), 
	.D(n2068), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][13]  (.Q(\ram[92][13] ), 
	.D(n2067), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][12]  (.Q(\ram[92][12] ), 
	.D(n2066), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][11]  (.Q(\ram[92][11] ), 
	.D(n2065), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][10]  (.Q(\ram[92][10] ), 
	.D(n2064), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][9]  (.Q(\ram[92][9] ), 
	.D(n2063), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][8]  (.Q(\ram[92][8] ), 
	.D(n2062), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[92][7]  (.Q(\ram[92][7] ), 
	.D(n2061), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[92][6]  (.Q(\ram[92][6] ), 
	.D(n2060), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][5]  (.Q(\ram[92][5] ), 
	.D(n2059), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[92][4]  (.Q(\ram[92][4] ), 
	.D(n2058), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][3]  (.Q(\ram[92][3] ), 
	.D(n2057), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[92][2]  (.Q(\ram[92][2] ), 
	.D(n2056), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[92][1]  (.Q(\ram[92][1] ), 
	.D(n2055), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][0]  (.Q(\ram[92][0] ), 
	.D(n2054), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[88][15]  (.Q(\ram[88][15] ), 
	.D(n2005), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[88][14]  (.Q(\ram[88][14] ), 
	.D(n2004), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[88][13]  (.Q(\ram[88][13] ), 
	.D(n2003), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[88][12]  (.Q(\ram[88][12] ), 
	.D(n2002), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[88][11]  (.Q(\ram[88][11] ), 
	.D(n2001), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[88][10]  (.Q(\ram[88][10] ), 
	.D(n2000), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[88][9]  (.Q(\ram[88][9] ), 
	.D(n1999), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[88][8]  (.Q(\ram[88][8] ), 
	.D(n1998), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][7]  (.Q(\ram[88][7] ), 
	.D(n1997), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[88][6]  (.Q(\ram[88][6] ), 
	.D(n1996), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][5]  (.Q(\ram[88][5] ), 
	.D(n1995), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][4]  (.Q(\ram[88][4] ), 
	.D(n1994), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[88][3]  (.Q(\ram[88][3] ), 
	.D(n1993), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][2]  (.Q(\ram[88][2] ), 
	.D(n1992), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][1]  (.Q(\ram[88][1] ), 
	.D(n1991), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[88][0]  (.Q(\ram[88][0] ), 
	.D(n1990), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[84][15]  (.Q(\ram[84][15] ), 
	.D(n1941), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][14]  (.Q(\ram[84][14] ), 
	.D(n1940), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][13]  (.Q(\ram[84][13] ), 
	.D(n1939), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[84][12]  (.Q(\ram[84][12] ), 
	.D(n1938), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[84][11]  (.Q(\ram[84][11] ), 
	.D(n1937), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][10]  (.Q(\ram[84][10] ), 
	.D(n1936), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[84][9]  (.Q(\ram[84][9] ), 
	.D(n1935), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][8]  (.Q(\ram[84][8] ), 
	.D(n1934), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[84][7]  (.Q(\ram[84][7] ), 
	.D(n1933), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[84][6]  (.Q(\ram[84][6] ), 
	.D(n1932), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][5]  (.Q(\ram[84][5] ), 
	.D(n1931), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[84][4]  (.Q(\ram[84][4] ), 
	.D(n1930), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][3]  (.Q(\ram[84][3] ), 
	.D(n1929), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][2]  (.Q(\ram[84][2] ), 
	.D(n1928), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][1]  (.Q(\ram[84][1] ), 
	.D(n1927), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[84][0]  (.Q(\ram[84][0] ), 
	.D(n1926), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[80][15]  (.Q(\ram[80][15] ), 
	.D(n1877), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][14]  (.Q(\ram[80][14] ), 
	.D(n1876), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][13]  (.Q(\ram[80][13] ), 
	.D(n1875), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][12]  (.Q(\ram[80][12] ), 
	.D(n1874), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][11]  (.Q(\ram[80][11] ), 
	.D(n1873), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][10]  (.Q(\ram[80][10] ), 
	.D(n1872), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[80][9]  (.Q(\ram[80][9] ), 
	.D(n1871), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[80][8]  (.Q(\ram[80][8] ), 
	.D(n1870), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[80][7]  (.Q(\ram[80][7] ), 
	.D(n1869), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[80][6]  (.Q(\ram[80][6] ), 
	.D(n1868), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][5]  (.Q(\ram[80][5] ), 
	.D(n1867), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][4]  (.Q(\ram[80][4] ), 
	.D(n1866), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][3]  (.Q(\ram[80][3] ), 
	.D(n1865), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][2]  (.Q(\ram[80][2] ), 
	.D(n1864), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][1]  (.Q(\ram[80][1] ), 
	.D(n1863), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[80][0]  (.Q(\ram[80][0] ), 
	.D(n1862), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[76][15]  (.Q(\ram[76][15] ), 
	.D(n1813), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][14]  (.Q(\ram[76][14] ), 
	.D(n1812), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[76][13]  (.Q(\ram[76][13] ), 
	.D(n1811), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[76][12]  (.Q(\ram[76][12] ), 
	.D(n1810), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[76][11]  (.Q(\ram[76][11] ), 
	.D(n1809), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][10]  (.Q(\ram[76][10] ), 
	.D(n1808), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][9]  (.Q(\ram[76][9] ), 
	.D(n1807), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][8]  (.Q(\ram[76][8] ), 
	.D(n1806), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[76][7]  (.Q(\ram[76][7] ), 
	.D(n1805), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[76][6]  (.Q(\ram[76][6] ), 
	.D(n1804), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][5]  (.Q(\ram[76][5] ), 
	.D(n1803), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[76][4]  (.Q(\ram[76][4] ), 
	.D(n1802), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][3]  (.Q(\ram[76][3] ), 
	.D(n1801), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][2]  (.Q(\ram[76][2] ), 
	.D(n1800), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][1]  (.Q(\ram[76][1] ), 
	.D(n1799), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][0]  (.Q(\ram[76][0] ), 
	.D(n1798), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[72][15]  (.Q(\ram[72][15] ), 
	.D(n1749), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][14]  (.Q(\ram[72][14] ), 
	.D(n1748), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][13]  (.Q(\ram[72][13] ), 
	.D(n1747), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[72][12]  (.Q(\ram[72][12] ), 
	.D(n1746), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][11]  (.Q(\ram[72][11] ), 
	.D(n1745), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][10]  (.Q(\ram[72][10] ), 
	.D(n1744), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][9]  (.Q(\ram[72][9] ), 
	.D(n1743), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][8]  (.Q(\ram[72][8] ), 
	.D(n1742), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[72][7]  (.Q(\ram[72][7] ), 
	.D(n1741), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][6]  (.Q(\ram[72][6] ), 
	.D(n1740), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][5]  (.Q(\ram[72][5] ), 
	.D(n1739), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][4]  (.Q(\ram[72][4] ), 
	.D(n1738), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][3]  (.Q(\ram[72][3] ), 
	.D(n1737), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[72][2]  (.Q(\ram[72][2] ), 
	.D(n1736), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][1]  (.Q(\ram[72][1] ), 
	.D(n1735), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][0]  (.Q(\ram[72][0] ), 
	.D(n1734), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[68][15]  (.Q(\ram[68][15] ), 
	.D(n1685), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][14]  (.Q(\ram[68][14] ), 
	.D(n1684), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][13]  (.Q(\ram[68][13] ), 
	.D(n1683), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][12]  (.Q(\ram[68][12] ), 
	.D(n1682), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][11]  (.Q(\ram[68][11] ), 
	.D(n1681), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][10]  (.Q(\ram[68][10] ), 
	.D(n1680), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][9]  (.Q(\ram[68][9] ), 
	.D(n1679), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][8]  (.Q(\ram[68][8] ), 
	.D(n1678), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][7]  (.Q(\ram[68][7] ), 
	.D(n1677), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[68][6]  (.Q(\ram[68][6] ), 
	.D(n1676), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][5]  (.Q(\ram[68][5] ), 
	.D(n1675), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][4]  (.Q(\ram[68][4] ), 
	.D(n1674), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][3]  (.Q(\ram[68][3] ), 
	.D(n1673), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][2]  (.Q(\ram[68][2] ), 
	.D(n1672), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][1]  (.Q(\ram[68][1] ), 
	.D(n1671), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[68][0]  (.Q(\ram[68][0] ), 
	.D(n1670), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[64][15]  (.Q(\ram[64][15] ), 
	.D(n1621), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][14]  (.Q(\ram[64][14] ), 
	.D(n1620), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][13]  (.Q(\ram[64][13] ), 
	.D(n1619), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[64][12]  (.Q(\ram[64][12] ), 
	.D(n1618), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[64][11]  (.Q(\ram[64][11] ), 
	.D(n1617), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][10]  (.Q(\ram[64][10] ), 
	.D(n1616), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][9]  (.Q(\ram[64][9] ), 
	.D(n1615), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[64][8]  (.Q(\ram[64][8] ), 
	.D(n1614), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][7]  (.Q(\ram[64][7] ), 
	.D(n1613), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[64][6]  (.Q(\ram[64][6] ), 
	.D(n1612), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][5]  (.Q(\ram[64][5] ), 
	.D(n1611), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][4]  (.Q(\ram[64][4] ), 
	.D(n1610), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][3]  (.Q(\ram[64][3] ), 
	.D(n1609), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][2]  (.Q(\ram[64][2] ), 
	.D(n1608), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][1]  (.Q(\ram[64][1] ), 
	.D(n1607), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][0]  (.Q(\ram[64][0] ), 
	.D(n1606), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[60][15]  (.Q(\ram[60][15] ), 
	.D(n1557), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][14]  (.Q(\ram[60][14] ), 
	.D(n1556), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][13]  (.Q(\ram[60][13] ), 
	.D(n1555), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[60][12]  (.Q(\ram[60][12] ), 
	.D(n1554), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][11]  (.Q(\ram[60][11] ), 
	.D(n1553), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][10]  (.Q(\ram[60][10] ), 
	.D(n1552), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][9]  (.Q(\ram[60][9] ), 
	.D(n1551), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[60][8]  (.Q(\ram[60][8] ), 
	.D(n1550), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[60][7]  (.Q(\ram[60][7] ), 
	.D(n1549), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[60][6]  (.Q(\ram[60][6] ), 
	.D(n1548), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][5]  (.Q(\ram[60][5] ), 
	.D(n1547), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][4]  (.Q(\ram[60][4] ), 
	.D(n1546), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][3]  (.Q(\ram[60][3] ), 
	.D(n1545), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][2]  (.Q(\ram[60][2] ), 
	.D(n1544), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][1]  (.Q(\ram[60][1] ), 
	.D(n1543), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[60][0]  (.Q(\ram[60][0] ), 
	.D(n1542), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[56][15]  (.Q(\ram[56][15] ), 
	.D(n1493), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[56][14]  (.Q(\ram[56][14] ), 
	.D(n1492), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[56][13]  (.Q(\ram[56][13] ), 
	.D(n1491), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][12]  (.Q(\ram[56][12] ), 
	.D(n1490), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[56][11]  (.Q(\ram[56][11] ), 
	.D(n1489), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][10]  (.Q(\ram[56][10] ), 
	.D(n1488), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][9]  (.Q(\ram[56][9] ), 
	.D(n1487), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[56][8]  (.Q(\ram[56][8] ), 
	.D(n1486), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[56][7]  (.Q(\ram[56][7] ), 
	.D(n1485), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][6]  (.Q(\ram[56][6] ), 
	.D(n1484), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[56][5]  (.Q(\ram[56][5] ), 
	.D(n1483), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][4]  (.Q(\ram[56][4] ), 
	.D(n1482), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[56][3]  (.Q(\ram[56][3] ), 
	.D(n1481), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][2]  (.Q(\ram[56][2] ), 
	.D(n1480), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[56][1]  (.Q(\ram[56][1] ), 
	.D(n1479), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[56][0]  (.Q(\ram[56][0] ), 
	.D(n1478), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[52][15]  (.Q(\ram[52][15] ), 
	.D(n1429), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][14]  (.Q(\ram[52][14] ), 
	.D(n1428), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][13]  (.Q(\ram[52][13] ), 
	.D(n1427), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][12]  (.Q(\ram[52][12] ), 
	.D(n1426), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][11]  (.Q(\ram[52][11] ), 
	.D(n1425), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][10]  (.Q(\ram[52][10] ), 
	.D(n1424), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][9]  (.Q(\ram[52][9] ), 
	.D(n1423), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][8]  (.Q(\ram[52][8] ), 
	.D(n1422), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][7]  (.Q(\ram[52][7] ), 
	.D(n1421), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][6]  (.Q(\ram[52][6] ), 
	.D(n1420), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][5]  (.Q(\ram[52][5] ), 
	.D(n1419), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][4]  (.Q(\ram[52][4] ), 
	.D(n1418), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][3]  (.Q(\ram[52][3] ), 
	.D(n1417), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][2]  (.Q(\ram[52][2] ), 
	.D(n1416), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][1]  (.Q(\ram[52][1] ), 
	.D(n1415), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][0]  (.Q(\ram[52][0] ), 
	.D(n1414), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[48][15]  (.Q(\ram[48][15] ), 
	.D(n1365), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[48][14]  (.Q(\ram[48][14] ), 
	.D(n1364), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[48][13]  (.Q(\ram[48][13] ), 
	.D(n1363), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][12]  (.Q(\ram[48][12] ), 
	.D(n1362), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][11]  (.Q(\ram[48][11] ), 
	.D(n1361), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][10]  (.Q(\ram[48][10] ), 
	.D(n1360), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][9]  (.Q(\ram[48][9] ), 
	.D(n1359), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[48][8]  (.Q(\ram[48][8] ), 
	.D(n1358), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[48][7]  (.Q(\ram[48][7] ), 
	.D(n1357), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[48][6]  (.Q(\ram[48][6] ), 
	.D(n1356), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[48][5]  (.Q(\ram[48][5] ), 
	.D(n1355), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][4]  (.Q(\ram[48][4] ), 
	.D(n1354), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][3]  (.Q(\ram[48][3] ), 
	.D(n1353), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][2]  (.Q(\ram[48][2] ), 
	.D(n1352), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[48][1]  (.Q(\ram[48][1] ), 
	.D(n1351), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[48][0]  (.Q(\ram[48][0] ), 
	.D(n1350), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[44][15]  (.Q(\ram[44][15] ), 
	.D(n1301), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[44][14]  (.Q(\ram[44][14] ), 
	.D(n1300), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][13]  (.Q(\ram[44][13] ), 
	.D(n1299), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[44][12]  (.Q(\ram[44][12] ), 
	.D(n1298), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[44][11]  (.Q(\ram[44][11] ), 
	.D(n1297), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][10]  (.Q(\ram[44][10] ), 
	.D(n1296), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[44][9]  (.Q(\ram[44][9] ), 
	.D(n1295), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[44][8]  (.Q(\ram[44][8] ), 
	.D(n1294), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[44][7]  (.Q(\ram[44][7] ), 
	.D(n1293), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[44][6]  (.Q(\ram[44][6] ), 
	.D(n1292), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][5]  (.Q(\ram[44][5] ), 
	.D(n1291), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][4]  (.Q(\ram[44][4] ), 
	.D(n1290), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][3]  (.Q(\ram[44][3] ), 
	.D(n1289), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][2]  (.Q(\ram[44][2] ), 
	.D(n1288), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][1]  (.Q(\ram[44][1] ), 
	.D(n1287), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][0]  (.Q(\ram[44][0] ), 
	.D(n1286), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[40][15]  (.Q(\ram[40][15] ), 
	.D(n1237), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][14]  (.Q(\ram[40][14] ), 
	.D(n1236), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][13]  (.Q(\ram[40][13] ), 
	.D(n1235), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][12]  (.Q(\ram[40][12] ), 
	.D(n1234), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[40][11]  (.Q(\ram[40][11] ), 
	.D(n1233), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[40][10]  (.Q(\ram[40][10] ), 
	.D(n1232), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][9]  (.Q(\ram[40][9] ), 
	.D(n1231), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][8]  (.Q(\ram[40][8] ), 
	.D(n1230), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][7]  (.Q(\ram[40][7] ), 
	.D(n1229), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[40][6]  (.Q(\ram[40][6] ), 
	.D(n1228), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[40][5]  (.Q(\ram[40][5] ), 
	.D(n1227), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[40][4]  (.Q(\ram[40][4] ), 
	.D(n1226), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][3]  (.Q(\ram[40][3] ), 
	.D(n1225), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[40][2]  (.Q(\ram[40][2] ), 
	.D(n1224), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][1]  (.Q(\ram[40][1] ), 
	.D(n1223), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][0]  (.Q(\ram[40][0] ), 
	.D(n1222), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[36][15]  (.Q(\ram[36][15] ), 
	.D(n1173), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][14]  (.Q(\ram[36][14] ), 
	.D(n1172), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[36][13]  (.Q(\ram[36][13] ), 
	.D(n1171), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[36][12]  (.Q(\ram[36][12] ), 
	.D(n1170), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[36][11]  (.Q(\ram[36][11] ), 
	.D(n1169), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][10]  (.Q(\ram[36][10] ), 
	.D(n1168), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][9]  (.Q(\ram[36][9] ), 
	.D(n1167), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][8]  (.Q(\ram[36][8] ), 
	.D(n1166), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][7]  (.Q(\ram[36][7] ), 
	.D(n1165), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][6]  (.Q(\ram[36][6] ), 
	.D(n1164), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][5]  (.Q(\ram[36][5] ), 
	.D(n1163), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[36][4]  (.Q(\ram[36][4] ), 
	.D(n1162), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[36][3]  (.Q(\ram[36][3] ), 
	.D(n1161), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][2]  (.Q(\ram[36][2] ), 
	.D(n1160), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[36][1]  (.Q(\ram[36][1] ), 
	.D(n1159), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[36][0]  (.Q(\ram[36][0] ), 
	.D(n1158), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[32][15]  (.Q(\ram[32][15] ), 
	.D(n1109), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][14]  (.Q(\ram[32][14] ), 
	.D(n1108), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][13]  (.Q(\ram[32][13] ), 
	.D(n1107), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][12]  (.Q(\ram[32][12] ), 
	.D(n1106), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[32][11]  (.Q(\ram[32][11] ), 
	.D(n1105), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][10]  (.Q(\ram[32][10] ), 
	.D(n1104), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[32][9]  (.Q(\ram[32][9] ), 
	.D(n1103), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][8]  (.Q(\ram[32][8] ), 
	.D(n1102), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][7]  (.Q(\ram[32][7] ), 
	.D(n1101), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][6]  (.Q(\ram[32][6] ), 
	.D(n1100), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][5]  (.Q(\ram[32][5] ), 
	.D(n1099), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][4]  (.Q(\ram[32][4] ), 
	.D(n1098), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][3]  (.Q(\ram[32][3] ), 
	.D(n1097), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][2]  (.Q(\ram[32][2] ), 
	.D(n1096), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][1]  (.Q(\ram[32][1] ), 
	.D(n1095), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[32][0]  (.Q(\ram[32][0] ), 
	.D(n1094), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[28][15]  (.Q(\ram[28][15] ), 
	.D(n1045), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[28][14]  (.Q(\ram[28][14] ), 
	.D(n1044), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[28][13]  (.Q(\ram[28][13] ), 
	.D(n1043), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[28][12]  (.Q(\ram[28][12] ), 
	.D(n1042), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[28][11]  (.Q(\ram[28][11] ), 
	.D(n1041), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][10]  (.Q(\ram[28][10] ), 
	.D(n1040), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[28][9]  (.Q(\ram[28][9] ), 
	.D(n1039), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[28][8]  (.Q(\ram[28][8] ), 
	.D(n1038), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][7]  (.Q(\ram[28][7] ), 
	.D(n1037), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[28][6]  (.Q(\ram[28][6] ), 
	.D(n1036), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[28][5]  (.Q(\ram[28][5] ), 
	.D(n1035), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][4]  (.Q(\ram[28][4] ), 
	.D(n1034), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[28][3]  (.Q(\ram[28][3] ), 
	.D(n1033), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[28][2]  (.Q(\ram[28][2] ), 
	.D(n1032), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[28][1]  (.Q(\ram[28][1] ), 
	.D(n1031), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][0]  (.Q(\ram[28][0] ), 
	.D(n1030), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[24][15]  (.Q(\ram[24][15] ), 
	.D(n981), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][14]  (.Q(\ram[24][14] ), 
	.D(n980), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][13]  (.Q(\ram[24][13] ), 
	.D(n979), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[24][12]  (.Q(\ram[24][12] ), 
	.D(n978), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[24][11]  (.Q(\ram[24][11] ), 
	.D(n977), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[24][10]  (.Q(\ram[24][10] ), 
	.D(n976), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[24][9]  (.Q(\ram[24][9] ), 
	.D(n975), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[24][8]  (.Q(\ram[24][8] ), 
	.D(n974), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][7]  (.Q(\ram[24][7] ), 
	.D(n973), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][6]  (.Q(\ram[24][6] ), 
	.D(n972), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[24][5]  (.Q(\ram[24][5] ), 
	.D(n971), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[24][4]  (.Q(\ram[24][4] ), 
	.D(n970), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[24][3]  (.Q(\ram[24][3] ), 
	.D(n969), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][2]  (.Q(\ram[24][2] ), 
	.D(n968), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[24][1]  (.Q(\ram[24][1] ), 
	.D(n967), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][0]  (.Q(\ram[24][0] ), 
	.D(n966), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[20][15]  (.Q(\ram[20][15] ), 
	.D(n917), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][14]  (.Q(\ram[20][14] ), 
	.D(n916), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][13]  (.Q(\ram[20][13] ), 
	.D(n915), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][12]  (.Q(\ram[20][12] ), 
	.D(n914), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][11]  (.Q(\ram[20][11] ), 
	.D(n913), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][10]  (.Q(\ram[20][10] ), 
	.D(n912), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[20][9]  (.Q(\ram[20][9] ), 
	.D(n911), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][8]  (.Q(\ram[20][8] ), 
	.D(n910), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][7]  (.Q(\ram[20][7] ), 
	.D(n909), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][6]  (.Q(\ram[20][6] ), 
	.D(n908), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][5]  (.Q(\ram[20][5] ), 
	.D(n907), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[20][4]  (.Q(\ram[20][4] ), 
	.D(n906), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[20][3]  (.Q(\ram[20][3] ), 
	.D(n905), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][2]  (.Q(\ram[20][2] ), 
	.D(n904), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][1]  (.Q(\ram[20][1] ), 
	.D(n903), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][0]  (.Q(\ram[20][0] ), 
	.D(n902), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[16][15]  (.Q(\ram[16][15] ), 
	.D(n853), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[16][14]  (.Q(\ram[16][14] ), 
	.D(n852), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][13]  (.Q(\ram[16][13] ), 
	.D(n851), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[16][12]  (.Q(\ram[16][12] ), 
	.D(n850), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[16][11]  (.Q(\ram[16][11] ), 
	.D(n849), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][10]  (.Q(\ram[16][10] ), 
	.D(n848), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][9]  (.Q(\ram[16][9] ), 
	.D(n847), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][8]  (.Q(\ram[16][8] ), 
	.D(n846), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][7]  (.Q(\ram[16][7] ), 
	.D(n845), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][6]  (.Q(\ram[16][6] ), 
	.D(n844), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[16][5]  (.Q(\ram[16][5] ), 
	.D(n843), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[16][4]  (.Q(\ram[16][4] ), 
	.D(n842), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[16][3]  (.Q(\ram[16][3] ), 
	.D(n841), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[16][2]  (.Q(\ram[16][2] ), 
	.D(n840), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[16][1]  (.Q(\ram[16][1] ), 
	.D(n839), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[16][0]  (.Q(\ram[16][0] ), 
	.D(n838), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[12][15]  (.Q(\ram[12][15] ), 
	.D(n789), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[12][14]  (.Q(\ram[12][14] ), 
	.D(n788), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[12][13]  (.Q(\ram[12][13] ), 
	.D(n787), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][12]  (.Q(\ram[12][12] ), 
	.D(n786), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[12][11]  (.Q(\ram[12][11] ), 
	.D(n785), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][10]  (.Q(\ram[12][10] ), 
	.D(n784), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[12][9]  (.Q(\ram[12][9] ), 
	.D(n783), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][8]  (.Q(\ram[12][8] ), 
	.D(n782), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][7]  (.Q(\ram[12][7] ), 
	.D(n781), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][6]  (.Q(\ram[12][6] ), 
	.D(n780), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][5]  (.Q(\ram[12][5] ), 
	.D(n779), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][4]  (.Q(\ram[12][4] ), 
	.D(n778), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][3]  (.Q(\ram[12][3] ), 
	.D(n777), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][2]  (.Q(\ram[12][2] ), 
	.D(n776), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][1]  (.Q(\ram[12][1] ), 
	.D(n775), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[12][0]  (.Q(\ram[12][0] ), 
	.D(n774), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[8][15]  (.Q(\ram[8][15] ), 
	.D(n725), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[8][14]  (.Q(\ram[8][14] ), 
	.D(n724), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[8][13]  (.Q(\ram[8][13] ), 
	.D(n723), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[8][12]  (.Q(\ram[8][12] ), 
	.D(n722), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[8][11]  (.Q(\ram[8][11] ), 
	.D(n721), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][10]  (.Q(\ram[8][10] ), 
	.D(n720), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[8][9]  (.Q(\ram[8][9] ), 
	.D(n719), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][8]  (.Q(\ram[8][8] ), 
	.D(n718), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[8][7]  (.Q(\ram[8][7] ), 
	.D(n717), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[8][6]  (.Q(\ram[8][6] ), 
	.D(n716), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[8][5]  (.Q(\ram[8][5] ), 
	.D(n715), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][4]  (.Q(\ram[8][4] ), 
	.D(n714), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[8][3]  (.Q(\ram[8][3] ), 
	.D(n713), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][2]  (.Q(\ram[8][2] ), 
	.D(n712), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[8][1]  (.Q(\ram[8][1] ), 
	.D(n711), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[8][0]  (.Q(\ram[8][0] ), 
	.D(n710), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[4][15]  (.Q(\ram[4][15] ), 
	.D(n661), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[4][14]  (.Q(\ram[4][14] ), 
	.D(n660), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[4][13]  (.Q(\ram[4][13] ), 
	.D(n659), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[4][12]  (.Q(\ram[4][12] ), 
	.D(n658), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[4][11]  (.Q(\ram[4][11] ), 
	.D(n657), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][10]  (.Q(\ram[4][10] ), 
	.D(n656), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[4][9]  (.Q(\ram[4][9] ), 
	.D(n655), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[4][8]  (.Q(\ram[4][8] ), 
	.D(n654), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[4][7]  (.Q(\ram[4][7] ), 
	.D(n653), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[4][6]  (.Q(\ram[4][6] ), 
	.D(n652), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][5]  (.Q(\ram[4][5] ), 
	.D(n651), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][4]  (.Q(\ram[4][4] ), 
	.D(n650), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[4][3]  (.Q(\ram[4][3] ), 
	.D(n649), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][2]  (.Q(\ram[4][2] ), 
	.D(n648), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[4][1]  (.Q(\ram[4][1] ), 
	.D(n647), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[4][0]  (.Q(\ram[4][0] ), 
	.D(n646), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[0][15]  (.Q(\ram[0][15] ), 
	.D(n597), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][14]  (.Q(\ram[0][14] ), 
	.D(n596), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][13]  (.Q(\ram[0][13] ), 
	.D(n595), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[0][12]  (.Q(\ram[0][12] ), 
	.D(n594), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[0][11]  (.Q(\ram[0][11] ), 
	.D(n593), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[0][10]  (.Q(\ram[0][10] ), 
	.D(n592), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[0][9]  (.Q(\ram[0][9] ), 
	.D(n591), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[0][8]  (.Q(\ram[0][8] ), 
	.D(n590), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][7]  (.Q(\ram[0][7] ), 
	.D(n589), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[0][6]  (.Q(\ram[0][6] ), 
	.D(n588), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[0][5]  (.Q(\ram[0][5] ), 
	.D(n587), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[0][4]  (.Q(\ram[0][4] ), 
	.D(n586), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[0][3]  (.Q(\ram[0][3] ), 
	.D(n585), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[0][2]  (.Q(\ram[0][2] ), 
	.D(n584), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][1]  (.Q(\ram[0][1] ), 
	.D(n583), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[0][0]  (.Q(\ram[0][0] ), 
	.D(n582), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[255][15]  (.Q(\ram[255][15] ), 
	.D(n4677), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[255][14]  (.Q(\ram[255][14] ), 
	.D(n4676), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[255][13]  (.Q(\ram[255][13] ), 
	.D(n4675), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][12]  (.Q(\ram[255][12] ), 
	.D(n4674), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[255][11]  (.Q(\ram[255][11] ), 
	.D(n4673), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[255][10]  (.Q(\ram[255][10] ), 
	.D(n4672), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][9]  (.Q(\ram[255][9] ), 
	.D(n4671), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][8]  (.Q(\ram[255][8] ), 
	.D(n4670), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][7]  (.Q(\ram[255][7] ), 
	.D(n4669), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[255][6]  (.Q(\ram[255][6] ), 
	.D(n4668), 
	.CK(clk));
   QDFFEHD \ram_reg[255][5]  (.Q(\ram[255][5] ), 
	.D(n4667), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[255][4]  (.Q(\ram[255][4] ), 
	.D(n4666), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[255][3]  (.Q(\ram[255][3] ), 
	.D(n4665), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][2]  (.Q(\ram[255][2] ), 
	.D(n4664), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[255][1]  (.Q(\ram[255][1] ), 
	.D(n4663), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[255][0]  (.Q(\ram[255][0] ), 
	.D(n4662), 
	.CK(clk));
   QDFFEHD \ram_reg[251][15]  (.Q(\ram[251][15] ), 
	.D(n4613), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][14]  (.Q(\ram[251][14] ), 
	.D(n4612), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][13]  (.Q(\ram[251][13] ), 
	.D(n4611), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][12]  (.Q(\ram[251][12] ), 
	.D(n4610), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][11]  (.Q(\ram[251][11] ), 
	.D(n4609), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][10]  (.Q(\ram[251][10] ), 
	.D(n4608), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][9]  (.Q(\ram[251][9] ), 
	.D(n4607), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][8]  (.Q(\ram[251][8] ), 
	.D(n4606), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][7]  (.Q(\ram[251][7] ), 
	.D(n4605), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][6]  (.Q(\ram[251][6] ), 
	.D(n4604), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][5]  (.Q(\ram[251][5] ), 
	.D(n4603), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][4]  (.Q(\ram[251][4] ), 
	.D(n4602), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][3]  (.Q(\ram[251][3] ), 
	.D(n4601), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[251][2]  (.Q(\ram[251][2] ), 
	.D(n4600), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][1]  (.Q(\ram[251][1] ), 
	.D(n4599), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[251][0]  (.Q(\ram[251][0] ), 
	.D(n4598), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[247][15]  (.Q(\ram[247][15] ), 
	.D(n4549), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][14]  (.Q(\ram[247][14] ), 
	.D(n4548), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[247][13]  (.Q(\ram[247][13] ), 
	.D(n4547), 
	.CK(clk));
   QDFFEHD \ram_reg[247][12]  (.Q(\ram[247][12] ), 
	.D(n4546), 
	.CK(clk));
   QDFFEHD \ram_reg[247][11]  (.Q(\ram[247][11] ), 
	.D(n4545), 
	.CK(clk));
   QDFFEHD \ram_reg[247][10]  (.Q(\ram[247][10] ), 
	.D(n4544), 
	.CK(clk));
   QDFFEHD \ram_reg[247][9]  (.Q(\ram[247][9] ), 
	.D(n4543), 
	.CK(clk));
   QDFFEHD \ram_reg[247][8]  (.Q(\ram[247][8] ), 
	.D(n4542), 
	.CK(clk));
   QDFFEHD \ram_reg[247][7]  (.Q(\ram[247][7] ), 
	.D(n4541), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[247][6]  (.Q(\ram[247][6] ), 
	.D(n4540), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][5]  (.Q(\ram[247][5] ), 
	.D(n4539), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][4]  (.Q(\ram[247][4] ), 
	.D(n4538), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][3]  (.Q(\ram[247][3] ), 
	.D(n4537), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[247][2]  (.Q(\ram[247][2] ), 
	.D(n4536), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][1]  (.Q(\ram[247][1] ), 
	.D(n4535), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[247][0]  (.Q(\ram[247][0] ), 
	.D(n4534), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[243][15]  (.Q(\ram[243][15] ), 
	.D(n4485), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][14]  (.Q(\ram[243][14] ), 
	.D(n4484), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][13]  (.Q(\ram[243][13] ), 
	.D(n4483), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][12]  (.Q(\ram[243][12] ), 
	.D(n4482), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[243][11]  (.Q(\ram[243][11] ), 
	.D(n4481), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[243][10]  (.Q(\ram[243][10] ), 
	.D(n4480), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][9]  (.Q(\ram[243][9] ), 
	.D(n4479), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[243][8]  (.Q(\ram[243][8] ), 
	.D(n4478), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[243][7]  (.Q(\ram[243][7] ), 
	.D(n4477), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[243][6]  (.Q(\ram[243][6] ), 
	.D(n4476), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][5]  (.Q(\ram[243][5] ), 
	.D(n4475), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][4]  (.Q(\ram[243][4] ), 
	.D(n4474), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][3]  (.Q(\ram[243][3] ), 
	.D(n4473), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][2]  (.Q(\ram[243][2] ), 
	.D(n4472), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][1]  (.Q(\ram[243][1] ), 
	.D(n4471), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][0]  (.Q(\ram[243][0] ), 
	.D(n4470), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[239][15]  (.Q(\ram[239][15] ), 
	.D(n4421), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][14]  (.Q(\ram[239][14] ), 
	.D(n4420), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][13]  (.Q(\ram[239][13] ), 
	.D(n4419), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][12]  (.Q(\ram[239][12] ), 
	.D(n4418), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][11]  (.Q(\ram[239][11] ), 
	.D(n4417), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][10]  (.Q(\ram[239][10] ), 
	.D(n4416), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[239][9]  (.Q(\ram[239][9] ), 
	.D(n4415), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[239][8]  (.Q(\ram[239][8] ), 
	.D(n4414), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[239][7]  (.Q(\ram[239][7] ), 
	.D(n4413), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][6]  (.Q(\ram[239][6] ), 
	.D(n4412), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[239][5]  (.Q(\ram[239][5] ), 
	.D(n4411), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][4]  (.Q(\ram[239][4] ), 
	.D(n4410), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][3]  (.Q(\ram[239][3] ), 
	.D(n4409), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[239][2]  (.Q(\ram[239][2] ), 
	.D(n4408), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][1]  (.Q(\ram[239][1] ), 
	.D(n4407), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][0]  (.Q(\ram[239][0] ), 
	.D(n4406), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[235][15]  (.Q(\ram[235][15] ), 
	.D(n4357), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][14]  (.Q(\ram[235][14] ), 
	.D(n4356), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[235][13]  (.Q(\ram[235][13] ), 
	.D(n4355), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[235][12]  (.Q(\ram[235][12] ), 
	.D(n4354), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][11]  (.Q(\ram[235][11] ), 
	.D(n4353), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][10]  (.Q(\ram[235][10] ), 
	.D(n4352), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][9]  (.Q(\ram[235][9] ), 
	.D(n4351), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][8]  (.Q(\ram[235][8] ), 
	.D(n4350), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[235][7]  (.Q(\ram[235][7] ), 
	.D(n4349), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][6]  (.Q(\ram[235][6] ), 
	.D(n4348), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][5]  (.Q(\ram[235][5] ), 
	.D(n4347), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[235][4]  (.Q(\ram[235][4] ), 
	.D(n4346), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][3]  (.Q(\ram[235][3] ), 
	.D(n4345), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][2]  (.Q(\ram[235][2] ), 
	.D(n4344), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][1]  (.Q(\ram[235][1] ), 
	.D(n4343), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[235][0]  (.Q(\ram[235][0] ), 
	.D(n4342), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[231][15]  (.Q(\ram[231][15] ), 
	.D(n4293), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][14]  (.Q(\ram[231][14] ), 
	.D(n4292), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][13]  (.Q(\ram[231][13] ), 
	.D(n4291), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][12]  (.Q(\ram[231][12] ), 
	.D(n4290), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][11]  (.Q(\ram[231][11] ), 
	.D(n4289), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[231][10]  (.Q(\ram[231][10] ), 
	.D(n4288), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][9]  (.Q(\ram[231][9] ), 
	.D(n4287), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][8]  (.Q(\ram[231][8] ), 
	.D(n4286), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[231][7]  (.Q(\ram[231][7] ), 
	.D(n4285), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][6]  (.Q(\ram[231][6] ), 
	.D(n4284), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[231][5]  (.Q(\ram[231][5] ), 
	.D(n4283), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][4]  (.Q(\ram[231][4] ), 
	.D(n4282), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][3]  (.Q(\ram[231][3] ), 
	.D(n4281), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[231][2]  (.Q(\ram[231][2] ), 
	.D(n4280), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[231][1]  (.Q(\ram[231][1] ), 
	.D(n4279), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][0]  (.Q(\ram[231][0] ), 
	.D(n4278), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[227][15]  (.Q(\ram[227][15] ), 
	.D(n4229), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][14]  (.Q(\ram[227][14] ), 
	.D(n4228), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][13]  (.Q(\ram[227][13] ), 
	.D(n4227), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[227][12]  (.Q(\ram[227][12] ), 
	.D(n4226), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][11]  (.Q(\ram[227][11] ), 
	.D(n4225), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][10]  (.Q(\ram[227][10] ), 
	.D(n4224), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[227][9]  (.Q(\ram[227][9] ), 
	.D(n4223), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[227][8]  (.Q(\ram[227][8] ), 
	.D(n4222), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][7]  (.Q(\ram[227][7] ), 
	.D(n4221), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[227][6]  (.Q(\ram[227][6] ), 
	.D(n4220), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][5]  (.Q(\ram[227][5] ), 
	.D(n4219), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[227][4]  (.Q(\ram[227][4] ), 
	.D(n4218), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][3]  (.Q(\ram[227][3] ), 
	.D(n4217), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][2]  (.Q(\ram[227][2] ), 
	.D(n4216), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[227][1]  (.Q(\ram[227][1] ), 
	.D(n4215), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][0]  (.Q(\ram[227][0] ), 
	.D(n4214), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[223][15]  (.Q(\ram[223][15] ), 
	.D(n4165), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[223][14]  (.Q(\ram[223][14] ), 
	.D(n4164), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][13]  (.Q(\ram[223][13] ), 
	.D(n4163), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][12]  (.Q(\ram[223][12] ), 
	.D(n4162), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][11]  (.Q(\ram[223][11] ), 
	.D(n4161), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[223][10]  (.Q(\ram[223][10] ), 
	.D(n4160), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[223][9]  (.Q(\ram[223][9] ), 
	.D(n4159), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][8]  (.Q(\ram[223][8] ), 
	.D(n4158), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][7]  (.Q(\ram[223][7] ), 
	.D(n4157), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[223][6]  (.Q(\ram[223][6] ), 
	.D(n4156), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][5]  (.Q(\ram[223][5] ), 
	.D(n4155), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][4]  (.Q(\ram[223][4] ), 
	.D(n4154), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[223][3]  (.Q(\ram[223][3] ), 
	.D(n4153), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][2]  (.Q(\ram[223][2] ), 
	.D(n4152), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[223][1]  (.Q(\ram[223][1] ), 
	.D(n4151), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][0]  (.Q(\ram[223][0] ), 
	.D(n4150), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[219][15]  (.Q(\ram[219][15] ), 
	.D(n4101), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][14]  (.Q(\ram[219][14] ), 
	.D(n4100), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][13]  (.Q(\ram[219][13] ), 
	.D(n4099), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][12]  (.Q(\ram[219][12] ), 
	.D(n4098), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][11]  (.Q(\ram[219][11] ), 
	.D(n4097), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][10]  (.Q(\ram[219][10] ), 
	.D(n4096), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[219][9]  (.Q(\ram[219][9] ), 
	.D(n4095), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][8]  (.Q(\ram[219][8] ), 
	.D(n4094), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][7]  (.Q(\ram[219][7] ), 
	.D(n4093), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][6]  (.Q(\ram[219][6] ), 
	.D(n4092), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][5]  (.Q(\ram[219][5] ), 
	.D(n4091), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][4]  (.Q(\ram[219][4] ), 
	.D(n4090), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][3]  (.Q(\ram[219][3] ), 
	.D(n4089), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][2]  (.Q(\ram[219][2] ), 
	.D(n4088), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][1]  (.Q(\ram[219][1] ), 
	.D(n4087), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][0]  (.Q(\ram[219][0] ), 
	.D(n4086), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[215][15]  (.Q(\ram[215][15] ), 
	.D(n4037), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][14]  (.Q(\ram[215][14] ), 
	.D(n4036), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][13]  (.Q(\ram[215][13] ), 
	.D(n4035), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[215][12]  (.Q(\ram[215][12] ), 
	.D(n4034), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[215][11]  (.Q(\ram[215][11] ), 
	.D(n4033), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][10]  (.Q(\ram[215][10] ), 
	.D(n4032), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][9]  (.Q(\ram[215][9] ), 
	.D(n4031), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[215][8]  (.Q(\ram[215][8] ), 
	.D(n4030), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[215][7]  (.Q(\ram[215][7] ), 
	.D(n4029), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][6]  (.Q(\ram[215][6] ), 
	.D(n4028), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[215][5]  (.Q(\ram[215][5] ), 
	.D(n4027), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[215][4]  (.Q(\ram[215][4] ), 
	.D(n4026), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][3]  (.Q(\ram[215][3] ), 
	.D(n4025), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][2]  (.Q(\ram[215][2] ), 
	.D(n4024), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][1]  (.Q(\ram[215][1] ), 
	.D(n4023), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][0]  (.Q(\ram[215][0] ), 
	.D(n4022), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[211][15]  (.Q(\ram[211][15] ), 
	.D(n3973), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[211][14]  (.Q(\ram[211][14] ), 
	.D(n3972), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[211][13]  (.Q(\ram[211][13] ), 
	.D(n3971), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][12]  (.Q(\ram[211][12] ), 
	.D(n3970), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][11]  (.Q(\ram[211][11] ), 
	.D(n3969), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[211][10]  (.Q(\ram[211][10] ), 
	.D(n3968), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][9]  (.Q(\ram[211][9] ), 
	.D(n3967), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][8]  (.Q(\ram[211][8] ), 
	.D(n3966), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][7]  (.Q(\ram[211][7] ), 
	.D(n3965), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][6]  (.Q(\ram[211][6] ), 
	.D(n3964), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][5]  (.Q(\ram[211][5] ), 
	.D(n3963), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][4]  (.Q(\ram[211][4] ), 
	.D(n3962), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[211][3]  (.Q(\ram[211][3] ), 
	.D(n3961), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[211][2]  (.Q(\ram[211][2] ), 
	.D(n3960), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][1]  (.Q(\ram[211][1] ), 
	.D(n3959), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[211][0]  (.Q(\ram[211][0] ), 
	.D(n3958), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[207][15]  (.Q(\ram[207][15] ), 
	.D(n3909), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][14]  (.Q(\ram[207][14] ), 
	.D(n3908), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][13]  (.Q(\ram[207][13] ), 
	.D(n3907), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[207][12]  (.Q(\ram[207][12] ), 
	.D(n3906), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][11]  (.Q(\ram[207][11] ), 
	.D(n3905), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][10]  (.Q(\ram[207][10] ), 
	.D(n3904), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][9]  (.Q(\ram[207][9] ), 
	.D(n3903), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[207][8]  (.Q(\ram[207][8] ), 
	.D(n3902), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[207][7]  (.Q(\ram[207][7] ), 
	.D(n3901), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][6]  (.Q(\ram[207][6] ), 
	.D(n3900), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[207][5]  (.Q(\ram[207][5] ), 
	.D(n3899), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][4]  (.Q(\ram[207][4] ), 
	.D(n3898), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][3]  (.Q(\ram[207][3] ), 
	.D(n3897), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][2]  (.Q(\ram[207][2] ), 
	.D(n3896), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][1]  (.Q(\ram[207][1] ), 
	.D(n3895), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][0]  (.Q(\ram[207][0] ), 
	.D(n3894), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[203][15]  (.Q(\ram[203][15] ), 
	.D(n3845), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[203][14]  (.Q(\ram[203][14] ), 
	.D(n3844), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][13]  (.Q(\ram[203][13] ), 
	.D(n3843), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[203][12]  (.Q(\ram[203][12] ), 
	.D(n3842), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[203][11]  (.Q(\ram[203][11] ), 
	.D(n3841), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[203][10]  (.Q(\ram[203][10] ), 
	.D(n3840), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[203][9]  (.Q(\ram[203][9] ), 
	.D(n3839), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][8]  (.Q(\ram[203][8] ), 
	.D(n3838), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][7]  (.Q(\ram[203][7] ), 
	.D(n3837), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][6]  (.Q(\ram[203][6] ), 
	.D(n3836), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][5]  (.Q(\ram[203][5] ), 
	.D(n3835), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][4]  (.Q(\ram[203][4] ), 
	.D(n3834), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][3]  (.Q(\ram[203][3] ), 
	.D(n3833), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][2]  (.Q(\ram[203][2] ), 
	.D(n3832), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][1]  (.Q(\ram[203][1] ), 
	.D(n3831), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][0]  (.Q(\ram[203][0] ), 
	.D(n3830), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[199][15]  (.Q(\ram[199][15] ), 
	.D(n3781), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][14]  (.Q(\ram[199][14] ), 
	.D(n3780), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][13]  (.Q(\ram[199][13] ), 
	.D(n3779), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[199][12]  (.Q(\ram[199][12] ), 
	.D(n3778), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[199][11]  (.Q(\ram[199][11] ), 
	.D(n3777), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][10]  (.Q(\ram[199][10] ), 
	.D(n3776), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[199][9]  (.Q(\ram[199][9] ), 
	.D(n3775), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[199][8]  (.Q(\ram[199][8] ), 
	.D(n3774), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][7]  (.Q(\ram[199][7] ), 
	.D(n3773), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][6]  (.Q(\ram[199][6] ), 
	.D(n3772), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][5]  (.Q(\ram[199][5] ), 
	.D(n3771), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][4]  (.Q(\ram[199][4] ), 
	.D(n3770), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][3]  (.Q(\ram[199][3] ), 
	.D(n3769), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[199][2]  (.Q(\ram[199][2] ), 
	.D(n3768), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][1]  (.Q(\ram[199][1] ), 
	.D(n3767), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][0]  (.Q(\ram[199][0] ), 
	.D(n3766), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[195][15]  (.Q(\ram[195][15] ), 
	.D(n3717), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][14]  (.Q(\ram[195][14] ), 
	.D(n3716), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][13]  (.Q(\ram[195][13] ), 
	.D(n3715), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[195][12]  (.Q(\ram[195][12] ), 
	.D(n3714), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[195][11]  (.Q(\ram[195][11] ), 
	.D(n3713), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][10]  (.Q(\ram[195][10] ), 
	.D(n3712), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][9]  (.Q(\ram[195][9] ), 
	.D(n3711), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][8]  (.Q(\ram[195][8] ), 
	.D(n3710), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[195][7]  (.Q(\ram[195][7] ), 
	.D(n3709), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][6]  (.Q(\ram[195][6] ), 
	.D(n3708), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][5]  (.Q(\ram[195][5] ), 
	.D(n3707), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][4]  (.Q(\ram[195][4] ), 
	.D(n3706), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][3]  (.Q(\ram[195][3] ), 
	.D(n3705), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[195][2]  (.Q(\ram[195][2] ), 
	.D(n3704), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][1]  (.Q(\ram[195][1] ), 
	.D(n3703), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][0]  (.Q(\ram[195][0] ), 
	.D(n3702), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[191][15]  (.Q(\ram[191][15] ), 
	.D(n3653), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[191][14]  (.Q(\ram[191][14] ), 
	.D(n3652), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[191][13]  (.Q(\ram[191][13] ), 
	.D(n3651), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[191][12]  (.Q(\ram[191][12] ), 
	.D(n3650), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[191][11]  (.Q(\ram[191][11] ), 
	.D(n3649), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[191][10]  (.Q(\ram[191][10] ), 
	.D(n3648), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][9]  (.Q(\ram[191][9] ), 
	.D(n3647), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[191][8]  (.Q(\ram[191][8] ), 
	.D(n3646), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][7]  (.Q(\ram[191][7] ), 
	.D(n3645), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][6]  (.Q(\ram[191][6] ), 
	.D(n3644), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[191][5]  (.Q(\ram[191][5] ), 
	.D(n3643), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[191][4]  (.Q(\ram[191][4] ), 
	.D(n3642), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][3]  (.Q(\ram[191][3] ), 
	.D(n3641), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[191][2]  (.Q(\ram[191][2] ), 
	.D(n3640), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[191][1]  (.Q(\ram[191][1] ), 
	.D(n3639), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][0]  (.Q(\ram[191][0] ), 
	.D(n3638), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[187][15]  (.Q(\ram[187][15] ), 
	.D(n3589), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][14]  (.Q(\ram[187][14] ), 
	.D(n3588), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][13]  (.Q(\ram[187][13] ), 
	.D(n3587), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[187][12]  (.Q(\ram[187][12] ), 
	.D(n3586), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[187][11]  (.Q(\ram[187][11] ), 
	.D(n3585), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[187][10]  (.Q(\ram[187][10] ), 
	.D(n3584), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[187][9]  (.Q(\ram[187][9] ), 
	.D(n3583), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[187][8]  (.Q(\ram[187][8] ), 
	.D(n3582), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[187][7]  (.Q(\ram[187][7] ), 
	.D(n3581), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[187][6]  (.Q(\ram[187][6] ), 
	.D(n3580), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[187][5]  (.Q(\ram[187][5] ), 
	.D(n3579), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[187][4]  (.Q(\ram[187][4] ), 
	.D(n3578), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[187][3]  (.Q(\ram[187][3] ), 
	.D(n3577), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[187][2]  (.Q(\ram[187][2] ), 
	.D(n3576), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][1]  (.Q(\ram[187][1] ), 
	.D(n3575), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][0]  (.Q(\ram[187][0] ), 
	.D(n3574), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[183][15]  (.Q(\ram[183][15] ), 
	.D(n3525), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[183][14]  (.Q(\ram[183][14] ), 
	.D(n3524), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[183][13]  (.Q(\ram[183][13] ), 
	.D(n3523), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[183][12]  (.Q(\ram[183][12] ), 
	.D(n3522), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][11]  (.Q(\ram[183][11] ), 
	.D(n3521), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[183][10]  (.Q(\ram[183][10] ), 
	.D(n3520), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][9]  (.Q(\ram[183][9] ), 
	.D(n3519), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][8]  (.Q(\ram[183][8] ), 
	.D(n3518), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][7]  (.Q(\ram[183][7] ), 
	.D(n3517), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[183][6]  (.Q(\ram[183][6] ), 
	.D(n3516), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[183][5]  (.Q(\ram[183][5] ), 
	.D(n3515), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[183][4]  (.Q(\ram[183][4] ), 
	.D(n3514), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][3]  (.Q(\ram[183][3] ), 
	.D(n3513), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[183][2]  (.Q(\ram[183][2] ), 
	.D(n3512), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][1]  (.Q(\ram[183][1] ), 
	.D(n3511), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][0]  (.Q(\ram[183][0] ), 
	.D(n3510), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[179][15]  (.Q(\ram[179][15] ), 
	.D(n3461), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][14]  (.Q(\ram[179][14] ), 
	.D(n3460), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][13]  (.Q(\ram[179][13] ), 
	.D(n3459), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[179][12]  (.Q(\ram[179][12] ), 
	.D(n3458), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][11]  (.Q(\ram[179][11] ), 
	.D(n3457), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][10]  (.Q(\ram[179][10] ), 
	.D(n3456), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][9]  (.Q(\ram[179][9] ), 
	.D(n3455), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][8]  (.Q(\ram[179][8] ), 
	.D(n3454), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][7]  (.Q(\ram[179][7] ), 
	.D(n3453), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][6]  (.Q(\ram[179][6] ), 
	.D(n3452), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[179][5]  (.Q(\ram[179][5] ), 
	.D(n3451), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[179][4]  (.Q(\ram[179][4] ), 
	.D(n3450), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][3]  (.Q(\ram[179][3] ), 
	.D(n3449), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[179][2]  (.Q(\ram[179][2] ), 
	.D(n3448), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[179][1]  (.Q(\ram[179][1] ), 
	.D(n3447), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][0]  (.Q(\ram[179][0] ), 
	.D(n3446), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[175][15]  (.Q(\ram[175][15] ), 
	.D(n3397), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][14]  (.Q(\ram[175][14] ), 
	.D(n3396), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][13]  (.Q(\ram[175][13] ), 
	.D(n3395), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[175][12]  (.Q(\ram[175][12] ), 
	.D(n3394), 
	.CK(clk));
   QDFFEHD \ram_reg[175][11]  (.Q(\ram[175][11] ), 
	.D(n3393), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][10]  (.Q(\ram[175][10] ), 
	.D(n3392), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][9]  (.Q(\ram[175][9] ), 
	.D(n3391), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][8]  (.Q(\ram[175][8] ), 
	.D(n3390), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][7]  (.Q(\ram[175][7] ), 
	.D(n3389), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][6]  (.Q(\ram[175][6] ), 
	.D(n3388), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][5]  (.Q(\ram[175][5] ), 
	.D(n3387), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][4]  (.Q(\ram[175][4] ), 
	.D(n3386), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[175][3]  (.Q(\ram[175][3] ), 
	.D(n3385), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][2]  (.Q(\ram[175][2] ), 
	.D(n3384), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][1]  (.Q(\ram[175][1] ), 
	.D(n3383), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][0]  (.Q(\ram[175][0] ), 
	.D(n3382), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[171][15]  (.Q(\ram[171][15] ), 
	.D(n3333), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][14]  (.Q(\ram[171][14] ), 
	.D(n3332), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][13]  (.Q(\ram[171][13] ), 
	.D(n3331), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][12]  (.Q(\ram[171][12] ), 
	.D(n3330), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][11]  (.Q(\ram[171][11] ), 
	.D(n3329), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][10]  (.Q(\ram[171][10] ), 
	.D(n3328), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][9]  (.Q(\ram[171][9] ), 
	.D(n3327), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][8]  (.Q(\ram[171][8] ), 
	.D(n3326), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][7]  (.Q(\ram[171][7] ), 
	.D(n3325), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][6]  (.Q(\ram[171][6] ), 
	.D(n3324), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][5]  (.Q(\ram[171][5] ), 
	.D(n3323), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][4]  (.Q(\ram[171][4] ), 
	.D(n3322), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][3]  (.Q(\ram[171][3] ), 
	.D(n3321), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][2]  (.Q(\ram[171][2] ), 
	.D(n3320), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][1]  (.Q(\ram[171][1] ), 
	.D(n3319), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][0]  (.Q(\ram[171][0] ), 
	.D(n3318), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[167][15]  (.Q(\ram[167][15] ), 
	.D(n3269), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[167][14]  (.Q(\ram[167][14] ), 
	.D(n3268), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][13]  (.Q(\ram[167][13] ), 
	.D(n3267), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][12]  (.Q(\ram[167][12] ), 
	.D(n3266), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][11]  (.Q(\ram[167][11] ), 
	.D(n3265), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][10]  (.Q(\ram[167][10] ), 
	.D(n3264), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][9]  (.Q(\ram[167][9] ), 
	.D(n3263), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][8]  (.Q(\ram[167][8] ), 
	.D(n3262), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][7]  (.Q(\ram[167][7] ), 
	.D(n3261), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[167][6]  (.Q(\ram[167][6] ), 
	.D(n3260), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][5]  (.Q(\ram[167][5] ), 
	.D(n3259), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][4]  (.Q(\ram[167][4] ), 
	.D(n3258), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][3]  (.Q(\ram[167][3] ), 
	.D(n3257), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][2]  (.Q(\ram[167][2] ), 
	.D(n3256), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][1]  (.Q(\ram[167][1] ), 
	.D(n3255), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][0]  (.Q(\ram[167][0] ), 
	.D(n3254), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[163][15]  (.Q(\ram[163][15] ), 
	.D(n3205), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][14]  (.Q(\ram[163][14] ), 
	.D(n3204), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][13]  (.Q(\ram[163][13] ), 
	.D(n3203), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][12]  (.Q(\ram[163][12] ), 
	.D(n3202), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][11]  (.Q(\ram[163][11] ), 
	.D(n3201), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][10]  (.Q(\ram[163][10] ), 
	.D(n3200), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][9]  (.Q(\ram[163][9] ), 
	.D(n3199), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][8]  (.Q(\ram[163][8] ), 
	.D(n3198), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][7]  (.Q(\ram[163][7] ), 
	.D(n3197), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[163][6]  (.Q(\ram[163][6] ), 
	.D(n3196), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[163][5]  (.Q(\ram[163][5] ), 
	.D(n3195), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][4]  (.Q(\ram[163][4] ), 
	.D(n3194), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][3]  (.Q(\ram[163][3] ), 
	.D(n3193), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][2]  (.Q(\ram[163][2] ), 
	.D(n3192), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][1]  (.Q(\ram[163][1] ), 
	.D(n3191), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[163][0]  (.Q(\ram[163][0] ), 
	.D(n3190), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[159][15]  (.Q(\ram[159][15] ), 
	.D(n3141), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[159][14]  (.Q(\ram[159][14] ), 
	.D(n3140), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][13]  (.Q(\ram[159][13] ), 
	.D(n3139), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][12]  (.Q(\ram[159][12] ), 
	.D(n3138), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][11]  (.Q(\ram[159][11] ), 
	.D(n3137), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][10]  (.Q(\ram[159][10] ), 
	.D(n3136), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[159][9]  (.Q(\ram[159][9] ), 
	.D(n3135), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[159][8]  (.Q(\ram[159][8] ), 
	.D(n3134), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[159][7]  (.Q(\ram[159][7] ), 
	.D(n3133), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[159][6]  (.Q(\ram[159][6] ), 
	.D(n3132), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[159][5]  (.Q(\ram[159][5] ), 
	.D(n3131), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[159][4]  (.Q(\ram[159][4] ), 
	.D(n3130), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[159][3]  (.Q(\ram[159][3] ), 
	.D(n3129), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[159][2]  (.Q(\ram[159][2] ), 
	.D(n3128), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[159][1]  (.Q(\ram[159][1] ), 
	.D(n3127), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[159][0]  (.Q(\ram[159][0] ), 
	.D(n3126), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[155][15]  (.Q(\ram[155][15] ), 
	.D(n3077), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[155][14]  (.Q(\ram[155][14] ), 
	.D(n3076), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][13]  (.Q(\ram[155][13] ), 
	.D(n3075), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][12]  (.Q(\ram[155][12] ), 
	.D(n3074), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][11]  (.Q(\ram[155][11] ), 
	.D(n3073), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][10]  (.Q(\ram[155][10] ), 
	.D(n3072), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][9]  (.Q(\ram[155][9] ), 
	.D(n3071), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[155][8]  (.Q(\ram[155][8] ), 
	.D(n3070), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[155][7]  (.Q(\ram[155][7] ), 
	.D(n3069), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][6]  (.Q(\ram[155][6] ), 
	.D(n3068), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][5]  (.Q(\ram[155][5] ), 
	.D(n3067), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[155][4]  (.Q(\ram[155][4] ), 
	.D(n3066), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[155][3]  (.Q(\ram[155][3] ), 
	.D(n3065), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][2]  (.Q(\ram[155][2] ), 
	.D(n3064), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][1]  (.Q(\ram[155][1] ), 
	.D(n3063), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][0]  (.Q(\ram[155][0] ), 
	.D(n3062), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[151][15]  (.Q(\ram[151][15] ), 
	.D(n3013), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][14]  (.Q(\ram[151][14] ), 
	.D(n3012), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][13]  (.Q(\ram[151][13] ), 
	.D(n3011), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][12]  (.Q(\ram[151][12] ), 
	.D(n3010), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[151][11]  (.Q(\ram[151][11] ), 
	.D(n3009), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][10]  (.Q(\ram[151][10] ), 
	.D(n3008), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[151][9]  (.Q(\ram[151][9] ), 
	.D(n3007), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[151][8]  (.Q(\ram[151][8] ), 
	.D(n3006), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[151][7]  (.Q(\ram[151][7] ), 
	.D(n3005), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[151][6]  (.Q(\ram[151][6] ), 
	.D(n3004), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[151][5]  (.Q(\ram[151][5] ), 
	.D(n3003), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[151][4]  (.Q(\ram[151][4] ), 
	.D(n3002), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[151][3]  (.Q(\ram[151][3] ), 
	.D(n3001), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[151][2]  (.Q(\ram[151][2] ), 
	.D(n3000), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[151][1]  (.Q(\ram[151][1] ), 
	.D(n2999), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[151][0]  (.Q(\ram[151][0] ), 
	.D(n2998), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[147][15]  (.Q(\ram[147][15] ), 
	.D(n2949), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[147][14]  (.Q(\ram[147][14] ), 
	.D(n2948), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[147][13]  (.Q(\ram[147][13] ), 
	.D(n2947), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[147][12]  (.Q(\ram[147][12] ), 
	.D(n2946), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][11]  (.Q(\ram[147][11] ), 
	.D(n2945), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][10]  (.Q(\ram[147][10] ), 
	.D(n2944), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[147][9]  (.Q(\ram[147][9] ), 
	.D(n2943), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][8]  (.Q(\ram[147][8] ), 
	.D(n2942), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][7]  (.Q(\ram[147][7] ), 
	.D(n2941), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][6]  (.Q(\ram[147][6] ), 
	.D(n2940), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][5]  (.Q(\ram[147][5] ), 
	.D(n2939), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][4]  (.Q(\ram[147][4] ), 
	.D(n2938), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][3]  (.Q(\ram[147][3] ), 
	.D(n2937), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][2]  (.Q(\ram[147][2] ), 
	.D(n2936), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[147][1]  (.Q(\ram[147][1] ), 
	.D(n2935), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][0]  (.Q(\ram[147][0] ), 
	.D(n2934), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[143][15]  (.Q(\ram[143][15] ), 
	.D(n2885), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[143][14]  (.Q(\ram[143][14] ), 
	.D(n2884), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[143][13]  (.Q(\ram[143][13] ), 
	.D(n2883), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[143][12]  (.Q(\ram[143][12] ), 
	.D(n2882), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[143][11]  (.Q(\ram[143][11] ), 
	.D(n2881), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[143][10]  (.Q(\ram[143][10] ), 
	.D(n2880), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[143][9]  (.Q(\ram[143][9] ), 
	.D(n2879), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[143][8]  (.Q(\ram[143][8] ), 
	.D(n2878), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[143][7]  (.Q(\ram[143][7] ), 
	.D(n2877), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[143][6]  (.Q(\ram[143][6] ), 
	.D(n2876), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[143][5]  (.Q(\ram[143][5] ), 
	.D(n2875), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[143][4]  (.Q(\ram[143][4] ), 
	.D(n2874), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[143][3]  (.Q(\ram[143][3] ), 
	.D(n2873), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[143][2]  (.Q(\ram[143][2] ), 
	.D(n2872), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[143][1]  (.Q(\ram[143][1] ), 
	.D(n2871), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[143][0]  (.Q(\ram[143][0] ), 
	.D(n2870), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[139][15]  (.Q(\ram[139][15] ), 
	.D(n2821), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][14]  (.Q(\ram[139][14] ), 
	.D(n2820), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][13]  (.Q(\ram[139][13] ), 
	.D(n2819), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][12]  (.Q(\ram[139][12] ), 
	.D(n2818), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][11]  (.Q(\ram[139][11] ), 
	.D(n2817), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][10]  (.Q(\ram[139][10] ), 
	.D(n2816), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][9]  (.Q(\ram[139][9] ), 
	.D(n2815), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][8]  (.Q(\ram[139][8] ), 
	.D(n2814), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][7]  (.Q(\ram[139][7] ), 
	.D(n2813), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][6]  (.Q(\ram[139][6] ), 
	.D(n2812), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[139][5]  (.Q(\ram[139][5] ), 
	.D(n2811), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[139][4]  (.Q(\ram[139][4] ), 
	.D(n2810), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[139][3]  (.Q(\ram[139][3] ), 
	.D(n2809), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[139][2]  (.Q(\ram[139][2] ), 
	.D(n2808), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][1]  (.Q(\ram[139][1] ), 
	.D(n2807), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[139][0]  (.Q(\ram[139][0] ), 
	.D(n2806), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[135][15]  (.Q(\ram[135][15] ), 
	.D(n2757), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[135][14]  (.Q(\ram[135][14] ), 
	.D(n2756), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[135][13]  (.Q(\ram[135][13] ), 
	.D(n2755), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[135][12]  (.Q(\ram[135][12] ), 
	.D(n2754), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][11]  (.Q(\ram[135][11] ), 
	.D(n2753), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[135][10]  (.Q(\ram[135][10] ), 
	.D(n2752), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][9]  (.Q(\ram[135][9] ), 
	.D(n2751), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[135][8]  (.Q(\ram[135][8] ), 
	.D(n2750), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][7]  (.Q(\ram[135][7] ), 
	.D(n2749), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][6]  (.Q(\ram[135][6] ), 
	.D(n2748), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][5]  (.Q(\ram[135][5] ), 
	.D(n2747), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][4]  (.Q(\ram[135][4] ), 
	.D(n2746), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][3]  (.Q(\ram[135][3] ), 
	.D(n2745), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[135][2]  (.Q(\ram[135][2] ), 
	.D(n2744), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][1]  (.Q(\ram[135][1] ), 
	.D(n2743), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][0]  (.Q(\ram[135][0] ), 
	.D(n2742), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[131][15]  (.Q(\ram[131][15] ), 
	.D(n2693), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][14]  (.Q(\ram[131][14] ), 
	.D(n2692), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][13]  (.Q(\ram[131][13] ), 
	.D(n2691), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][12]  (.Q(\ram[131][12] ), 
	.D(n2690), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[131][11]  (.Q(\ram[131][11] ), 
	.D(n2689), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[131][10]  (.Q(\ram[131][10] ), 
	.D(n2688), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[131][9]  (.Q(\ram[131][9] ), 
	.D(n2687), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][8]  (.Q(\ram[131][8] ), 
	.D(n2686), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[131][7]  (.Q(\ram[131][7] ), 
	.D(n2685), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[131][6]  (.Q(\ram[131][6] ), 
	.D(n2684), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][5]  (.Q(\ram[131][5] ), 
	.D(n2683), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[131][4]  (.Q(\ram[131][4] ), 
	.D(n2682), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][3]  (.Q(\ram[131][3] ), 
	.D(n2681), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][2]  (.Q(\ram[131][2] ), 
	.D(n2680), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[131][1]  (.Q(\ram[131][1] ), 
	.D(n2679), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][0]  (.Q(\ram[131][0] ), 
	.D(n2678), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[127][15]  (.Q(\ram[127][15] ), 
	.D(n2629), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[127][14]  (.Q(\ram[127][14] ), 
	.D(n2628), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[127][13]  (.Q(\ram[127][13] ), 
	.D(n2627), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[127][12]  (.Q(\ram[127][12] ), 
	.D(n2626), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][11]  (.Q(\ram[127][11] ), 
	.D(n2625), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][10]  (.Q(\ram[127][10] ), 
	.D(n2624), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][9]  (.Q(\ram[127][9] ), 
	.D(n2623), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[127][8]  (.Q(\ram[127][8] ), 
	.D(n2622), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][7]  (.Q(\ram[127][7] ), 
	.D(n2621), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][6]  (.Q(\ram[127][6] ), 
	.D(n2620), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[127][5]  (.Q(\ram[127][5] ), 
	.D(n2619), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][4]  (.Q(\ram[127][4] ), 
	.D(n2618), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[127][3]  (.Q(\ram[127][3] ), 
	.D(n2617), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[127][2]  (.Q(\ram[127][2] ), 
	.D(n2616), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][1]  (.Q(\ram[127][1] ), 
	.D(n2615), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[127][0]  (.Q(\ram[127][0] ), 
	.D(n2614), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[123][15]  (.Q(\ram[123][15] ), 
	.D(n2565), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][14]  (.Q(\ram[123][14] ), 
	.D(n2564), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][13]  (.Q(\ram[123][13] ), 
	.D(n2563), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[123][12]  (.Q(\ram[123][12] ), 
	.D(n2562), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][11]  (.Q(\ram[123][11] ), 
	.D(n2561), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[123][10]  (.Q(\ram[123][10] ), 
	.D(n2560), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[123][9]  (.Q(\ram[123][9] ), 
	.D(n2559), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][8]  (.Q(\ram[123][8] ), 
	.D(n2558), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[123][7]  (.Q(\ram[123][7] ), 
	.D(n2557), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[123][6]  (.Q(\ram[123][6] ), 
	.D(n2556), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[123][5]  (.Q(\ram[123][5] ), 
	.D(n2555), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[123][4]  (.Q(\ram[123][4] ), 
	.D(n2554), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[123][3]  (.Q(\ram[123][3] ), 
	.D(n2553), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[123][2]  (.Q(\ram[123][2] ), 
	.D(n2552), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[123][1]  (.Q(\ram[123][1] ), 
	.D(n2551), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[123][0]  (.Q(\ram[123][0] ), 
	.D(n2550), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[119][15]  (.Q(\ram[119][15] ), 
	.D(n2501), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[119][14]  (.Q(\ram[119][14] ), 
	.D(n2500), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][13]  (.Q(\ram[119][13] ), 
	.D(n2499), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[119][12]  (.Q(\ram[119][12] ), 
	.D(n2498), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[119][11]  (.Q(\ram[119][11] ), 
	.D(n2497), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][10]  (.Q(\ram[119][10] ), 
	.D(n2496), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[119][9]  (.Q(\ram[119][9] ), 
	.D(n2495), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][8]  (.Q(\ram[119][8] ), 
	.D(n2494), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][7]  (.Q(\ram[119][7] ), 
	.D(n2493), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][6]  (.Q(\ram[119][6] ), 
	.D(n2492), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][5]  (.Q(\ram[119][5] ), 
	.D(n2491), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[119][4]  (.Q(\ram[119][4] ), 
	.D(n2490), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][3]  (.Q(\ram[119][3] ), 
	.D(n2489), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][2]  (.Q(\ram[119][2] ), 
	.D(n2488), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][1]  (.Q(\ram[119][1] ), 
	.D(n2487), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[119][0]  (.Q(\ram[119][0] ), 
	.D(n2486), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[115][15]  (.Q(\ram[115][15] ), 
	.D(n2437), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[115][14]  (.Q(\ram[115][14] ), 
	.D(n2436), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[115][13]  (.Q(\ram[115][13] ), 
	.D(n2435), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[115][12]  (.Q(\ram[115][12] ), 
	.D(n2434), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][11]  (.Q(\ram[115][11] ), 
	.D(n2433), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][10]  (.Q(\ram[115][10] ), 
	.D(n2432), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[115][9]  (.Q(\ram[115][9] ), 
	.D(n2431), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[115][8]  (.Q(\ram[115][8] ), 
	.D(n2430), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][7]  (.Q(\ram[115][7] ), 
	.D(n2429), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][6]  (.Q(\ram[115][6] ), 
	.D(n2428), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[115][5]  (.Q(\ram[115][5] ), 
	.D(n2427), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[115][4]  (.Q(\ram[115][4] ), 
	.D(n2426), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[115][3]  (.Q(\ram[115][3] ), 
	.D(n2425), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[115][2]  (.Q(\ram[115][2] ), 
	.D(n2424), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[115][1]  (.Q(\ram[115][1] ), 
	.D(n2423), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][0]  (.Q(\ram[115][0] ), 
	.D(n2422), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[111][15]  (.Q(\ram[111][15] ), 
	.D(n2373), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][14]  (.Q(\ram[111][14] ), 
	.D(n2372), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][13]  (.Q(\ram[111][13] ), 
	.D(n2371), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][12]  (.Q(\ram[111][12] ), 
	.D(n2370), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][11]  (.Q(\ram[111][11] ), 
	.D(n2369), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][10]  (.Q(\ram[111][10] ), 
	.D(n2368), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][9]  (.Q(\ram[111][9] ), 
	.D(n2367), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][8]  (.Q(\ram[111][8] ), 
	.D(n2366), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][7]  (.Q(\ram[111][7] ), 
	.D(n2365), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][6]  (.Q(\ram[111][6] ), 
	.D(n2364), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][5]  (.Q(\ram[111][5] ), 
	.D(n2363), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][4]  (.Q(\ram[111][4] ), 
	.D(n2362), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][3]  (.Q(\ram[111][3] ), 
	.D(n2361), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][2]  (.Q(\ram[111][2] ), 
	.D(n2360), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][1]  (.Q(\ram[111][1] ), 
	.D(n2359), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][0]  (.Q(\ram[111][0] ), 
	.D(n2358), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[107][15]  (.Q(\ram[107][15] ), 
	.D(n2309), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][14]  (.Q(\ram[107][14] ), 
	.D(n2308), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[107][13]  (.Q(\ram[107][13] ), 
	.D(n2307), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[107][12]  (.Q(\ram[107][12] ), 
	.D(n2306), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[107][11]  (.Q(\ram[107][11] ), 
	.D(n2305), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[107][10]  (.Q(\ram[107][10] ), 
	.D(n2304), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][9]  (.Q(\ram[107][9] ), 
	.D(n2303), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][8]  (.Q(\ram[107][8] ), 
	.D(n2302), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[107][7]  (.Q(\ram[107][7] ), 
	.D(n2301), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[107][6]  (.Q(\ram[107][6] ), 
	.D(n2300), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][5]  (.Q(\ram[107][5] ), 
	.D(n2299), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[107][4]  (.Q(\ram[107][4] ), 
	.D(n2298), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][3]  (.Q(\ram[107][3] ), 
	.D(n2297), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[107][2]  (.Q(\ram[107][2] ), 
	.D(n2296), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][1]  (.Q(\ram[107][1] ), 
	.D(n2295), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[107][0]  (.Q(\ram[107][0] ), 
	.D(n2294), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[103][15]  (.Q(\ram[103][15] ), 
	.D(n2245), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[103][14]  (.Q(\ram[103][14] ), 
	.D(n2244), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[103][13]  (.Q(\ram[103][13] ), 
	.D(n2243), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][12]  (.Q(\ram[103][12] ), 
	.D(n2242), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][11]  (.Q(\ram[103][11] ), 
	.D(n2241), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][10]  (.Q(\ram[103][10] ), 
	.D(n2240), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][9]  (.Q(\ram[103][9] ), 
	.D(n2239), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][8]  (.Q(\ram[103][8] ), 
	.D(n2238), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][7]  (.Q(\ram[103][7] ), 
	.D(n2237), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[103][6]  (.Q(\ram[103][6] ), 
	.D(n2236), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][5]  (.Q(\ram[103][5] ), 
	.D(n2235), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][4]  (.Q(\ram[103][4] ), 
	.D(n2234), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][3]  (.Q(\ram[103][3] ), 
	.D(n2233), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[103][2]  (.Q(\ram[103][2] ), 
	.D(n2232), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][1]  (.Q(\ram[103][1] ), 
	.D(n2231), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[103][0]  (.Q(\ram[103][0] ), 
	.D(n2230), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[99][15]  (.Q(\ram[99][15] ), 
	.D(n2181), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[99][14]  (.Q(\ram[99][14] ), 
	.D(n2180), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][13]  (.Q(\ram[99][13] ), 
	.D(n2179), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[99][12]  (.Q(\ram[99][12] ), 
	.D(n2178), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[99][11]  (.Q(\ram[99][11] ), 
	.D(n2177), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[99][10]  (.Q(\ram[99][10] ), 
	.D(n2176), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][9]  (.Q(\ram[99][9] ), 
	.D(n2175), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][8]  (.Q(\ram[99][8] ), 
	.D(n2174), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][7]  (.Q(\ram[99][7] ), 
	.D(n2173), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[99][6]  (.Q(\ram[99][6] ), 
	.D(n2172), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][5]  (.Q(\ram[99][5] ), 
	.D(n2171), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][4]  (.Q(\ram[99][4] ), 
	.D(n2170), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][3]  (.Q(\ram[99][3] ), 
	.D(n2169), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[99][2]  (.Q(\ram[99][2] ), 
	.D(n2168), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[99][1]  (.Q(\ram[99][1] ), 
	.D(n2167), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[99][0]  (.Q(\ram[99][0] ), 
	.D(n2166), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[95][15]  (.Q(\ram[95][15] ), 
	.D(n2117), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][14]  (.Q(\ram[95][14] ), 
	.D(n2116), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[95][13]  (.Q(\ram[95][13] ), 
	.D(n2115), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][12]  (.Q(\ram[95][12] ), 
	.D(n2114), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[95][11]  (.Q(\ram[95][11] ), 
	.D(n2113), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[95][10]  (.Q(\ram[95][10] ), 
	.D(n2112), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][9]  (.Q(\ram[95][9] ), 
	.D(n2111), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][8]  (.Q(\ram[95][8] ), 
	.D(n2110), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[95][7]  (.Q(\ram[95][7] ), 
	.D(n2109), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][6]  (.Q(\ram[95][6] ), 
	.D(n2108), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[95][5]  (.Q(\ram[95][5] ), 
	.D(n2107), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[95][4]  (.Q(\ram[95][4] ), 
	.D(n2106), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][3]  (.Q(\ram[95][3] ), 
	.D(n2105), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][2]  (.Q(\ram[95][2] ), 
	.D(n2104), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][1]  (.Q(\ram[95][1] ), 
	.D(n2103), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][0]  (.Q(\ram[95][0] ), 
	.D(n2102), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[91][15]  (.Q(\ram[91][15] ), 
	.D(n2053), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][14]  (.Q(\ram[91][14] ), 
	.D(n2052), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[91][13]  (.Q(\ram[91][13] ), 
	.D(n2051), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][12]  (.Q(\ram[91][12] ), 
	.D(n2050), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][11]  (.Q(\ram[91][11] ), 
	.D(n2049), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][10]  (.Q(\ram[91][10] ), 
	.D(n2048), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][9]  (.Q(\ram[91][9] ), 
	.D(n2047), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][8]  (.Q(\ram[91][8] ), 
	.D(n2046), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][7]  (.Q(\ram[91][7] ), 
	.D(n2045), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][6]  (.Q(\ram[91][6] ), 
	.D(n2044), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][5]  (.Q(\ram[91][5] ), 
	.D(n2043), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][4]  (.Q(\ram[91][4] ), 
	.D(n2042), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][3]  (.Q(\ram[91][3] ), 
	.D(n2041), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][2]  (.Q(\ram[91][2] ), 
	.D(n2040), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][1]  (.Q(\ram[91][1] ), 
	.D(n2039), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][0]  (.Q(\ram[91][0] ), 
	.D(n2038), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[87][15]  (.Q(\ram[87][15] ), 
	.D(n1989), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][14]  (.Q(\ram[87][14] ), 
	.D(n1988), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][13]  (.Q(\ram[87][13] ), 
	.D(n1987), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[87][12]  (.Q(\ram[87][12] ), 
	.D(n1986), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[87][11]  (.Q(\ram[87][11] ), 
	.D(n1985), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][10]  (.Q(\ram[87][10] ), 
	.D(n1984), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][9]  (.Q(\ram[87][9] ), 
	.D(n1983), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][8]  (.Q(\ram[87][8] ), 
	.D(n1982), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][7]  (.Q(\ram[87][7] ), 
	.D(n1981), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][6]  (.Q(\ram[87][6] ), 
	.D(n1980), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][5]  (.Q(\ram[87][5] ), 
	.D(n1979), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][4]  (.Q(\ram[87][4] ), 
	.D(n1978), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][3]  (.Q(\ram[87][3] ), 
	.D(n1977), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][2]  (.Q(\ram[87][2] ), 
	.D(n1976), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][1]  (.Q(\ram[87][1] ), 
	.D(n1975), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[87][0]  (.Q(\ram[87][0] ), 
	.D(n1974), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[83][15]  (.Q(\ram[83][15] ), 
	.D(n1925), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][14]  (.Q(\ram[83][14] ), 
	.D(n1924), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][13]  (.Q(\ram[83][13] ), 
	.D(n1923), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][12]  (.Q(\ram[83][12] ), 
	.D(n1922), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][11]  (.Q(\ram[83][11] ), 
	.D(n1921), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[83][10]  (.Q(\ram[83][10] ), 
	.D(n1920), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][9]  (.Q(\ram[83][9] ), 
	.D(n1919), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][8]  (.Q(\ram[83][8] ), 
	.D(n1918), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][7]  (.Q(\ram[83][7] ), 
	.D(n1917), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][6]  (.Q(\ram[83][6] ), 
	.D(n1916), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][5]  (.Q(\ram[83][5] ), 
	.D(n1915), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[83][4]  (.Q(\ram[83][4] ), 
	.D(n1914), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[83][3]  (.Q(\ram[83][3] ), 
	.D(n1913), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][2]  (.Q(\ram[83][2] ), 
	.D(n1912), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[83][1]  (.Q(\ram[83][1] ), 
	.D(n1911), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[83][0]  (.Q(\ram[83][0] ), 
	.D(n1910), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[79][15]  (.Q(\ram[79][15] ), 
	.D(n1861), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][14]  (.Q(\ram[79][14] ), 
	.D(n1860), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][13]  (.Q(\ram[79][13] ), 
	.D(n1859), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][12]  (.Q(\ram[79][12] ), 
	.D(n1858), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][11]  (.Q(\ram[79][11] ), 
	.D(n1857), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][10]  (.Q(\ram[79][10] ), 
	.D(n1856), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[79][9]  (.Q(\ram[79][9] ), 
	.D(n1855), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][8]  (.Q(\ram[79][8] ), 
	.D(n1854), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][7]  (.Q(\ram[79][7] ), 
	.D(n1853), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[79][6]  (.Q(\ram[79][6] ), 
	.D(n1852), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][5]  (.Q(\ram[79][5] ), 
	.D(n1851), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][4]  (.Q(\ram[79][4] ), 
	.D(n1850), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][3]  (.Q(\ram[79][3] ), 
	.D(n1849), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[79][2]  (.Q(\ram[79][2] ), 
	.D(n1848), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[79][1]  (.Q(\ram[79][1] ), 
	.D(n1847), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[79][0]  (.Q(\ram[79][0] ), 
	.D(n1846), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[75][15]  (.Q(\ram[75][15] ), 
	.D(n1797), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][14]  (.Q(\ram[75][14] ), 
	.D(n1796), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][13]  (.Q(\ram[75][13] ), 
	.D(n1795), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][12]  (.Q(\ram[75][12] ), 
	.D(n1794), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][11]  (.Q(\ram[75][11] ), 
	.D(n1793), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][10]  (.Q(\ram[75][10] ), 
	.D(n1792), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][9]  (.Q(\ram[75][9] ), 
	.D(n1791), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][8]  (.Q(\ram[75][8] ), 
	.D(n1790), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[75][7]  (.Q(\ram[75][7] ), 
	.D(n1789), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][6]  (.Q(\ram[75][6] ), 
	.D(n1788), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][5]  (.Q(\ram[75][5] ), 
	.D(n1787), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][4]  (.Q(\ram[75][4] ), 
	.D(n1786), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][3]  (.Q(\ram[75][3] ), 
	.D(n1785), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[75][2]  (.Q(\ram[75][2] ), 
	.D(n1784), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][1]  (.Q(\ram[75][1] ), 
	.D(n1783), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][0]  (.Q(\ram[75][0] ), 
	.D(n1782), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[71][15]  (.Q(\ram[71][15] ), 
	.D(n1733), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][14]  (.Q(\ram[71][14] ), 
	.D(n1732), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][13]  (.Q(\ram[71][13] ), 
	.D(n1731), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][12]  (.Q(\ram[71][12] ), 
	.D(n1730), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][11]  (.Q(\ram[71][11] ), 
	.D(n1729), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][10]  (.Q(\ram[71][10] ), 
	.D(n1728), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][9]  (.Q(\ram[71][9] ), 
	.D(n1727), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][8]  (.Q(\ram[71][8] ), 
	.D(n1726), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][7]  (.Q(\ram[71][7] ), 
	.D(n1725), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][6]  (.Q(\ram[71][6] ), 
	.D(n1724), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][5]  (.Q(\ram[71][5] ), 
	.D(n1723), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][4]  (.Q(\ram[71][4] ), 
	.D(n1722), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][3]  (.Q(\ram[71][3] ), 
	.D(n1721), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[71][2]  (.Q(\ram[71][2] ), 
	.D(n1720), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][1]  (.Q(\ram[71][1] ), 
	.D(n1719), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[71][0]  (.Q(\ram[71][0] ), 
	.D(n1718), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[67][15]  (.Q(\ram[67][15] ), 
	.D(n1669), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[67][14]  (.Q(\ram[67][14] ), 
	.D(n1668), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[67][13]  (.Q(\ram[67][13] ), 
	.D(n1667), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[67][12]  (.Q(\ram[67][12] ), 
	.D(n1666), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[67][11]  (.Q(\ram[67][11] ), 
	.D(n1665), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][10]  (.Q(\ram[67][10] ), 
	.D(n1664), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[67][9]  (.Q(\ram[67][9] ), 
	.D(n1663), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[67][8]  (.Q(\ram[67][8] ), 
	.D(n1662), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][7]  (.Q(\ram[67][7] ), 
	.D(n1661), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[67][6]  (.Q(\ram[67][6] ), 
	.D(n1660), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[67][5]  (.Q(\ram[67][5] ), 
	.D(n1659), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][4]  (.Q(\ram[67][4] ), 
	.D(n1658), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][3]  (.Q(\ram[67][3] ), 
	.D(n1657), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][2]  (.Q(\ram[67][2] ), 
	.D(n1656), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[67][1]  (.Q(\ram[67][1] ), 
	.D(n1655), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[67][0]  (.Q(\ram[67][0] ), 
	.D(n1654), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[63][15]  (.Q(\ram[63][15] ), 
	.D(n1605), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][14]  (.Q(\ram[63][14] ), 
	.D(n1604), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][13]  (.Q(\ram[63][13] ), 
	.D(n1603), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][12]  (.Q(\ram[63][12] ), 
	.D(n1602), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[63][11]  (.Q(\ram[63][11] ), 
	.D(n1601), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[63][10]  (.Q(\ram[63][10] ), 
	.D(n1600), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][9]  (.Q(\ram[63][9] ), 
	.D(n1599), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[63][8]  (.Q(\ram[63][8] ), 
	.D(n1598), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][7]  (.Q(\ram[63][7] ), 
	.D(n1597), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][6]  (.Q(\ram[63][6] ), 
	.D(n1596), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][5]  (.Q(\ram[63][5] ), 
	.D(n1595), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][4]  (.Q(\ram[63][4] ), 
	.D(n1594), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[63][3]  (.Q(\ram[63][3] ), 
	.D(n1593), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][2]  (.Q(\ram[63][2] ), 
	.D(n1592), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[63][1]  (.Q(\ram[63][1] ), 
	.D(n1591), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[63][0]  (.Q(\ram[63][0] ), 
	.D(n1590), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[59][15]  (.Q(\ram[59][15] ), 
	.D(n1541), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][14]  (.Q(\ram[59][14] ), 
	.D(n1540), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][13]  (.Q(\ram[59][13] ), 
	.D(n1539), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][12]  (.Q(\ram[59][12] ), 
	.D(n1538), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[59][11]  (.Q(\ram[59][11] ), 
	.D(n1537), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][10]  (.Q(\ram[59][10] ), 
	.D(n1536), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][9]  (.Q(\ram[59][9] ), 
	.D(n1535), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][8]  (.Q(\ram[59][8] ), 
	.D(n1534), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][7]  (.Q(\ram[59][7] ), 
	.D(n1533), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][6]  (.Q(\ram[59][6] ), 
	.D(n1532), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][5]  (.Q(\ram[59][5] ), 
	.D(n1531), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][4]  (.Q(\ram[59][4] ), 
	.D(n1530), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[59][3]  (.Q(\ram[59][3] ), 
	.D(n1529), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][2]  (.Q(\ram[59][2] ), 
	.D(n1528), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][1]  (.Q(\ram[59][1] ), 
	.D(n1527), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[59][0]  (.Q(\ram[59][0] ), 
	.D(n1526), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[55][15]  (.Q(\ram[55][15] ), 
	.D(n1477), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][14]  (.Q(\ram[55][14] ), 
	.D(n1476), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][13]  (.Q(\ram[55][13] ), 
	.D(n1475), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][12]  (.Q(\ram[55][12] ), 
	.D(n1474), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[55][11]  (.Q(\ram[55][11] ), 
	.D(n1473), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][10]  (.Q(\ram[55][10] ), 
	.D(n1472), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][9]  (.Q(\ram[55][9] ), 
	.D(n1471), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][8]  (.Q(\ram[55][8] ), 
	.D(n1470), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][7]  (.Q(\ram[55][7] ), 
	.D(n1469), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][6]  (.Q(\ram[55][6] ), 
	.D(n1468), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][5]  (.Q(\ram[55][5] ), 
	.D(n1467), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][4]  (.Q(\ram[55][4] ), 
	.D(n1466), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][3]  (.Q(\ram[55][3] ), 
	.D(n1465), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][2]  (.Q(\ram[55][2] ), 
	.D(n1464), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][1]  (.Q(\ram[55][1] ), 
	.D(n1463), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][0]  (.Q(\ram[55][0] ), 
	.D(n1462), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[51][15]  (.Q(\ram[51][15] ), 
	.D(n1413), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[51][14]  (.Q(\ram[51][14] ), 
	.D(n1412), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][13]  (.Q(\ram[51][13] ), 
	.D(n1411), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][12]  (.Q(\ram[51][12] ), 
	.D(n1410), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[51][11]  (.Q(\ram[51][11] ), 
	.D(n1409), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][10]  (.Q(\ram[51][10] ), 
	.D(n1408), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][9]  (.Q(\ram[51][9] ), 
	.D(n1407), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[51][8]  (.Q(\ram[51][8] ), 
	.D(n1406), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][7]  (.Q(\ram[51][7] ), 
	.D(n1405), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[51][6]  (.Q(\ram[51][6] ), 
	.D(n1404), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[51][5]  (.Q(\ram[51][5] ), 
	.D(n1403), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][4]  (.Q(\ram[51][4] ), 
	.D(n1402), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][3]  (.Q(\ram[51][3] ), 
	.D(n1401), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][2]  (.Q(\ram[51][2] ), 
	.D(n1400), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[51][1]  (.Q(\ram[51][1] ), 
	.D(n1399), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[51][0]  (.Q(\ram[51][0] ), 
	.D(n1398), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[47][15]  (.Q(\ram[47][15] ), 
	.D(n1349), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[47][14]  (.Q(\ram[47][14] ), 
	.D(n1348), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][13]  (.Q(\ram[47][13] ), 
	.D(n1347), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[47][12]  (.Q(\ram[47][12] ), 
	.D(n1346), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][11]  (.Q(\ram[47][11] ), 
	.D(n1345), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][10]  (.Q(\ram[47][10] ), 
	.D(n1344), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][9]  (.Q(\ram[47][9] ), 
	.D(n1343), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[47][8]  (.Q(\ram[47][8] ), 
	.D(n1342), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[47][7]  (.Q(\ram[47][7] ), 
	.D(n1341), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][6]  (.Q(\ram[47][6] ), 
	.D(n1340), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][5]  (.Q(\ram[47][5] ), 
	.D(n1339), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][4]  (.Q(\ram[47][4] ), 
	.D(n1338), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][3]  (.Q(\ram[47][3] ), 
	.D(n1337), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][2]  (.Q(\ram[47][2] ), 
	.D(n1336), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][1]  (.Q(\ram[47][1] ), 
	.D(n1335), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][0]  (.Q(\ram[47][0] ), 
	.D(n1334), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[43][15]  (.Q(\ram[43][15] ), 
	.D(n1285), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][14]  (.Q(\ram[43][14] ), 
	.D(n1284), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[43][13]  (.Q(\ram[43][13] ), 
	.D(n1283), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[43][12]  (.Q(\ram[43][12] ), 
	.D(n1282), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[43][11]  (.Q(\ram[43][11] ), 
	.D(n1281), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[43][10]  (.Q(\ram[43][10] ), 
	.D(n1280), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][9]  (.Q(\ram[43][9] ), 
	.D(n1279), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][8]  (.Q(\ram[43][8] ), 
	.D(n1278), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][7]  (.Q(\ram[43][7] ), 
	.D(n1277), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[43][6]  (.Q(\ram[43][6] ), 
	.D(n1276), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[43][5]  (.Q(\ram[43][5] ), 
	.D(n1275), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[43][4]  (.Q(\ram[43][4] ), 
	.D(n1274), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[43][3]  (.Q(\ram[43][3] ), 
	.D(n1273), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[43][2]  (.Q(\ram[43][2] ), 
	.D(n1272), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[43][1]  (.Q(\ram[43][1] ), 
	.D(n1271), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[43][0]  (.Q(\ram[43][0] ), 
	.D(n1270), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[39][15]  (.Q(\ram[39][15] ), 
	.D(n1221), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][14]  (.Q(\ram[39][14] ), 
	.D(n1220), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[39][13]  (.Q(\ram[39][13] ), 
	.D(n1219), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[39][12]  (.Q(\ram[39][12] ), 
	.D(n1218), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[39][11]  (.Q(\ram[39][11] ), 
	.D(n1217), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[39][10]  (.Q(\ram[39][10] ), 
	.D(n1216), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][9]  (.Q(\ram[39][9] ), 
	.D(n1215), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][8]  (.Q(\ram[39][8] ), 
	.D(n1214), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[39][7]  (.Q(\ram[39][7] ), 
	.D(n1213), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][6]  (.Q(\ram[39][6] ), 
	.D(n1212), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[39][5]  (.Q(\ram[39][5] ), 
	.D(n1211), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[39][4]  (.Q(\ram[39][4] ), 
	.D(n1210), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[39][3]  (.Q(\ram[39][3] ), 
	.D(n1209), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[39][2]  (.Q(\ram[39][2] ), 
	.D(n1208), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[39][1]  (.Q(\ram[39][1] ), 
	.D(n1207), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[39][0]  (.Q(\ram[39][0] ), 
	.D(n1206), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[35][15]  (.Q(\ram[35][15] ), 
	.D(n1157), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[35][14]  (.Q(\ram[35][14] ), 
	.D(n1156), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][13]  (.Q(\ram[35][13] ), 
	.D(n1155), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][12]  (.Q(\ram[35][12] ), 
	.D(n1154), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][11]  (.Q(\ram[35][11] ), 
	.D(n1153), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][10]  (.Q(\ram[35][10] ), 
	.D(n1152), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][9]  (.Q(\ram[35][9] ), 
	.D(n1151), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[35][8]  (.Q(\ram[35][8] ), 
	.D(n1150), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][7]  (.Q(\ram[35][7] ), 
	.D(n1149), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[35][6]  (.Q(\ram[35][6] ), 
	.D(n1148), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][5]  (.Q(\ram[35][5] ), 
	.D(n1147), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][4]  (.Q(\ram[35][4] ), 
	.D(n1146), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][3]  (.Q(\ram[35][3] ), 
	.D(n1145), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][2]  (.Q(\ram[35][2] ), 
	.D(n1144), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][1]  (.Q(\ram[35][1] ), 
	.D(n1143), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][0]  (.Q(\ram[35][0] ), 
	.D(n1142), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[31][15]  (.Q(\ram[31][15] ), 
	.D(n1093), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[31][14]  (.Q(\ram[31][14] ), 
	.D(n1092), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][13]  (.Q(\ram[31][13] ), 
	.D(n1091), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[31][12]  (.Q(\ram[31][12] ), 
	.D(n1090), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[31][11]  (.Q(\ram[31][11] ), 
	.D(n1089), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][10]  (.Q(\ram[31][10] ), 
	.D(n1088), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[31][9]  (.Q(\ram[31][9] ), 
	.D(n1087), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][8]  (.Q(\ram[31][8] ), 
	.D(n1086), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][7]  (.Q(\ram[31][7] ), 
	.D(n1085), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][6]  (.Q(\ram[31][6] ), 
	.D(n1084), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][5]  (.Q(\ram[31][5] ), 
	.D(n1083), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][4]  (.Q(\ram[31][4] ), 
	.D(n1082), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[31][3]  (.Q(\ram[31][3] ), 
	.D(n1081), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][2]  (.Q(\ram[31][2] ), 
	.D(n1080), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[31][1]  (.Q(\ram[31][1] ), 
	.D(n1079), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][0]  (.Q(\ram[31][0] ), 
	.D(n1078), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[27][15]  (.Q(\ram[27][15] ), 
	.D(n1029), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[27][14]  (.Q(\ram[27][14] ), 
	.D(n1028), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][13]  (.Q(\ram[27][13] ), 
	.D(n1027), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[27][12]  (.Q(\ram[27][12] ), 
	.D(n1026), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[27][11]  (.Q(\ram[27][11] ), 
	.D(n1025), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][10]  (.Q(\ram[27][10] ), 
	.D(n1024), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[27][9]  (.Q(\ram[27][9] ), 
	.D(n1023), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][8]  (.Q(\ram[27][8] ), 
	.D(n1022), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][7]  (.Q(\ram[27][7] ), 
	.D(n1021), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[27][6]  (.Q(\ram[27][6] ), 
	.D(n1020), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][5]  (.Q(\ram[27][5] ), 
	.D(n1019), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[27][4]  (.Q(\ram[27][4] ), 
	.D(n1018), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[27][3]  (.Q(\ram[27][3] ), 
	.D(n1017), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[27][2]  (.Q(\ram[27][2] ), 
	.D(n1016), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[27][1]  (.Q(\ram[27][1] ), 
	.D(n1015), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][0]  (.Q(\ram[27][0] ), 
	.D(n1014), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[23][15]  (.Q(\ram[23][15] ), 
	.D(n965), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][14]  (.Q(\ram[23][14] ), 
	.D(n964), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][13]  (.Q(\ram[23][13] ), 
	.D(n963), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[23][12]  (.Q(\ram[23][12] ), 
	.D(n962), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][11]  (.Q(\ram[23][11] ), 
	.D(n961), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[23][10]  (.Q(\ram[23][10] ), 
	.D(n960), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[23][9]  (.Q(\ram[23][9] ), 
	.D(n959), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][8]  (.Q(\ram[23][8] ), 
	.D(n958), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[23][7]  (.Q(\ram[23][7] ), 
	.D(n957), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][6]  (.Q(\ram[23][6] ), 
	.D(n956), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[23][5]  (.Q(\ram[23][5] ), 
	.D(n955), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[23][4]  (.Q(\ram[23][4] ), 
	.D(n954), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][3]  (.Q(\ram[23][3] ), 
	.D(n953), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[23][2]  (.Q(\ram[23][2] ), 
	.D(n952), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][1]  (.Q(\ram[23][1] ), 
	.D(n951), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][0]  (.Q(\ram[23][0] ), 
	.D(n950), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[19][15]  (.Q(\ram[19][15] ), 
	.D(n901), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[19][14]  (.Q(\ram[19][14] ), 
	.D(n900), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][13]  (.Q(\ram[19][13] ), 
	.D(n899), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[19][12]  (.Q(\ram[19][12] ), 
	.D(n898), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[19][11]  (.Q(\ram[19][11] ), 
	.D(n897), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][10]  (.Q(\ram[19][10] ), 
	.D(n896), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[19][9]  (.Q(\ram[19][9] ), 
	.D(n895), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][8]  (.Q(\ram[19][8] ), 
	.D(n894), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[19][7]  (.Q(\ram[19][7] ), 
	.D(n893), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][6]  (.Q(\ram[19][6] ), 
	.D(n892), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[19][5]  (.Q(\ram[19][5] ), 
	.D(n891), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[19][4]  (.Q(\ram[19][4] ), 
	.D(n890), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][3]  (.Q(\ram[19][3] ), 
	.D(n889), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[19][2]  (.Q(\ram[19][2] ), 
	.D(n888), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[19][1]  (.Q(\ram[19][1] ), 
	.D(n887), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[19][0]  (.Q(\ram[19][0] ), 
	.D(n886), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[15][15]  (.Q(\ram[15][15] ), 
	.D(n837), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][14]  (.Q(\ram[15][14] ), 
	.D(n836), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[15][13]  (.Q(\ram[15][13] ), 
	.D(n835), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][12]  (.Q(\ram[15][12] ), 
	.D(n834), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[15][11]  (.Q(\ram[15][11] ), 
	.D(n833), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[15][10]  (.Q(\ram[15][10] ), 
	.D(n832), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[15][9]  (.Q(\ram[15][9] ), 
	.D(n831), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][8]  (.Q(\ram[15][8] ), 
	.D(n830), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[15][7]  (.Q(\ram[15][7] ), 
	.D(n829), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[15][6]  (.Q(\ram[15][6] ), 
	.D(n828), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][5]  (.Q(\ram[15][5] ), 
	.D(n827), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[15][4]  (.Q(\ram[15][4] ), 
	.D(n826), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[15][3]  (.Q(\ram[15][3] ), 
	.D(n825), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[15][2]  (.Q(\ram[15][2] ), 
	.D(n824), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[15][1]  (.Q(\ram[15][1] ), 
	.D(n823), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[15][0]  (.Q(\ram[15][0] ), 
	.D(n822), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][15]  (.Q(\ram[11][15] ), 
	.D(n773), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[11][14]  (.Q(\ram[11][14] ), 
	.D(n772), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[11][13]  (.Q(\ram[11][13] ), 
	.D(n771), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[11][12]  (.Q(\ram[11][12] ), 
	.D(n770), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][11]  (.Q(\ram[11][11] ), 
	.D(n769), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][10]  (.Q(\ram[11][10] ), 
	.D(n768), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[11][9]  (.Q(\ram[11][9] ), 
	.D(n767), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][8]  (.Q(\ram[11][8] ), 
	.D(n766), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[11][7]  (.Q(\ram[11][7] ), 
	.D(n765), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[11][6]  (.Q(\ram[11][6] ), 
	.D(n764), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[11][5]  (.Q(\ram[11][5] ), 
	.D(n763), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][4]  (.Q(\ram[11][4] ), 
	.D(n762), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][3]  (.Q(\ram[11][3] ), 
	.D(n761), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][2]  (.Q(\ram[11][2] ), 
	.D(n760), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[11][1]  (.Q(\ram[11][1] ), 
	.D(n759), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][0]  (.Q(\ram[11][0] ), 
	.D(n758), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[7][15]  (.Q(\ram[7][15] ), 
	.D(n709), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][14]  (.Q(\ram[7][14] ), 
	.D(n708), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][13]  (.Q(\ram[7][13] ), 
	.D(n707), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[7][12]  (.Q(\ram[7][12] ), 
	.D(n706), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[7][11]  (.Q(\ram[7][11] ), 
	.D(n705), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][10]  (.Q(\ram[7][10] ), 
	.D(n704), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][9]  (.Q(\ram[7][9] ), 
	.D(n703), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[7][8]  (.Q(\ram[7][8] ), 
	.D(n702), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[7][7]  (.Q(\ram[7][7] ), 
	.D(n701), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][6]  (.Q(\ram[7][6] ), 
	.D(n700), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][5]  (.Q(\ram[7][5] ), 
	.D(n699), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[7][4]  (.Q(\ram[7][4] ), 
	.D(n698), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][3]  (.Q(\ram[7][3] ), 
	.D(n697), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[7][2]  (.Q(\ram[7][2] ), 
	.D(n696), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][1]  (.Q(\ram[7][1] ), 
	.D(n695), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[7][0]  (.Q(\ram[7][0] ), 
	.D(n694), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[3][15]  (.Q(\ram[3][15] ), 
	.D(n645), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][14]  (.Q(\ram[3][14] ), 
	.D(n644), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][13]  (.Q(\ram[3][13] ), 
	.D(n643), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][12]  (.Q(\ram[3][12] ), 
	.D(n642), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][11]  (.Q(\ram[3][11] ), 
	.D(n641), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[3][10]  (.Q(\ram[3][10] ), 
	.D(n640), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[3][9]  (.Q(\ram[3][9] ), 
	.D(n639), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[3][8]  (.Q(\ram[3][8] ), 
	.D(n638), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][7]  (.Q(\ram[3][7] ), 
	.D(n637), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][6]  (.Q(\ram[3][6] ), 
	.D(n636), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[3][5]  (.Q(\ram[3][5] ), 
	.D(n635), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[3][4]  (.Q(\ram[3][4] ), 
	.D(n634), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][3]  (.Q(\ram[3][3] ), 
	.D(n633), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[3][2]  (.Q(\ram[3][2] ), 
	.D(n632), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][1]  (.Q(\ram[3][1] ), 
	.D(n631), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][0]  (.Q(\ram[3][0] ), 
	.D(n630), 
	.CK(clk_m__L3_N131));
   AN2EHD U2 (.O(n1), 
	.I2(n545), 
	.I1(n544));
   AN2EHD U3 (.O(n2), 
	.I2(n544), 
	.I1(n548));
   AN2HHD U4 (.O(n3), 
	.I2(n545), 
	.I1(n557));
   AN2HHD U5 (.O(n4), 
	.I2(n548), 
	.I1(n557));
   AN2HHD U6 (.O(n5), 
	.I2(n551), 
	.I1(n557));
   AN2HHD U7 (.O(n7), 
	.I2(n554), 
	.I1(n557));
   AN2HHD U8 (.O(n24), 
	.I2(n545), 
	.I1(n566));
   AN2HHD U9 (.O(n25), 
	.I2(n545), 
	.I1(n575));
   AN2EHD U10 (.O(n26), 
	.I2(n544), 
	.I1(n551));
   AN2EHD U11 (.O(n28), 
	.I2(n544), 
	.I1(n554));
   AN2HHD U12 (.O(n29), 
	.I2(n548), 
	.I1(n566));
   AN2EHD U13 (.O(n31), 
	.I2(n548), 
	.I1(n575));
   AN2HHD U14 (.O(n32), 
	.I2(n551), 
	.I1(n566));
   AN2HHD U15 (.O(n34), 
	.I2(n554), 
	.I1(n566));
   AN2EHD U16 (.O(n35), 
	.I2(n551), 
	.I1(n575));
   AN2HHD U17 (.O(n37), 
	.I2(n554), 
	.I1(n575));
   AN2EHD U18 (.O(n38), 
	.I2(n72), 
	.I1(n208));
   AN2EHD U19 (.O(n40), 
	.I2(n106), 
	.I1(n208));
   AN2EHD U20 (.O(n41), 
	.I2(n140), 
	.I1(n208));
   AN2EHD U21 (.O(n43), 
	.I2(n174), 
	.I1(n208));
   AN2EHD U22 (.O(n44), 
	.I2(n72), 
	.I1(n341));
   AN2EHD U23 (.O(n46), 
	.I2(n72), 
	.I1(n474));
   AN2EHD U24 (.O(n47), 
	.I2(n106), 
	.I1(n341));
   AN2EHD U25 (.O(n49), 
	.I2(n106), 
	.I1(n474));
   AN2EHD U26 (.O(n50), 
	.I2(n140), 
	.I1(n341));
   AN2EHD U27 (.O(n52), 
	.I2(n174), 
	.I1(n341));
   AN2EHD U28 (.O(n53), 
	.I2(n140), 
	.I1(n474));
   AN2EHD U29 (.O(n55), 
	.I2(n174), 
	.I1(n474));
   AN2EHD U30 (.O(n56), 
	.I2(n1), 
	.I1(n38));
   AN2EHD U31 (.O(n58), 
	.I2(n2), 
	.I1(n38));
   AN2EHD U32 (.O(n59), 
	.I2(n26), 
	.I1(n38));
   AN2EHD U33 (.O(n61), 
	.I2(n28), 
	.I1(n38));
   AN2EHD U34 (.O(n62), 
	.I2(n3), 
	.I1(n38));
   AN2EHD U35 (.O(n64), 
	.I2(n4), 
	.I1(n38));
   AN2EHD U36 (.O(n65), 
	.I2(n5), 
	.I1(n38));
   AN2EHD U37 (.O(n67), 
	.I2(n7), 
	.I1(n38));
   AN2EHD U38 (.O(n68), 
	.I2(n24), 
	.I1(n38));
   AN2EHD U39 (.O(n70), 
	.I2(n29), 
	.I1(n38));
   AN2EHD U40 (.O(n73), 
	.I2(n32), 
	.I1(n38));
   AN2EHD U41 (.O(n75), 
	.I2(n34), 
	.I1(n38));
   AN2EHD U42 (.O(n76), 
	.I2(n25), 
	.I1(n38));
   AN2EHD U43 (.O(n78), 
	.I2(n31), 
	.I1(n38));
   AN2EHD U44 (.O(n80), 
	.I2(n35), 
	.I1(n38));
   AN2EHD U45 (.O(n82), 
	.I2(n37), 
	.I1(n38));
   AN2EHD U46 (.O(n84), 
	.I2(n1), 
	.I1(n40));
   AN2EHD U47 (.O(n86), 
	.I2(n2), 
	.I1(n40));
   AN2EHD U48 (.O(n88), 
	.I2(n26), 
	.I1(n40));
   AN2EHD U49 (.O(n90), 
	.I2(n28), 
	.I1(n40));
   AN2EHD U50 (.O(n92), 
	.I2(n3), 
	.I1(n40));
   AN2EHD U51 (.O(n94), 
	.I2(n4), 
	.I1(n40));
   AN2EHD U52 (.O(n96), 
	.I2(n5), 
	.I1(n40));
   AN2EHD U53 (.O(n98), 
	.I2(n7), 
	.I1(n40));
   AN2EHD U54 (.O(n100), 
	.I2(n24), 
	.I1(n40));
   AN2EHD U55 (.O(n102), 
	.I2(n29), 
	.I1(n40));
   AN2EHD U56 (.O(n104), 
	.I2(n32), 
	.I1(n40));
   AN2EHD U57 (.O(n107), 
	.I2(n34), 
	.I1(n40));
   AN2EHD U58 (.O(n109), 
	.I2(n25), 
	.I1(n40));
   AN2EHD U59 (.O(n110), 
	.I2(n31), 
	.I1(n40));
   AN2EHD U60 (.O(n112), 
	.I2(n35), 
	.I1(n40));
   AN2EHD U61 (.O(n114), 
	.I2(n37), 
	.I1(n40));
   AN2EHD U62 (.O(n116), 
	.I2(n1), 
	.I1(n41));
   AN2EHD U63 (.O(n118), 
	.I2(n2), 
	.I1(n41));
   AN2EHD U64 (.O(n120), 
	.I2(n26), 
	.I1(n41));
   AN2EHD U65 (.O(n122), 
	.I2(n28), 
	.I1(n41));
   AN2EHD U66 (.O(n124), 
	.I2(n3), 
	.I1(n41));
   AN2EHD U67 (.O(n126), 
	.I2(n4), 
	.I1(n41));
   AN2EHD U68 (.O(n128), 
	.I2(n5), 
	.I1(n41));
   AN2EHD U69 (.O(n130), 
	.I2(n7), 
	.I1(n41));
   AN2EHD U70 (.O(n132), 
	.I2(n24), 
	.I1(n41));
   AN2EHD U71 (.O(n134), 
	.I2(n29), 
	.I1(n41));
   AN2EHD U72 (.O(n136), 
	.I2(n32), 
	.I1(n41));
   AN2EHD U73 (.O(n138), 
	.I2(n34), 
	.I1(n41));
   AN2EHD U74 (.O(n141), 
	.I2(n25), 
	.I1(n41));
   AN2EHD U75 (.O(n143), 
	.I2(n31), 
	.I1(n41));
   AN2EHD U76 (.O(n144), 
	.I2(n35), 
	.I1(n41));
   AN2EHD U77 (.O(n146), 
	.I2(n37), 
	.I1(n41));
   AN2EHD U78 (.O(n148), 
	.I2(n1), 
	.I1(n43));
   AN2EHD U79 (.O(n150), 
	.I2(n2), 
	.I1(n43));
   AN2EHD U80 (.O(n152), 
	.I2(n26), 
	.I1(n43));
   AN2EHD U81 (.O(n154), 
	.I2(n28), 
	.I1(n43));
   AN2EHD U82 (.O(n156), 
	.I2(n3), 
	.I1(n43));
   AN2EHD U83 (.O(n158), 
	.I2(n4), 
	.I1(n43));
   AN2EHD U84 (.O(n160), 
	.I2(n5), 
	.I1(n43));
   AN2EHD U85 (.O(n162), 
	.I2(n7), 
	.I1(n43));
   AN2EHD U86 (.O(n164), 
	.I2(n24), 
	.I1(n43));
   AN2EHD U87 (.O(n166), 
	.I2(n29), 
	.I1(n43));
   AN2EHD U88 (.O(n168), 
	.I2(n32), 
	.I1(n43));
   AN2EHD U89 (.O(n170), 
	.I2(n34), 
	.I1(n43));
   AN2EHD U90 (.O(n172), 
	.I2(n25), 
	.I1(n43));
   AN2EHD U91 (.O(n175), 
	.I2(n31), 
	.I1(n43));
   AN2EHD U92 (.O(n177), 
	.I2(n35), 
	.I1(n43));
   AN2EHD U93 (.O(n178), 
	.I2(n37), 
	.I1(n43));
   AN2EHD U94 (.O(n180), 
	.I2(n1), 
	.I1(n44));
   AN2EHD U95 (.O(n182), 
	.I2(n2), 
	.I1(n44));
   AN2EHD U96 (.O(n184), 
	.I2(n26), 
	.I1(n44));
   AN2EHD U97 (.O(n186), 
	.I2(n28), 
	.I1(n44));
   AN2EHD U98 (.O(n188), 
	.I2(n3), 
	.I1(n44));
   AN2EHD U99 (.O(n190), 
	.I2(n4), 
	.I1(n44));
   AN2EHD U100 (.O(n192), 
	.I2(n5), 
	.I1(n44));
   AN2EHD U101 (.O(n194), 
	.I2(n7), 
	.I1(n44));
   AN2EHD U102 (.O(n196), 
	.I2(n24), 
	.I1(n44));
   AN2EHD U103 (.O(n198), 
	.I2(n29), 
	.I1(n44));
   AN2EHD U104 (.O(n200), 
	.I2(n32), 
	.I1(n44));
   AN2EHD U105 (.O(n202), 
	.I2(n34), 
	.I1(n44));
   AN2EHD U106 (.O(n204), 
	.I2(n25), 
	.I1(n44));
   AN2EHD U107 (.O(n206), 
	.I2(n31), 
	.I1(n44));
   AN2EHD U108 (.O(n209), 
	.I2(n35), 
	.I1(n44));
   AN2EHD U109 (.O(n211), 
	.I2(n37), 
	.I1(n44));
   AN2EHD U110 (.O(n212), 
	.I2(n1), 
	.I1(n47));
   AN2EHD U111 (.O(n214), 
	.I2(n2), 
	.I1(n47));
   AN2EHD U112 (.O(n216), 
	.I2(n26), 
	.I1(n47));
   AN2EHD U113 (.O(n218), 
	.I2(n28), 
	.I1(n47));
   AN2EHD U114 (.O(n220), 
	.I2(n3), 
	.I1(n47));
   AN2EHD U115 (.O(n222), 
	.I2(n4), 
	.I1(n47));
   AN2EHD U116 (.O(n224), 
	.I2(n5), 
	.I1(n47));
   AN2EHD U117 (.O(n226), 
	.I2(n7), 
	.I1(n47));
   AN2EHD U118 (.O(n228), 
	.I2(n24), 
	.I1(n47));
   AN2EHD U119 (.O(n230), 
	.I2(n29), 
	.I1(n47));
   AN2EHD U120 (.O(n232), 
	.I2(n32), 
	.I1(n47));
   AN2EHD U121 (.O(n234), 
	.I2(n34), 
	.I1(n47));
   AN2EHD U122 (.O(n236), 
	.I2(n25), 
	.I1(n47));
   AN2EHD U123 (.O(n238), 
	.I2(n31), 
	.I1(n47));
   AN2EHD U124 (.O(n240), 
	.I2(n35), 
	.I1(n47));
   AN2EHD U125 (.O(n242), 
	.I2(n37), 
	.I1(n47));
   AN2EHD U126 (.O(n244), 
	.I2(n1), 
	.I1(n50));
   AN2EHD U127 (.O(n245), 
	.I2(n2), 
	.I1(n50));
   AN2EHD U128 (.O(n247), 
	.I2(n26), 
	.I1(n50));
   AN2EHD U129 (.O(n249), 
	.I2(n28), 
	.I1(n50));
   AN2EHD U130 (.O(n251), 
	.I2(n3), 
	.I1(n50));
   AN2EHD U131 (.O(n253), 
	.I2(n4), 
	.I1(n50));
   AN2EHD U132 (.O(n255), 
	.I2(n5), 
	.I1(n50));
   AN2EHD U133 (.O(n257), 
	.I2(n7), 
	.I1(n50));
   AN2EHD U134 (.O(n259), 
	.I2(n24), 
	.I1(n50));
   AN2EHD U135 (.O(n261), 
	.I2(n29), 
	.I1(n50));
   AN2EHD U136 (.O(n263), 
	.I2(n32), 
	.I1(n50));
   AN2EHD U137 (.O(n265), 
	.I2(n34), 
	.I1(n50));
   AN2EHD U138 (.O(n267), 
	.I2(n25), 
	.I1(n50));
   AN2EHD U139 (.O(n269), 
	.I2(n31), 
	.I1(n50));
   AN2EHD U140 (.O(n271), 
	.I2(n35), 
	.I1(n50));
   AN2EHD U141 (.O(n273), 
	.I2(n37), 
	.I1(n50));
   AN2EHD U142 (.O(n275), 
	.I2(n1), 
	.I1(n52));
   AN2EHD U143 (.O(n277), 
	.I2(n2), 
	.I1(n52));
   AN2EHD U144 (.O(n278), 
	.I2(n26), 
	.I1(n52));
   AN2EHD U145 (.O(n280), 
	.I2(n28), 
	.I1(n52));
   AN2EHD U146 (.O(n282), 
	.I2(n3), 
	.I1(n52));
   AN2EHD U147 (.O(n284), 
	.I2(n4), 
	.I1(n52));
   AN2EHD U148 (.O(n286), 
	.I2(n5), 
	.I1(n52));
   AN2EHD U149 (.O(n288), 
	.I2(n7), 
	.I1(n52));
   AN2EHD U150 (.O(n290), 
	.I2(n24), 
	.I1(n52));
   AN2EHD U151 (.O(n292), 
	.I2(n29), 
	.I1(n52));
   AN2EHD U152 (.O(n294), 
	.I2(n32), 
	.I1(n52));
   AN2EHD U153 (.O(n296), 
	.I2(n34), 
	.I1(n52));
   AN2EHD U154 (.O(n298), 
	.I2(n25), 
	.I1(n52));
   AN2EHD U155 (.O(n300), 
	.I2(n31), 
	.I1(n52));
   AN2EHD U156 (.O(n302), 
	.I2(n35), 
	.I1(n52));
   AN2EHD U157 (.O(n304), 
	.I2(n37), 
	.I1(n52));
   AN2EHD U158 (.O(n306), 
	.I2(n1), 
	.I1(n46));
   AN2EHD U159 (.O(n308), 
	.I2(n2), 
	.I1(n46));
   AN2EHD U160 (.O(n310), 
	.I2(n26), 
	.I1(n46));
   AN2EHD U161 (.O(n311), 
	.I2(n28), 
	.I1(n46));
   AN2EHD U162 (.O(n313), 
	.I2(n3), 
	.I1(n46));
   AN2EHD U163 (.O(n315), 
	.I2(n4), 
	.I1(n46));
   AN2EHD U164 (.O(n317), 
	.I2(n5), 
	.I1(n46));
   AN2EHD U165 (.O(n319), 
	.I2(n7), 
	.I1(n46));
   AN2EHD U166 (.O(n321), 
	.I2(n24), 
	.I1(n46));
   AN2EHD U167 (.O(n323), 
	.I2(n29), 
	.I1(n46));
   AN2EHD U168 (.O(n325), 
	.I2(n32), 
	.I1(n46));
   AN2EHD U169 (.O(n327), 
	.I2(n34), 
	.I1(n46));
   AN2EHD U170 (.O(n329), 
	.I2(n25), 
	.I1(n46));
   AN2EHD U171 (.O(n331), 
	.I2(n31), 
	.I1(n46));
   AN2EHD U172 (.O(n333), 
	.I2(n35), 
	.I1(n46));
   AN2EHD U173 (.O(n335), 
	.I2(n37), 
	.I1(n46));
   AN2EHD U174 (.O(n337), 
	.I2(n1), 
	.I1(n49));
   AN2EHD U175 (.O(n339), 
	.I2(n2), 
	.I1(n49));
   AN2EHD U176 (.O(n342), 
	.I2(n26), 
	.I1(n49));
   AN2EHD U177 (.O(n344), 
	.I2(n28), 
	.I1(n49));
   AN2EHD U178 (.O(n345), 
	.I2(n3), 
	.I1(n49));
   AN2EHD U179 (.O(n347), 
	.I2(n4), 
	.I1(n49));
   AN2EHD U180 (.O(n349), 
	.I2(n5), 
	.I1(n49));
   AN2EHD U181 (.O(n351), 
	.I2(n7), 
	.I1(n49));
   AN2EHD U182 (.O(n353), 
	.I2(n24), 
	.I1(n49));
   AN2EHD U183 (.O(n355), 
	.I2(n29), 
	.I1(n49));
   AN2EHD U184 (.O(n357), 
	.I2(n32), 
	.I1(n49));
   AN2EHD U185 (.O(n359), 
	.I2(n34), 
	.I1(n49));
   AN2EHD U186 (.O(n361), 
	.I2(n25), 
	.I1(n49));
   AN2EHD U187 (.O(n363), 
	.I2(n31), 
	.I1(n49));
   AN2EHD U188 (.O(n365), 
	.I2(n35), 
	.I1(n49));
   AN2EHD U189 (.O(n367), 
	.I2(n37), 
	.I1(n49));
   AN2EHD U190 (.O(n369), 
	.I2(n1), 
	.I1(n53));
   AN2EHD U191 (.O(n371), 
	.I2(n2), 
	.I1(n53));
   AN2EHD U192 (.O(n373), 
	.I2(n26), 
	.I1(n53));
   AN2EHD U193 (.O(n375), 
	.I2(n28), 
	.I1(n53));
   AN2EHD U194 (.O(n377), 
	.I2(n3), 
	.I1(n53));
   AN2EHD U195 (.O(n378), 
	.I2(n4), 
	.I1(n53));
   AN2EHD U196 (.O(n380), 
	.I2(n5), 
	.I1(n53));
   AN2EHD U197 (.O(n382), 
	.I2(n7), 
	.I1(n53));
   AN2EHD U198 (.O(n384), 
	.I2(n24), 
	.I1(n53));
   AN2EHD U199 (.O(n386), 
	.I2(n29), 
	.I1(n53));
   AN2EHD U200 (.O(n388), 
	.I2(n32), 
	.I1(n53));
   AN2EHD U201 (.O(n390), 
	.I2(n34), 
	.I1(n53));
   AN2EHD U202 (.O(n392), 
	.I2(n25), 
	.I1(n53));
   AN2EHD U203 (.O(n394), 
	.I2(n31), 
	.I1(n53));
   AN2EHD U204 (.O(n396), 
	.I2(n35), 
	.I1(n53));
   AN2EHD U205 (.O(n398), 
	.I2(n37), 
	.I1(n53));
   AN2EHD U206 (.O(n400), 
	.I2(n1), 
	.I1(n55));
   AN2EHD U207 (.O(n402), 
	.I2(n2), 
	.I1(n55));
   AN2EHD U208 (.O(n404), 
	.I2(n26), 
	.I1(n55));
   AN2EHD U209 (.O(n406), 
	.I2(n28), 
	.I1(n55));
   AN2EHD U210 (.O(n408), 
	.I2(n3), 
	.I1(n55));
   AN2EHD U211 (.O(n410), 
	.I2(n4), 
	.I1(n55));
   AN2EHD U212 (.O(n411), 
	.I2(n5), 
	.I1(n55));
   AN2EHD U213 (.O(n413), 
	.I2(n7), 
	.I1(n55));
   AN2EHD U214 (.O(n415), 
	.I2(n24), 
	.I1(n55));
   AN2EHD U215 (.O(n417), 
	.I2(n29), 
	.I1(n55));
   AN2EHD U216 (.O(n419), 
	.I2(n32), 
	.I1(n55));
   AN2EHD U217 (.O(n421), 
	.I2(n34), 
	.I1(n55));
   AN2EHD U218 (.O(n423), 
	.I2(n25), 
	.I1(n55));
   AN2EHD U219 (.O(n425), 
	.I2(n31), 
	.I1(n55));
   AN2EHD U220 (.O(n427), 
	.I2(n35), 
	.I1(n55));
   AN2EHD U221 (.O(n429), 
	.I2(n37), 
	.I1(n55));
   AN2EHD U222 (.O(n431), 
	.I2(n72), 
	.I1(n71));
   AN2EHD U223 (.O(n433), 
	.I2(n431), 
	.I1(n1));
   AN2EHD U224 (.O(n435), 
	.I2(n71), 
	.I1(n106));
   AN2EHD U225 (.O(n437), 
	.I2(n71), 
	.I1(n140));
   AN2EHD U226 (.O(n439), 
	.I2(n71), 
	.I1(n174));
   AN2EHD U227 (.O(n441), 
	.I2(n431), 
	.I1(n2));
   AN2EHD U228 (.O(n443), 
	.I2(n431), 
	.I1(n26));
   AN2EHD U229 (.O(n444), 
	.I2(n431), 
	.I1(n28));
   AN2EHD U230 (.O(n446), 
	.I2(n431), 
	.I1(n3));
   AN2EHD U231 (.O(n448), 
	.I2(n431), 
	.I1(n4));
   AN2EHD U232 (.O(n450), 
	.I2(n431), 
	.I1(n5));
   AN2EHD U233 (.O(n452), 
	.I2(n431), 
	.I1(n7));
   AN2EHD U234 (.O(n454), 
	.I2(n431), 
	.I1(n24));
   AN2EHD U235 (.O(n456), 
	.I2(n431), 
	.I1(n29));
   AN2EHD U236 (.O(n458), 
	.I2(n431), 
	.I1(n32));
   AN2EHD U237 (.O(n460), 
	.I2(n431), 
	.I1(n34));
   AN2EHD U238 (.O(n462), 
	.I2(n431), 
	.I1(n25));
   AN2EHD U239 (.O(n464), 
	.I2(n431), 
	.I1(n31));
   AN2EHD U240 (.O(n466), 
	.I2(n431), 
	.I1(n35));
   AN2EHD U241 (.O(n468), 
	.I2(n431), 
	.I1(n37));
   AN2EHD U242 (.O(n470), 
	.I2(n1), 
	.I1(n435));
   AN2EHD U243 (.O(n472), 
	.I2(n2), 
	.I1(n435));
   AN2EHD U244 (.O(n475), 
	.I2(n26), 
	.I1(n435));
   AN2EHD U245 (.O(n477), 
	.I2(n28), 
	.I1(n435));
   AN2EHD U246 (.O(n478), 
	.I2(n3), 
	.I1(n435));
   AN2EHD U247 (.O(n480), 
	.I2(n4), 
	.I1(n435));
   AN2EHD U248 (.O(n482), 
	.I2(n5), 
	.I1(n435));
   AN2EHD U249 (.O(n484), 
	.I2(n7), 
	.I1(n435));
   AN2EHD U250 (.O(n486), 
	.I2(n24), 
	.I1(n435));
   AN2EHD U251 (.O(n488), 
	.I2(n29), 
	.I1(n435));
   AN2EHD U252 (.O(n490), 
	.I2(n32), 
	.I1(n435));
   AN2EHD U253 (.O(n492), 
	.I2(n34), 
	.I1(n435));
   AN2EHD U254 (.O(n494), 
	.I2(n25), 
	.I1(n435));
   AN2EHD U255 (.O(n496), 
	.I2(n31), 
	.I1(n435));
   AN2EHD U256 (.O(n498), 
	.I2(n35), 
	.I1(n435));
   AN2EHD U257 (.O(n500), 
	.I2(n37), 
	.I1(n435));
   AN2EHD U258 (.O(n502), 
	.I2(n1), 
	.I1(n437));
   AN2EHD U259 (.O(n504), 
	.I2(n2), 
	.I1(n437));
   AN2EHD U260 (.O(n506), 
	.I2(n26), 
	.I1(n437));
   AN2EHD U261 (.O(n508), 
	.I2(n28), 
	.I1(n437));
   AN2EHD U262 (.O(n510), 
	.I2(n3), 
	.I1(n437));
   AN2EHD U263 (.O(n511), 
	.I2(n4), 
	.I1(n437));
   AN2EHD U264 (.O(n513), 
	.I2(n5), 
	.I1(n437));
   AN2EHD U265 (.O(n515), 
	.I2(n7), 
	.I1(n437));
   AN2EHD U266 (.O(n517), 
	.I2(n24), 
	.I1(n437));
   AN2EHD U267 (.O(n519), 
	.I2(n29), 
	.I1(n437));
   AN2EHD U268 (.O(n521), 
	.I2(n32), 
	.I1(n437));
   AN2EHD U269 (.O(n523), 
	.I2(n34), 
	.I1(n437));
   AN2EHD U270 (.O(n525), 
	.I2(n25), 
	.I1(n437));
   AN2EHD U271 (.O(n527), 
	.I2(n31), 
	.I1(n437));
   AN2EHD U272 (.O(n529), 
	.I2(n35), 
	.I1(n437));
   AN2EHD U273 (.O(n531), 
	.I2(n37), 
	.I1(n437));
   AN2EHD U274 (.O(n533), 
	.I2(n1), 
	.I1(n439));
   AN2EHD U275 (.O(n535), 
	.I2(n2), 
	.I1(n439));
   AN2EHD U276 (.O(n537), 
	.I2(n26), 
	.I1(n439));
   AN2EHD U277 (.O(n539), 
	.I2(n28), 
	.I1(n439));
   AN2EHD U278 (.O(n541), 
	.I2(n3), 
	.I1(n439));
   AN2EHD U279 (.O(n543), 
	.I2(n4), 
	.I1(n439));
   AN2EHD U280 (.O(n546), 
	.I2(n5), 
	.I1(n439));
   AN2EHD U281 (.O(n549), 
	.I2(n7), 
	.I1(n439));
   AN2EHD U282 (.O(n552), 
	.I2(n24), 
	.I1(n439));
   AN2EHD U283 (.O(n555), 
	.I2(n29), 
	.I1(n439));
   AN2EHD U284 (.O(n558), 
	.I2(n32), 
	.I1(n439));
   AN2EHD U285 (.O(n560), 
	.I2(n34), 
	.I1(n439));
   AN2EHD U286 (.O(n562), 
	.I2(n25), 
	.I1(n439));
   AN2EHD U287 (.O(n564), 
	.I2(n31), 
	.I1(n439));
   AN2EHD U288 (.O(n567), 
	.I2(n35), 
	.I1(n439));
   AN2EHD U289 (.O(n569), 
	.I2(n37), 
	.I1(n439));
   ND2DHD U751 (.O(n27), 
	.I2(mem_write_en), 
	.I1(n441));
   ND2DHD U753 (.O(n30), 
	.I2(mem_write_en), 
	.I1(n443));
   ND2DHD U755 (.O(n33), 
	.I2(mem_write_en), 
	.I1(n444));
   ND2DHD U757 (.O(n36), 
	.I2(mem_write_en), 
	.I1(n446));
   ND2DHD U759 (.O(n39), 
	.I2(mem_write_en), 
	.I1(n448));
   ND2DHD U761 (.O(n42), 
	.I2(mem_write_en), 
	.I1(n450));
   ND2DHD U763 (.O(n45), 
	.I2(mem_write_en), 
	.I1(n452));
   ND2DHD U765 (.O(n48), 
	.I2(mem_write_en), 
	.I1(n454));
   ND2DHD U767 (.O(n51), 
	.I2(mem_write_en), 
	.I1(n456));
   ND2DHD U769 (.O(n54), 
	.I2(mem_write_en), 
	.I1(n458));
   ND2DHD U771 (.O(n57), 
	.I2(mem_write_en), 
	.I1(n460));
   ND2DHD U773 (.O(n60), 
	.I2(mem_write_en), 
	.I1(n462));
   ND2DHD U775 (.O(n63), 
	.I2(mem_write_en), 
	.I1(n464));
   ND2DHD U777 (.O(n66), 
	.I2(mem_write_en), 
	.I1(n466));
   ND2DHD U779 (.O(n69), 
	.I2(mem_write_en), 
	.I1(n468));
   ND2DHD U781 (.O(n74), 
	.I2(mem_write_en), 
	.I1(n470));
   ND2DHD U783 (.O(n77), 
	.I2(mem_write_en), 
	.I1(n472));
   ND2DHD U785 (.O(n79), 
	.I2(mem_write_en), 
	.I1(n475));
   ND2DHD U787 (.O(n81), 
	.I2(mem_write_en), 
	.I1(n477));
   ND2DHD U789 (.O(n83), 
	.I2(FE_OFN94_mem_write), 
	.I1(n478));
   ND2DHD U791 (.O(n85), 
	.I2(FE_OFN94_mem_write), 
	.I1(n480));
   ND2DHD U793 (.O(n87), 
	.I2(FE_OFN94_mem_write), 
	.I1(n482));
   ND2DHD U795 (.O(n89), 
	.I2(FE_OFN94_mem_write), 
	.I1(n484));
   ND2DHD U797 (.O(n91), 
	.I2(mem_write_en), 
	.I1(n486));
   ND2DHD U799 (.O(n93), 
	.I2(mem_write_en), 
	.I1(n488));
   ND2DHD U801 (.O(n95), 
	.I2(mem_write_en), 
	.I1(n490));
   ND2DHD U803 (.O(n97), 
	.I2(mem_write_en), 
	.I1(n492));
   ND2DHD U805 (.O(n99), 
	.I2(mem_write_en), 
	.I1(n494));
   ND2DHD U807 (.O(n101), 
	.I2(mem_write_en), 
	.I1(n496));
   ND2DHD U809 (.O(n103), 
	.I2(mem_write_en), 
	.I1(n498));
   ND2DHD U811 (.O(n105), 
	.I2(mem_write_en), 
	.I1(n500));
   ND2DHD U813 (.O(n108), 
	.I2(mem_write_en), 
	.I1(n502));
   ND2DHD U815 (.O(n111), 
	.I2(mem_write_en), 
	.I1(n504));
   ND2DHD U817 (.O(n113), 
	.I2(mem_write_en), 
	.I1(n506));
   ND2DHD U819 (.O(n115), 
	.I2(mem_write_en), 
	.I1(n508));
   ND2DHD U821 (.O(n117), 
	.I2(mem_write_en), 
	.I1(n510));
   ND2DHD U823 (.O(n119), 
	.I2(mem_write_en), 
	.I1(n511));
   ND2DHD U825 (.O(n121), 
	.I2(mem_write_en), 
	.I1(n513));
   ND2DHD U827 (.O(n123), 
	.I2(mem_write_en), 
	.I1(n515));
   ND2DHD U829 (.O(n125), 
	.I2(FE_OFN94_mem_write), 
	.I1(n517));
   ND2DHD U831 (.O(n127), 
	.I2(FE_OFN94_mem_write), 
	.I1(n519));
   ND2DHD U833 (.O(n129), 
	.I2(FE_OFN94_mem_write), 
	.I1(n521));
   ND2DHD U835 (.O(n131), 
	.I2(FE_OFN94_mem_write), 
	.I1(n523));
   ND2DHD U837 (.O(n133), 
	.I2(FE_OFN94_mem_write), 
	.I1(n525));
   ND2DHD U839 (.O(n135), 
	.I2(FE_OFN94_mem_write), 
	.I1(n527));
   ND2DHD U841 (.O(n137), 
	.I2(mem_write_en), 
	.I1(n529));
   ND2DHD U843 (.O(n139), 
	.I2(FE_OFN94_mem_write), 
	.I1(n531));
   ND2DHD U845 (.O(n142), 
	.I2(FE_OFN94_mem_write), 
	.I1(n533));
   ND2DHD U847 (.O(n145), 
	.I2(FE_OFN94_mem_write), 
	.I1(n535));
   ND2DHD U849 (.O(n147), 
	.I2(FE_OFN94_mem_write), 
	.I1(n537));
   ND2DHD U851 (.O(n149), 
	.I2(FE_OFN94_mem_write), 
	.I1(n539));
   ND2DHD U853 (.O(n151), 
	.I2(FE_OFN94_mem_write), 
	.I1(n541));
   ND2DHD U855 (.O(n153), 
	.I2(FE_OFN94_mem_write), 
	.I1(n543));
   ND2DHD U857 (.O(n155), 
	.I2(FE_OFN94_mem_write), 
	.I1(n546));
   ND2DHD U859 (.O(n157), 
	.I2(FE_OFN94_mem_write), 
	.I1(n549));
   ND2DHD U861 (.O(n159), 
	.I2(FE_OFN94_mem_write), 
	.I1(n552));
   ND2DHD U863 (.O(n161), 
	.I2(FE_OFN94_mem_write), 
	.I1(n555));
   ND2DHD U865 (.O(n163), 
	.I2(FE_OFN94_mem_write), 
	.I1(n558));
   ND2DHD U867 (.O(n165), 
	.I2(FE_OFN94_mem_write), 
	.I1(n560));
   ND2DHD U869 (.O(n167), 
	.I2(FE_OFN94_mem_write), 
	.I1(n562));
   ND2DHD U871 (.O(n169), 
	.I2(FE_OFN94_mem_write), 
	.I1(n564));
   ND2DHD U873 (.O(n171), 
	.I2(FE_OFN94_mem_write), 
	.I1(n567));
   ND2DHD U875 (.O(n173), 
	.I2(FE_OFN94_mem_write), 
	.I1(n569));
   ND2DHD U877 (.O(n176), 
	.I2(FE_OFN94_mem_write), 
	.I1(n56));
   ND2DHD U879 (.O(n179), 
	.I2(FE_OFN94_mem_write), 
	.I1(n58));
   ND2DHD U881 (.O(n181), 
	.I2(FE_OFN94_mem_write), 
	.I1(n59));
   ND2DHD U883 (.O(n183), 
	.I2(FE_OFN94_mem_write), 
	.I1(n61));
   ND2DHD U885 (.O(n185), 
	.I2(FE_OFN94_mem_write), 
	.I1(n62));
   ND2DHD U887 (.O(n187), 
	.I2(FE_OFN94_mem_write), 
	.I1(n64));
   ND2DHD U889 (.O(n189), 
	.I2(FE_OFN94_mem_write), 
	.I1(n65));
   ND2DHD U891 (.O(n191), 
	.I2(FE_OFN94_mem_write), 
	.I1(n67));
   ND2DHD U893 (.O(n193), 
	.I2(FE_OFN92_mem_write), 
	.I1(n68));
   ND2DHD U895 (.O(n195), 
	.I2(FE_OFN92_mem_write), 
	.I1(n70));
   ND2DHD U897 (.O(n197), 
	.I2(FE_OFN92_mem_write), 
	.I1(n73));
   ND2DHD U899 (.O(n199), 
	.I2(FE_OFN92_mem_write), 
	.I1(n75));
   ND2DHD U901 (.O(n201), 
	.I2(FE_OFN92_mem_write), 
	.I1(n76));
   ND2DHD U903 (.O(n203), 
	.I2(FE_OFN92_mem_write), 
	.I1(n78));
   ND2DHD U905 (.O(n205), 
	.I2(FE_OFN92_mem_write), 
	.I1(n80));
   ND2DHD U907 (.O(n207), 
	.I2(FE_OFN92_mem_write), 
	.I1(n82));
   ND2DHD U909 (.O(n210), 
	.I2(FE_OFN94_mem_write), 
	.I1(n84));
   ND2DHD U911 (.O(n213), 
	.I2(FE_OFN94_mem_write), 
	.I1(n86));
   ND2DHD U913 (.O(n215), 
	.I2(FE_OFN94_mem_write), 
	.I1(n88));
   ND2DHD U915 (.O(n217), 
	.I2(FE_OFN94_mem_write), 
	.I1(n90));
   ND2DHD U917 (.O(n219), 
	.I2(FE_OFN94_mem_write), 
	.I1(n92));
   ND2DHD U919 (.O(n221), 
	.I2(FE_OFN94_mem_write), 
	.I1(n94));
   ND2DHD U921 (.O(n223), 
	.I2(FE_OFN94_mem_write), 
	.I1(n96));
   ND2DHD U923 (.O(n225), 
	.I2(FE_OFN94_mem_write), 
	.I1(n98));
   ND2DHD U925 (.O(n227), 
	.I2(FE_OFN94_mem_write), 
	.I1(n100));
   ND2DHD U927 (.O(n229), 
	.I2(FE_OFN94_mem_write), 
	.I1(n102));
   ND2DHD U929 (.O(n231), 
	.I2(FE_OFN94_mem_write), 
	.I1(n104));
   ND2DHD U931 (.O(n233), 
	.I2(FE_OFN94_mem_write), 
	.I1(n107));
   ND2DHD U933 (.O(n235), 
	.I2(FE_OFN94_mem_write), 
	.I1(n109));
   ND2DHD U935 (.O(n237), 
	.I2(FE_OFN94_mem_write), 
	.I1(n110));
   ND2DHD U937 (.O(n239), 
	.I2(FE_OFN94_mem_write), 
	.I1(n112));
   ND2DHD U939 (.O(n241), 
	.I2(FE_OFN94_mem_write), 
	.I1(n114));
   ND2DHD U941 (.O(n243), 
	.I2(FE_OFN92_mem_write), 
	.I1(n116));
   ND2DHD U943 (.O(n246), 
	.I2(FE_OFN92_mem_write), 
	.I1(n118));
   ND2DHD U945 (.O(n248), 
	.I2(FE_OFN92_mem_write), 
	.I1(n120));
   ND2DHD U947 (.O(n250), 
	.I2(FE_OFN92_mem_write), 
	.I1(n122));
   ND2DHD U949 (.O(n252), 
	.I2(FE_OFN94_mem_write), 
	.I1(n124));
   ND2DHD U951 (.O(n254), 
	.I2(FE_OFN94_mem_write), 
	.I1(n126));
   ND2DHD U953 (.O(n256), 
	.I2(FE_OFN94_mem_write), 
	.I1(n128));
   ND2DHD U955 (.O(n258), 
	.I2(FE_OFN94_mem_write), 
	.I1(n130));
   ND2DHD U957 (.O(n260), 
	.I2(FE_OFN94_mem_write), 
	.I1(n132));
   ND2DHD U959 (.O(n262), 
	.I2(FE_OFN94_mem_write), 
	.I1(n134));
   ND2DHD U961 (.O(n264), 
	.I2(FE_OFN94_mem_write), 
	.I1(n136));
   ND2DHD U963 (.O(n266), 
	.I2(FE_OFN94_mem_write), 
	.I1(n138));
   ND2DHD U965 (.O(n268), 
	.I2(FE_OFN94_mem_write), 
	.I1(n141));
   ND2DHD U967 (.O(n270), 
	.I2(FE_OFN94_mem_write), 
	.I1(n143));
   ND2DHD U969 (.O(n272), 
	.I2(FE_OFN94_mem_write), 
	.I1(n144));
   ND2DHD U971 (.O(n274), 
	.I2(FE_OFN94_mem_write), 
	.I1(n146));
   ND2DHD U973 (.O(n276), 
	.I2(FE_OFN92_mem_write), 
	.I1(n148));
   ND2DHD U975 (.O(n279), 
	.I2(FE_OFN92_mem_write), 
	.I1(n150));
   ND2DHD U977 (.O(n281), 
	.I2(FE_OFN92_mem_write), 
	.I1(n152));
   ND2DHD U979 (.O(n283), 
	.I2(FE_OFN92_mem_write), 
	.I1(n154));
   ND2DHD U981 (.O(n285), 
	.I2(FE_OFN94_mem_write), 
	.I1(n156));
   ND2DHD U983 (.O(n287), 
	.I2(FE_OFN94_mem_write), 
	.I1(n158));
   ND2DHD U985 (.O(n289), 
	.I2(FE_OFN94_mem_write), 
	.I1(n160));
   ND2DHD U987 (.O(n291), 
	.I2(FE_OFN94_mem_write), 
	.I1(n162));
   ND2DHD U989 (.O(n293), 
	.I2(FE_OFN94_mem_write), 
	.I1(n164));
   ND2DHD U991 (.O(n295), 
	.I2(FE_OFN94_mem_write), 
	.I1(n166));
   ND2DHD U993 (.O(n297), 
	.I2(FE_OFN94_mem_write), 
	.I1(n168));
   ND2DHD U995 (.O(n299), 
	.I2(FE_OFN94_mem_write), 
	.I1(n170));
   ND2DHD U997 (.O(n301), 
	.I2(FE_OFN94_mem_write), 
	.I1(n172));
   ND2DHD U999 (.O(n303), 
	.I2(FE_OFN94_mem_write), 
	.I1(n175));
   ND2DHD U1001 (.O(n305), 
	.I2(FE_OFN94_mem_write), 
	.I1(n177));
   ND2DHD U1003 (.O(n307), 
	.I2(FE_OFN94_mem_write), 
	.I1(n178));
   ND2DHD U1005 (.O(n309), 
	.I2(FE_OFN93_mem_write), 
	.I1(n180));
   ND2DHD U1007 (.O(n312), 
	.I2(FE_OFN93_mem_write), 
	.I1(n182));
   ND2DHD U1009 (.O(n314), 
	.I2(FE_OFN93_mem_write), 
	.I1(n184));
   ND2DHD U1011 (.O(n316), 
	.I2(FE_OFN93_mem_write), 
	.I1(n186));
   ND2DHD U1013 (.O(n318), 
	.I2(FE_OFN93_mem_write), 
	.I1(n188));
   ND2DHD U1015 (.O(n320), 
	.I2(FE_OFN93_mem_write), 
	.I1(n190));
   ND2DHD U1017 (.O(n322), 
	.I2(FE_OFN93_mem_write), 
	.I1(n192));
   ND2DHD U1019 (.O(n324), 
	.I2(FE_OFN93_mem_write), 
	.I1(n194));
   ND2DHD U1021 (.O(n326), 
	.I2(FE_OFN93_mem_write), 
	.I1(n196));
   ND2DHD U1023 (.O(n328), 
	.I2(FE_OFN93_mem_write), 
	.I1(n198));
   ND2DHD U1025 (.O(n334), 
	.I2(FE_OFN93_mem_write), 
	.I1(n204));
   ND2DHD U1027 (.O(n338), 
	.I2(FE_OFN93_mem_write), 
	.I1(n209));
   ND2DHD U1029 (.O(n340), 
	.I2(FE_OFN93_mem_write), 
	.I1(n211));
   ND2DHD U1031 (.O(n343), 
	.I2(FE_OFN93_mem_write), 
	.I1(n212));
   ND2DHD U1033 (.O(n346), 
	.I2(FE_OFN93_mem_write), 
	.I1(n214));
   ND2DHD U1035 (.O(n348), 
	.I2(FE_OFN93_mem_write), 
	.I1(n216));
   ND2DHD U1037 (.O(n350), 
	.I2(FE_OFN93_mem_write), 
	.I1(n218));
   ND2DHD U1039 (.O(n352), 
	.I2(mem_write_en), 
	.I1(n220));
   ND2DHD U1041 (.O(n354), 
	.I2(mem_write_en), 
	.I1(n222));
   ND2DHD U1043 (.O(n356), 
	.I2(mem_write_en), 
	.I1(n224));
   ND2DHD U1045 (.O(n358), 
	.I2(mem_write_en), 
	.I1(n226));
   ND2DHD U1047 (.O(n360), 
	.I2(mem_write_en), 
	.I1(n228));
   ND2DHD U1049 (.O(n362), 
	.I2(mem_write_en), 
	.I1(n230));
   ND2DHD U1051 (.O(n364), 
	.I2(mem_write_en), 
	.I1(n232));
   ND2DHD U1053 (.O(n366), 
	.I2(mem_write_en), 
	.I1(n234));
   ND2DHD U1055 (.O(n368), 
	.I2(FE_OFN93_mem_write), 
	.I1(n236));
   ND2DHD U1057 (.O(n370), 
	.I2(FE_OFN93_mem_write), 
	.I1(n238));
   ND2DHD U1059 (.O(n372), 
	.I2(FE_OFN93_mem_write), 
	.I1(n240));
   ND2DHD U1061 (.O(n374), 
	.I2(FE_OFN93_mem_write), 
	.I1(n242));
   ND2DHD U1063 (.O(n376), 
	.I2(FE_OFN93_mem_write), 
	.I1(n244));
   ND2DHD U1065 (.O(n379), 
	.I2(FE_OFN93_mem_write), 
	.I1(n245));
   ND2DHD U1067 (.O(n381), 
	.I2(FE_OFN93_mem_write), 
	.I1(n247));
   ND2DHD U1069 (.O(n383), 
	.I2(FE_OFN93_mem_write), 
	.I1(n249));
   ND2DHD U1071 (.O(n385), 
	.I2(FE_OFN93_mem_write), 
	.I1(n251));
   ND2DHD U1073 (.O(n387), 
	.I2(FE_OFN93_mem_write), 
	.I1(n253));
   ND2DHD U1075 (.O(n389), 
	.I2(FE_OFN93_mem_write), 
	.I1(n255));
   ND2DHD U1077 (.O(n391), 
	.I2(FE_OFN93_mem_write), 
	.I1(n257));
   ND2DHD U1079 (.O(n393), 
	.I2(FE_OFN93_mem_write), 
	.I1(n259));
   ND2DHD U1081 (.O(n395), 
	.I2(FE_OFN93_mem_write), 
	.I1(n261));
   ND2DHD U1083 (.O(n397), 
	.I2(FE_OFN93_mem_write), 
	.I1(n263));
   ND2DHD U1085 (.O(n399), 
	.I2(FE_OFN93_mem_write), 
	.I1(n265));
   ND2DHD U1087 (.O(n401), 
	.I2(FE_OFN93_mem_write), 
	.I1(n267));
   ND2DHD U1089 (.O(n403), 
	.I2(FE_OFN93_mem_write), 
	.I1(n269));
   ND2DHD U1091 (.O(n405), 
	.I2(FE_OFN93_mem_write), 
	.I1(n271));
   ND2DHD U1093 (.O(n407), 
	.I2(FE_OFN93_mem_write), 
	.I1(n273));
   ND2DHD U1095 (.O(n409), 
	.I2(mem_write_en), 
	.I1(n275));
   ND2DHD U1097 (.O(n412), 
	.I2(mem_write_en), 
	.I1(n277));
   ND2DHD U1099 (.O(n414), 
	.I2(mem_write_en), 
	.I1(n278));
   ND2DHD U1101 (.O(n416), 
	.I2(mem_write_en), 
	.I1(n280));
   ND2DHD U1103 (.O(n418), 
	.I2(FE_OFN93_mem_write), 
	.I1(n282));
   ND2DHD U1105 (.O(n420), 
	.I2(FE_OFN93_mem_write), 
	.I1(n284));
   ND2DHD U1107 (.O(n422), 
	.I2(FE_OFN93_mem_write), 
	.I1(n286));
   ND2DHD U1109 (.O(n424), 
	.I2(FE_OFN93_mem_write), 
	.I1(n288));
   ND2DHD U1111 (.O(n426), 
	.I2(FE_OFN93_mem_write), 
	.I1(n290));
   ND2DHD U1113 (.O(n428), 
	.I2(FE_OFN93_mem_write), 
	.I1(n292));
   ND2DHD U1115 (.O(n430), 
	.I2(FE_OFN93_mem_write), 
	.I1(n294));
   ND2DHD U1117 (.O(n432), 
	.I2(FE_OFN93_mem_write), 
	.I1(n296));
   ND2DHD U1119 (.O(n434), 
	.I2(FE_OFN93_mem_write), 
	.I1(n298));
   ND2DHD U1121 (.O(n436), 
	.I2(FE_OFN93_mem_write), 
	.I1(n300));
   ND2DHD U1123 (.O(n438), 
	.I2(FE_OFN93_mem_write), 
	.I1(n302));
   ND2DHD U1125 (.O(n440), 
	.I2(FE_OFN93_mem_write), 
	.I1(n304));
   ND2DHD U1127 (.O(n442), 
	.I2(FE_OFN92_mem_write), 
	.I1(n306));
   ND2DHD U1129 (.O(n445), 
	.I2(FE_OFN92_mem_write), 
	.I1(n308));
   ND2DHD U1131 (.O(n447), 
	.I2(FE_OFN92_mem_write), 
	.I1(n310));
   ND2DHD U1133 (.O(n449), 
	.I2(FE_OFN92_mem_write), 
	.I1(n311));
   ND2DHD U1135 (.O(n451), 
	.I2(FE_OFN92_mem_write), 
	.I1(n313));
   ND2DHD U1137 (.O(n453), 
	.I2(FE_OFN92_mem_write), 
	.I1(n315));
   ND2DHD U1139 (.O(n455), 
	.I2(FE_OFN92_mem_write), 
	.I1(n317));
   ND2DHD U1141 (.O(n457), 
	.I2(FE_OFN92_mem_write), 
	.I1(n319));
   ND2DHD U1143 (.O(n459), 
	.I2(FE_OFN92_mem_write), 
	.I1(n321));
   ND2DHD U1145 (.O(n461), 
	.I2(FE_OFN92_mem_write), 
	.I1(n323));
   ND2DHD U1147 (.O(n463), 
	.I2(FE_OFN92_mem_write), 
	.I1(n325));
   ND2DHD U1149 (.O(n465), 
	.I2(FE_OFN92_mem_write), 
	.I1(n327));
   ND2DHD U1151 (.O(n467), 
	.I2(FE_OFN92_mem_write), 
	.I1(n329));
   ND2DHD U1153 (.O(n469), 
	.I2(FE_OFN92_mem_write), 
	.I1(n331));
   ND2DHD U1155 (.O(n471), 
	.I2(FE_OFN92_mem_write), 
	.I1(n333));
   ND2DHD U1157 (.O(n473), 
	.I2(FE_OFN92_mem_write), 
	.I1(n335));
   ND2DHD U1159 (.O(n476), 
	.I2(FE_OFN92_mem_write), 
	.I1(n337));
   ND2DHD U1161 (.O(n479), 
	.I2(FE_OFN92_mem_write), 
	.I1(n339));
   ND2DHD U1163 (.O(n481), 
	.I2(FE_OFN92_mem_write), 
	.I1(n342));
   ND2DHD U1165 (.O(n483), 
	.I2(FE_OFN92_mem_write), 
	.I1(n344));
   ND2DHD U1167 (.O(n485), 
	.I2(FE_OFN92_mem_write), 
	.I1(n345));
   ND2DHD U1169 (.O(n487), 
	.I2(FE_OFN92_mem_write), 
	.I1(n347));
   ND2DHD U1171 (.O(n489), 
	.I2(FE_OFN92_mem_write), 
	.I1(n349));
   ND2DHD U1173 (.O(n491), 
	.I2(FE_OFN92_mem_write), 
	.I1(n351));
   ND2DHD U1175 (.O(n493), 
	.I2(FE_OFN92_mem_write), 
	.I1(n353));
   ND2DHD U1177 (.O(n495), 
	.I2(FE_OFN92_mem_write), 
	.I1(n355));
   ND2DHD U1179 (.O(n497), 
	.I2(FE_OFN92_mem_write), 
	.I1(n357));
   ND2DHD U1181 (.O(n499), 
	.I2(FE_OFN92_mem_write), 
	.I1(n359));
   ND2DHD U1183 (.O(n501), 
	.I2(FE_OFN92_mem_write), 
	.I1(n361));
   ND2DHD U1185 (.O(n503), 
	.I2(FE_OFN92_mem_write), 
	.I1(n363));
   ND2DHD U1187 (.O(n505), 
	.I2(FE_OFN92_mem_write), 
	.I1(n365));
   ND2DHD U1189 (.O(n507), 
	.I2(FE_OFN92_mem_write), 
	.I1(n367));
   ND2DHD U1191 (.O(n509), 
	.I2(FE_OFN92_mem_write), 
	.I1(n369));
   ND2DHD U1193 (.O(n512), 
	.I2(FE_OFN92_mem_write), 
	.I1(n371));
   ND2DHD U1195 (.O(n514), 
	.I2(FE_OFN92_mem_write), 
	.I1(n373));
   ND2DHD U1197 (.O(n516), 
	.I2(FE_OFN92_mem_write), 
	.I1(n375));
   ND2DHD U1199 (.O(n518), 
	.I2(FE_OFN92_mem_write), 
	.I1(n377));
   ND2DHD U1201 (.O(n520), 
	.I2(FE_OFN92_mem_write), 
	.I1(n378));
   ND2DHD U1203 (.O(n522), 
	.I2(FE_OFN92_mem_write), 
	.I1(n380));
   ND2DHD U1205 (.O(n524), 
	.I2(FE_OFN92_mem_write), 
	.I1(n382));
   ND2DHD U1207 (.O(n526), 
	.I2(FE_OFN93_mem_write), 
	.I1(n384));
   ND2DHD U1209 (.O(n528), 
	.I2(FE_OFN93_mem_write), 
	.I1(n386));
   ND2DHD U1211 (.O(n530), 
	.I2(FE_OFN93_mem_write), 
	.I1(n388));
   ND2DHD U1213 (.O(n532), 
	.I2(FE_OFN93_mem_write), 
	.I1(n390));
   ND2DHD U1215 (.O(n534), 
	.I2(FE_OFN93_mem_write), 
	.I1(n392));
   ND2DHD U1217 (.O(n536), 
	.I2(FE_OFN93_mem_write), 
	.I1(n394));
   ND2DHD U1219 (.O(n538), 
	.I2(FE_OFN93_mem_write), 
	.I1(n396));
   ND2DHD U1221 (.O(n540), 
	.I2(FE_OFN93_mem_write), 
	.I1(n398));
   ND2DHD U1223 (.O(n542), 
	.I2(FE_OFN93_mem_write), 
	.I1(n400));
   ND2DHD U1225 (.O(n547), 
	.I2(FE_OFN93_mem_write), 
	.I1(n402));
   ND2DHD U1227 (.O(n550), 
	.I2(FE_OFN93_mem_write), 
	.I1(n404));
   ND2DHD U1229 (.O(n553), 
	.I2(FE_OFN93_mem_write), 
	.I1(n406));
   ND2DHD U1231 (.O(n556), 
	.I2(FE_OFN93_mem_write), 
	.I1(n408));
   ND2DHD U1233 (.O(n559), 
	.I2(FE_OFN93_mem_write), 
	.I1(n410));
   ND2DHD U1235 (.O(n561), 
	.I2(FE_OFN93_mem_write), 
	.I1(n411));
   ND2DHD U1237 (.O(n563), 
	.I2(FE_OFN93_mem_write), 
	.I1(n413));
   ND2DHD U1239 (.O(n565), 
	.I2(FE_OFN92_mem_write), 
	.I1(n415));
   ND2DHD U1241 (.O(n568), 
	.I2(FE_OFN92_mem_write), 
	.I1(n417));
   ND2DHD U1243 (.O(n570), 
	.I2(FE_OFN92_mem_write), 
	.I1(n419));
   ND2DHD U1245 (.O(n572), 
	.I2(FE_OFN92_mem_write), 
	.I1(n421));
   ND2DHD U1247 (.O(n574), 
	.I2(FE_OFN92_mem_write), 
	.I1(n423));
   ND2DHD U1249 (.O(n577), 
	.I2(FE_OFN92_mem_write), 
	.I1(n425));
   ND2DHD U1251 (.O(n579), 
	.I2(FE_OFN92_mem_write), 
	.I1(n427));
   ND2DHD U1253 (.O(n581), 
	.I2(FE_OFN92_mem_write), 
	.I1(n429));
   ND2DHD U1255 (.O(n330), 
	.I2(FE_OFN93_mem_write), 
	.I1(n200));
   ND2DHD U1257 (.O(n332), 
	.I2(FE_OFN93_mem_write), 
	.I1(n202));
   ND2DHD U1259 (.O(n336), 
	.I2(FE_OFN93_mem_write), 
	.I1(n206));
   ND2DHD U1261 (.O(n8), 
	.I2(n433), 
	.I1(mem_write_en));
   BUFEHD U1267 (.O(n6459), 
	.I(N20));
   BUFHHD U1271 (.O(n6136), 
	.I(N22));
   BUFHHD U1272 (.O(n6038), 
	.I(N24));
   AN2EHD U1671 (.O(n140), 
	.I2(n7443), 
	.I1(n7444));
   AN2EHD U1672 (.O(n551), 
	.I2(n7439), 
	.I1(n7440));
   AN2EHD U1673 (.O(n174), 
	.I2(N24), 
	.I1(n7444));
   AN2EHD U1674 (.O(n554), 
	.I2(N20), 
	.I1(n7440));
   NR2CHD U1675 (.O(n72), 
	.I2(n7444), 
	.I1(N24));
   NR2CHD U1676 (.O(n106), 
	.I2(n7444), 
	.I1(n7443));
   NR2BHD U1677 (.O(n544), 
	.I2(n7442), 
	.I1(N22));
   AN2EHD U1678 (.O(n566), 
	.I2(n7441), 
	.I1(n7442));
   AN2EHD U1679 (.O(n575), 
	.I2(N22), 
	.I1(n7442));
   NR2BHD U1680 (.O(n557), 
	.I2(n7442), 
	.I1(n7441));
   NR2CHD U1681 (.O(n545), 
	.I2(n7440), 
	.I1(N20));
   NR2CHD U1682 (.O(n548), 
	.I2(n7440), 
	.I1(n7439));
   INVDHD U1879 (.O(n7443), 
	.I(N24));
   INVDHD U1880 (.O(n7441), 
	.I(N22));
   INVDHD U1881 (.O(n7439), 
	.I(N20));
   BUFIHD U1882 (.O(n7440), 
	.I(N21));
   BUFHHD U1883 (.O(n7442), 
	.I(N23));
   BUFIHD U1884 (.O(n7444), 
	.I(N25));
   NR2CHD U1951 (.O(n71), 
	.I2(N27), 
	.I1(N26));
   NR2CHD U1952 (.O(n208), 
	.I2(N27), 
	.I1(n7445));
   INVDHD U1953 (.O(n7445), 
	.I(N26));
   AN2EHD U1954 (.O(n341), 
	.I2(n7445), 
	.I1(N27));
   AN2EHD U1955 (.O(n474), 
	.I2(N26), 
	.I1(N27));
   BUFEHD U1956 (.O(n6470), 
	.I(N27));
   BUFEHD U1957 (.O(n6469), 
	.I(N26));
   AN2EHD U1990 (.O(mem_read_data[9]), 
	.I2(N4132), 
	.I1(n6471));
   AN2EHD U1991 (.O(mem_read_data[8]), 
	.I2(n6471), 
	.I1(N4133));
   AN2EHD U1992 (.O(mem_read_data[1]), 
	.I2(n6471), 
	.I1(N4140));
   AN2EHD U1993 (.O(mem_read_data[2]), 
	.I2(n6471), 
	.I1(N4139));
   AN2EHD U1994 (.O(mem_read_data[3]), 
	.I2(n6471), 
	.I1(N4138));
   AN2EHD U1995 (.O(mem_read_data[4]), 
	.I2(n6471), 
	.I1(N4137));
   AN2EHD U1996 (.O(mem_read_data[5]), 
	.I2(n6471), 
	.I1(N4136));
   AN2EHD U1997 (.O(mem_read_data[6]), 
	.I2(n6471), 
	.I1(N4135));
   AN2EHD U1998 (.O(mem_read_data[7]), 
	.I2(n6471), 
	.I1(N4134));
   AN2EHD U1999 (.O(mem_read_data[10]), 
	.I2(n6471), 
	.I1(N4131));
   AN2EHD U2000 (.O(mem_read_data[11]), 
	.I2(n6471), 
	.I1(N4130));
   AN2EHD U2001 (.O(mem_read_data[12]), 
	.I2(n6471), 
	.I1(N4129));
   AN2EHD U2002 (.O(mem_read_data[13]), 
	.I2(n6471), 
	.I1(N4128));
   AN2EHD U2003 (.O(mem_read_data[14]), 
	.I2(n6471), 
	.I1(N4127));
   AN2EHD U2004 (.O(mem_read_data[15]), 
	.I2(n6471), 
	.I1(N4126));
   AN2HHD U2005 (.O(n6), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[0]));
   AN2HHD U2006 (.O(n9), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[1]));
   AN2HHD U2007 (.O(n10), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[2]));
   AN2EHD U2008 (.O(n11), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[3]));
   AN2EHD U2009 (.O(n12), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[4]));
   AN2EHD U2010 (.O(n13), 
	.I2(mem_write_en), 
	.I1(mem_write_data[5]));
   AN2HHD U2011 (.O(n14), 
	.I2(mem_write_en), 
	.I1(mem_write_data[6]));
   AN2EHD U2012 (.O(n15), 
	.I2(mem_write_en), 
	.I1(mem_write_data[7]));
   AN2EHD U2013 (.O(n16), 
	.I2(mem_write_en), 
	.I1(mem_write_data[8]));
   AN2HHD U2014 (.O(n17), 
	.I2(mem_write_en), 
	.I1(mem_write_data[9]));
   AN2HHD U2015 (.O(n18), 
	.I2(mem_write_en), 
	.I1(mem_write_data[10]));
   AN2HHD U2016 (.O(n19), 
	.I2(mem_write_en), 
	.I1(mem_write_data[11]));
   AN2EHD U2017 (.O(n20), 
	.I2(mem_write_en), 
	.I1(mem_write_data[12]));
   AN2HHD U2018 (.O(n21), 
	.I2(mem_write_en), 
	.I1(mem_write_data[13]));
   AN2HHD U2019 (.O(n22), 
	.I2(mem_write_en), 
	.I1(mem_write_data[14]));
   AN2HHD U2020 (.O(n23), 
	.I2(mem_write_en), 
	.I1(mem_write_data[15]));
   BUFEHD U2021 (.O(n6471), 
	.I(mem_read));
   AN2EHD U2022 (.O(mem_read_data[0]), 
	.I2(n6471), 
	.I1(N4141));
   AO22CHD U2023 (.O(n598), 
	.B2(n27), 
	.B1(\ram[1][0] ), 
	.A2(n6), 
	.A1(n441));
   AO22CHD U2024 (.O(n599), 
	.B2(n27), 
	.B1(\ram[1][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n441));
   AO22CHD U2025 (.O(n600), 
	.B2(n27), 
	.B1(\ram[1][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n441));
   AO22CHD U2026 (.O(n601), 
	.B2(n27), 
	.B1(\ram[1][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n441));
   AO22CHD U2027 (.O(n602), 
	.B2(n27), 
	.B1(\ram[1][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n441));
   AO22CHD U2028 (.O(n603), 
	.B2(n27), 
	.B1(\ram[1][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n441));
   AO22CHD U2029 (.O(n604), 
	.B2(n27), 
	.B1(\ram[1][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n441));
   AO22CHD U2030 (.O(n605), 
	.B2(n27), 
	.B1(\ram[1][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n441));
   AO22CHD U2031 (.O(n606), 
	.B2(n27), 
	.B1(\ram[1][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n441));
   AO22CHD U2032 (.O(n607), 
	.B2(n27), 
	.B1(\ram[1][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n441));
   AO22CHD U2033 (.O(n608), 
	.B2(n27), 
	.B1(\ram[1][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n441));
   AO22CHD U2034 (.O(n609), 
	.B2(n27), 
	.B1(\ram[1][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n441));
   AO22CHD U2035 (.O(n610), 
	.B2(n27), 
	.B1(\ram[1][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n441));
   AO22CHD U2036 (.O(n611), 
	.B2(n27), 
	.B1(\ram[1][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n441));
   AO22CHD U2037 (.O(n612), 
	.B2(n27), 
	.B1(\ram[1][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n441));
   AO22CHD U2038 (.O(n613), 
	.B2(n27), 
	.B1(\ram[1][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n441));
   AO22CHD U2039 (.O(n614), 
	.B2(n30), 
	.B1(\ram[2][0] ), 
	.A2(n6), 
	.A1(n443));
   AO22CHD U2040 (.O(n615), 
	.B2(n30), 
	.B1(\ram[2][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n443));
   AO22CHD U2041 (.O(n616), 
	.B2(n30), 
	.B1(\ram[2][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n443));
   AO22CHD U2042 (.O(n617), 
	.B2(n30), 
	.B1(\ram[2][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n443));
   AO22CHD U2043 (.O(n618), 
	.B2(n30), 
	.B1(\ram[2][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n443));
   AO22CHD U2044 (.O(n619), 
	.B2(n30), 
	.B1(\ram[2][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n443));
   AO22CHD U2045 (.O(n620), 
	.B2(n30), 
	.B1(\ram[2][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n443));
   AO22CHD U2046 (.O(n621), 
	.B2(n30), 
	.B1(\ram[2][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n443));
   AO22CHD U2047 (.O(n622), 
	.B2(n30), 
	.B1(\ram[2][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n443));
   AO22CHD U2048 (.O(n623), 
	.B2(n30), 
	.B1(\ram[2][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n443));
   AO22CHD U2049 (.O(n624), 
	.B2(n30), 
	.B1(\ram[2][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n443));
   AO22CHD U2050 (.O(n625), 
	.B2(n30), 
	.B1(\ram[2][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n443));
   AO22CHD U2051 (.O(n626), 
	.B2(n30), 
	.B1(\ram[2][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n443));
   AO22CHD U2052 (.O(n627), 
	.B2(n30), 
	.B1(\ram[2][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n443));
   AO22CHD U2053 (.O(n628), 
	.B2(n30), 
	.B1(\ram[2][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n443));
   AO22CHD U2054 (.O(n629), 
	.B2(n30), 
	.B1(\ram[2][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n443));
   AO22CHD U2055 (.O(n630), 
	.B2(n33), 
	.B1(\ram[3][0] ), 
	.A2(n6), 
	.A1(n444));
   AO22CHD U2056 (.O(n631), 
	.B2(n33), 
	.B1(\ram[3][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n444));
   AO22CHD U2057 (.O(n632), 
	.B2(n33), 
	.B1(\ram[3][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n444));
   AO22CHD U2058 (.O(n633), 
	.B2(n33), 
	.B1(\ram[3][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n444));
   AO22CHD U2059 (.O(n634), 
	.B2(n33), 
	.B1(\ram[3][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n444));
   AO22CHD U2060 (.O(n635), 
	.B2(n33), 
	.B1(\ram[3][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n444));
   AO22CHD U2061 (.O(n636), 
	.B2(n33), 
	.B1(\ram[3][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n444));
   AO22CHD U2062 (.O(n637), 
	.B2(n33), 
	.B1(\ram[3][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n444));
   AO22CHD U2063 (.O(n638), 
	.B2(n33), 
	.B1(\ram[3][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n444));
   AO22CHD U2064 (.O(n639), 
	.B2(n33), 
	.B1(\ram[3][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n444));
   AO22CHD U2065 (.O(n640), 
	.B2(n33), 
	.B1(\ram[3][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n444));
   AO22CHD U2066 (.O(n641), 
	.B2(n33), 
	.B1(\ram[3][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n444));
   AO22CHD U2067 (.O(n642), 
	.B2(n33), 
	.B1(\ram[3][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n444));
   AO22CHD U2068 (.O(n643), 
	.B2(n33), 
	.B1(\ram[3][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n444));
   AO22CHD U2069 (.O(n644), 
	.B2(n33), 
	.B1(\ram[3][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n444));
   AO22CHD U2070 (.O(n645), 
	.B2(n33), 
	.B1(\ram[3][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n444));
   AO22CHD U2071 (.O(n646), 
	.B2(n36), 
	.B1(\ram[4][0] ), 
	.A2(n6), 
	.A1(n446));
   AO22CHD U2072 (.O(n647), 
	.B2(n36), 
	.B1(\ram[4][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n446));
   AO22CHD U2073 (.O(n648), 
	.B2(n36), 
	.B1(\ram[4][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n446));
   AO22CHD U2074 (.O(n649), 
	.B2(n36), 
	.B1(\ram[4][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n446));
   AO22CHD U2075 (.O(n650), 
	.B2(n36), 
	.B1(\ram[4][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n446));
   AO22CHD U2076 (.O(n651), 
	.B2(n36), 
	.B1(\ram[4][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n446));
   AO22CHD U2077 (.O(n652), 
	.B2(n36), 
	.B1(\ram[4][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n446));
   AO22CHD U2078 (.O(n653), 
	.B2(n36), 
	.B1(\ram[4][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n446));
   AO22CHD U2079 (.O(n654), 
	.B2(n36), 
	.B1(\ram[4][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n446));
   AO22CHD U2080 (.O(n655), 
	.B2(n36), 
	.B1(\ram[4][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n446));
   AO22CHD U2081 (.O(n656), 
	.B2(n36), 
	.B1(\ram[4][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n446));
   AO22CHD U2082 (.O(n657), 
	.B2(n36), 
	.B1(\ram[4][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n446));
   AO22CHD U2083 (.O(n658), 
	.B2(n36), 
	.B1(\ram[4][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n446));
   AO22CHD U2084 (.O(n659), 
	.B2(n36), 
	.B1(\ram[4][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n446));
   AO22CHD U2085 (.O(n660), 
	.B2(n36), 
	.B1(\ram[4][14] ), 
	.A2(n22), 
	.A1(n446));
   AO22CHD U2086 (.O(n661), 
	.B2(n36), 
	.B1(\ram[4][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n446));
   AO22CHD U2087 (.O(n662), 
	.B2(n39), 
	.B1(\ram[5][0] ), 
	.A2(n6), 
	.A1(n448));
   AO22CHD U2088 (.O(n663), 
	.B2(n39), 
	.B1(\ram[5][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n448));
   AO22CHD U2089 (.O(n664), 
	.B2(n39), 
	.B1(\ram[5][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n448));
   AO22CHD U2090 (.O(n665), 
	.B2(n39), 
	.B1(\ram[5][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n448));
   AO22CHD U2091 (.O(n666), 
	.B2(n39), 
	.B1(\ram[5][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n448));
   AO22CHD U2092 (.O(n667), 
	.B2(n39), 
	.B1(\ram[5][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n448));
   AO22CHD U2093 (.O(n668), 
	.B2(n39), 
	.B1(\ram[5][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n448));
   AO22CHD U2094 (.O(n669), 
	.B2(n39), 
	.B1(\ram[5][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n448));
   AO22CHD U2095 (.O(n670), 
	.B2(n39), 
	.B1(\ram[5][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n448));
   AO22CHD U2096 (.O(n671), 
	.B2(n39), 
	.B1(\ram[5][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n448));
   AO22CHD U2097 (.O(n672), 
	.B2(n39), 
	.B1(\ram[5][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n448));
   AO22CHD U2098 (.O(n673), 
	.B2(n39), 
	.B1(\ram[5][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n448));
   AO22CHD U2099 (.O(n674), 
	.B2(n39), 
	.B1(\ram[5][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n448));
   AO22CHD U2100 (.O(n675), 
	.B2(n39), 
	.B1(\ram[5][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n448));
   AO22CHD U2101 (.O(n676), 
	.B2(n39), 
	.B1(\ram[5][14] ), 
	.A2(n22), 
	.A1(n448));
   AO22CHD U2102 (.O(n677), 
	.B2(n39), 
	.B1(\ram[5][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n448));
   AO22CHD U2103 (.O(n678), 
	.B2(n42), 
	.B1(\ram[6][0] ), 
	.A2(n6), 
	.A1(n450));
   AO22CHD U2104 (.O(n679), 
	.B2(n42), 
	.B1(\ram[6][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n450));
   AO22CHD U2105 (.O(n680), 
	.B2(n42), 
	.B1(\ram[6][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n450));
   AO22CHD U2106 (.O(n681), 
	.B2(n42), 
	.B1(\ram[6][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n450));
   AO22CHD U2107 (.O(n682), 
	.B2(n42), 
	.B1(\ram[6][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n450));
   AO22CHD U2108 (.O(n683), 
	.B2(n42), 
	.B1(\ram[6][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n450));
   AO22CHD U2109 (.O(n684), 
	.B2(n42), 
	.B1(\ram[6][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n450));
   AO22CHD U2110 (.O(n685), 
	.B2(n42), 
	.B1(\ram[6][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n450));
   AO22CHD U2111 (.O(n686), 
	.B2(n42), 
	.B1(\ram[6][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n450));
   AO22CHD U2112 (.O(n687), 
	.B2(n42), 
	.B1(\ram[6][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n450));
   AO22CHD U2113 (.O(n688), 
	.B2(n42), 
	.B1(\ram[6][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n450));
   AO22CHD U2114 (.O(n689), 
	.B2(n42), 
	.B1(\ram[6][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n450));
   AO22CHD U2115 (.O(n690), 
	.B2(n42), 
	.B1(\ram[6][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n450));
   AO22CHD U2116 (.O(n691), 
	.B2(n42), 
	.B1(\ram[6][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n450));
   AO22CHD U2117 (.O(n692), 
	.B2(n42), 
	.B1(\ram[6][14] ), 
	.A2(n22), 
	.A1(n450));
   AO22CHD U2118 (.O(n693), 
	.B2(n42), 
	.B1(\ram[6][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n450));
   AO22CHD U2119 (.O(n694), 
	.B2(n45), 
	.B1(\ram[7][0] ), 
	.A2(n6), 
	.A1(n452));
   AO22CHD U2120 (.O(n695), 
	.B2(n45), 
	.B1(\ram[7][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n452));
   AO22CHD U2121 (.O(n696), 
	.B2(n45), 
	.B1(\ram[7][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n452));
   AO22CHD U2122 (.O(n697), 
	.B2(n45), 
	.B1(\ram[7][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n452));
   AO22CHD U2123 (.O(n698), 
	.B2(n45), 
	.B1(\ram[7][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n452));
   AO22CHD U2124 (.O(n699), 
	.B2(n45), 
	.B1(\ram[7][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n452));
   AO22CHD U2125 (.O(n700), 
	.B2(n45), 
	.B1(\ram[7][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n452));
   AO22CHD U2126 (.O(n701), 
	.B2(n45), 
	.B1(\ram[7][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n452));
   AO22CHD U2127 (.O(n702), 
	.B2(n45), 
	.B1(\ram[7][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n452));
   AO22CHD U2128 (.O(n703), 
	.B2(n45), 
	.B1(\ram[7][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n452));
   AO22CHD U2129 (.O(n704), 
	.B2(n45), 
	.B1(\ram[7][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n452));
   AO22CHD U2130 (.O(n705), 
	.B2(n45), 
	.B1(\ram[7][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n452));
   AO22CHD U2131 (.O(n706), 
	.B2(n45), 
	.B1(\ram[7][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n452));
   AO22CHD U2132 (.O(n707), 
	.B2(n45), 
	.B1(\ram[7][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n452));
   AO22CHD U2133 (.O(n708), 
	.B2(n45), 
	.B1(\ram[7][14] ), 
	.A2(n22), 
	.A1(n452));
   AO22CHD U2134 (.O(n709), 
	.B2(n45), 
	.B1(\ram[7][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n452));
   AO22CHD U2135 (.O(n710), 
	.B2(n48), 
	.B1(\ram[8][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n454));
   AO22CHD U2136 (.O(n711), 
	.B2(n48), 
	.B1(\ram[8][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n454));
   AO22CHD U2137 (.O(n712), 
	.B2(n48), 
	.B1(\ram[8][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n454));
   AO22CHD U2138 (.O(n713), 
	.B2(n48), 
	.B1(\ram[8][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n454));
   AO22CHD U2139 (.O(n714), 
	.B2(n48), 
	.B1(\ram[8][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n454));
   AO22CHD U2140 (.O(n715), 
	.B2(n48), 
	.B1(\ram[8][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n454));
   AO22CHD U2141 (.O(n716), 
	.B2(n48), 
	.B1(\ram[8][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n454));
   AO22CHD U2142 (.O(n717), 
	.B2(n48), 
	.B1(\ram[8][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n454));
   AO22CHD U2143 (.O(n718), 
	.B2(n48), 
	.B1(\ram[8][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n454));
   AO22CHD U2144 (.O(n719), 
	.B2(n48), 
	.B1(\ram[8][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n454));
   AO22CHD U2145 (.O(n720), 
	.B2(n48), 
	.B1(\ram[8][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n454));
   AO22CHD U2146 (.O(n721), 
	.B2(n48), 
	.B1(\ram[8][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n454));
   AO22CHD U2147 (.O(n722), 
	.B2(n48), 
	.B1(\ram[8][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n454));
   AO22CHD U2148 (.O(n723), 
	.B2(n48), 
	.B1(\ram[8][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n454));
   AO22CHD U2149 (.O(n724), 
	.B2(n48), 
	.B1(\ram[8][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n454));
   AO22CHD U2150 (.O(n725), 
	.B2(n48), 
	.B1(\ram[8][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n454));
   AO22CHD U2151 (.O(n726), 
	.B2(n51), 
	.B1(\ram[9][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n456));
   AO22CHD U2152 (.O(n727), 
	.B2(n51), 
	.B1(\ram[9][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n456));
   AO22CHD U2153 (.O(n728), 
	.B2(n51), 
	.B1(\ram[9][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n456));
   AO22CHD U2154 (.O(n729), 
	.B2(n51), 
	.B1(\ram[9][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n456));
   AO22CHD U2155 (.O(n730), 
	.B2(n51), 
	.B1(\ram[9][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n456));
   AO22CHD U2156 (.O(n731), 
	.B2(n51), 
	.B1(\ram[9][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n456));
   AO22CHD U2157 (.O(n732), 
	.B2(n51), 
	.B1(\ram[9][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n456));
   AO22CHD U2158 (.O(n733), 
	.B2(n51), 
	.B1(\ram[9][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n456));
   AO22CHD U2159 (.O(n734), 
	.B2(n51), 
	.B1(\ram[9][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n456));
   AO22CHD U2160 (.O(n735), 
	.B2(n51), 
	.B1(\ram[9][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n456));
   AO22CHD U2161 (.O(n736), 
	.B2(n51), 
	.B1(\ram[9][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n456));
   AO22CHD U2162 (.O(n737), 
	.B2(n51), 
	.B1(\ram[9][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n456));
   AO22CHD U2163 (.O(n738), 
	.B2(n51), 
	.B1(\ram[9][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n456));
   AO22CHD U2164 (.O(n739), 
	.B2(n51), 
	.B1(\ram[9][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n456));
   AO22CHD U2165 (.O(n740), 
	.B2(n51), 
	.B1(\ram[9][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n456));
   AO22CHD U2166 (.O(n741), 
	.B2(n51), 
	.B1(\ram[9][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n456));
   AO22CHD U2167 (.O(n742), 
	.B2(n54), 
	.B1(\ram[10][0] ), 
	.A2(n6), 
	.A1(n458));
   AO22CHD U2168 (.O(n743), 
	.B2(n54), 
	.B1(\ram[10][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n458));
   AO22CHD U2169 (.O(n744), 
	.B2(n54), 
	.B1(\ram[10][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n458));
   AO22CHD U2170 (.O(n745), 
	.B2(n54), 
	.B1(\ram[10][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n458));
   AO22CHD U2171 (.O(n746), 
	.B2(n54), 
	.B1(\ram[10][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n458));
   AO22CHD U2172 (.O(n747), 
	.B2(n54), 
	.B1(\ram[10][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n458));
   AO22CHD U2173 (.O(n748), 
	.B2(n54), 
	.B1(\ram[10][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n458));
   AO22CHD U2174 (.O(n749), 
	.B2(n54), 
	.B1(\ram[10][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n458));
   AO22CHD U2175 (.O(n750), 
	.B2(n54), 
	.B1(\ram[10][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n458));
   AO22CHD U2176 (.O(n751), 
	.B2(n54), 
	.B1(\ram[10][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n458));
   AO22CHD U2177 (.O(n752), 
	.B2(n54), 
	.B1(\ram[10][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n458));
   AO22CHD U2178 (.O(n753), 
	.B2(n54), 
	.B1(\ram[10][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n458));
   AO22CHD U2179 (.O(n754), 
	.B2(n54), 
	.B1(\ram[10][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n458));
   AO22CHD U2180 (.O(n755), 
	.B2(n54), 
	.B1(\ram[10][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n458));
   AO22CHD U2181 (.O(n756), 
	.B2(n54), 
	.B1(\ram[10][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n458));
   AO22CHD U2182 (.O(n757), 
	.B2(n54), 
	.B1(\ram[10][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n458));
   AO22CHD U2183 (.O(n758), 
	.B2(n57), 
	.B1(\ram[11][0] ), 
	.A2(n6), 
	.A1(n460));
   AO22CHD U2184 (.O(n759), 
	.B2(n57), 
	.B1(\ram[11][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n460));
   AO22CHD U2185 (.O(n760), 
	.B2(n57), 
	.B1(\ram[11][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n460));
   AO22CHD U2186 (.O(n761), 
	.B2(n57), 
	.B1(\ram[11][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n460));
   AO22CHD U2187 (.O(n762), 
	.B2(n57), 
	.B1(\ram[11][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n460));
   AO22CHD U2188 (.O(n763), 
	.B2(n57), 
	.B1(\ram[11][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n460));
   AO22CHD U2189 (.O(n764), 
	.B2(n57), 
	.B1(\ram[11][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n460));
   AO22CHD U2190 (.O(n765), 
	.B2(n57), 
	.B1(\ram[11][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n460));
   AO22CHD U2191 (.O(n766), 
	.B2(n57), 
	.B1(\ram[11][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n460));
   AO22CHD U2192 (.O(n767), 
	.B2(n57), 
	.B1(\ram[11][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n460));
   AO22CHD U2193 (.O(n768), 
	.B2(n57), 
	.B1(\ram[11][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n460));
   AO22CHD U2194 (.O(n769), 
	.B2(n57), 
	.B1(\ram[11][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n460));
   AO22CHD U2195 (.O(n770), 
	.B2(n57), 
	.B1(\ram[11][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n460));
   AO22CHD U2196 (.O(n771), 
	.B2(n57), 
	.B1(\ram[11][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n460));
   AO22CHD U2197 (.O(n772), 
	.B2(n57), 
	.B1(\ram[11][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n460));
   AO22CHD U2198 (.O(n773), 
	.B2(n57), 
	.B1(\ram[11][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n460));
   AO22CHD U2199 (.O(n774), 
	.B2(n60), 
	.B1(\ram[12][0] ), 
	.A2(n6), 
	.A1(n462));
   AO22CHD U2200 (.O(n775), 
	.B2(n60), 
	.B1(\ram[12][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n462));
   AO22CHD U2201 (.O(n776), 
	.B2(n60), 
	.B1(\ram[12][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n462));
   AO22CHD U2202 (.O(n777), 
	.B2(n60), 
	.B1(\ram[12][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n462));
   AO22CHD U2203 (.O(n778), 
	.B2(n60), 
	.B1(\ram[12][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n462));
   AO22CHD U2204 (.O(n779), 
	.B2(n60), 
	.B1(\ram[12][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n462));
   AO22CHD U2205 (.O(n780), 
	.B2(n60), 
	.B1(\ram[12][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n462));
   AO22CHD U2206 (.O(n781), 
	.B2(n60), 
	.B1(\ram[12][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n462));
   AO22CHD U2207 (.O(n782), 
	.B2(n60), 
	.B1(\ram[12][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n462));
   AO22CHD U2208 (.O(n783), 
	.B2(n60), 
	.B1(\ram[12][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n462));
   AO22CHD U2209 (.O(n784), 
	.B2(n60), 
	.B1(\ram[12][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n462));
   AO22CHD U2210 (.O(n785), 
	.B2(n60), 
	.B1(\ram[12][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n462));
   AO22CHD U2211 (.O(n786), 
	.B2(n60), 
	.B1(\ram[12][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n462));
   AO22CHD U2212 (.O(n787), 
	.B2(n60), 
	.B1(\ram[12][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n462));
   AO22CHD U2213 (.O(n788), 
	.B2(n60), 
	.B1(\ram[12][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n462));
   AO22CHD U2214 (.O(n789), 
	.B2(n60), 
	.B1(\ram[12][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n462));
   AO22CHD U2215 (.O(n790), 
	.B2(n63), 
	.B1(\ram[13][0] ), 
	.A2(n6), 
	.A1(n464));
   AO22CHD U2216 (.O(n791), 
	.B2(n63), 
	.B1(\ram[13][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n464));
   AO22CHD U2217 (.O(n792), 
	.B2(n63), 
	.B1(\ram[13][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n464));
   AO22CHD U2218 (.O(n793), 
	.B2(n63), 
	.B1(\ram[13][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n464));
   AO22CHD U2219 (.O(n794), 
	.B2(n63), 
	.B1(\ram[13][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n464));
   AO22CHD U2220 (.O(n795), 
	.B2(n63), 
	.B1(\ram[13][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n464));
   AO22CHD U2221 (.O(n796), 
	.B2(n63), 
	.B1(\ram[13][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n464));
   AO22CHD U2222 (.O(n797), 
	.B2(n63), 
	.B1(\ram[13][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n464));
   AO22CHD U2223 (.O(n798), 
	.B2(n63), 
	.B1(\ram[13][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n464));
   AO22CHD U2224 (.O(n799), 
	.B2(n63), 
	.B1(\ram[13][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n464));
   AO22CHD U2225 (.O(n800), 
	.B2(n63), 
	.B1(\ram[13][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n464));
   AO22CHD U2226 (.O(n801), 
	.B2(n63), 
	.B1(\ram[13][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n464));
   AO22CHD U2227 (.O(n802), 
	.B2(n63), 
	.B1(\ram[13][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n464));
   AO22CHD U2228 (.O(n803), 
	.B2(n63), 
	.B1(\ram[13][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n464));
   AO22CHD U2229 (.O(n804), 
	.B2(n63), 
	.B1(\ram[13][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n464));
   AO22CHD U2230 (.O(n805), 
	.B2(n63), 
	.B1(\ram[13][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n464));
   AO22CHD U2231 (.O(n806), 
	.B2(n66), 
	.B1(\ram[14][0] ), 
	.A2(n6), 
	.A1(n466));
   AO22CHD U2232 (.O(n807), 
	.B2(n66), 
	.B1(\ram[14][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n466));
   AO22CHD U2233 (.O(n808), 
	.B2(n66), 
	.B1(\ram[14][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n466));
   AO22CHD U2234 (.O(n809), 
	.B2(n66), 
	.B1(\ram[14][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n466));
   AO22CHD U2235 (.O(n810), 
	.B2(n66), 
	.B1(\ram[14][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n466));
   AO22CHD U2236 (.O(n811), 
	.B2(n66), 
	.B1(\ram[14][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n466));
   AO22CHD U2237 (.O(n812), 
	.B2(n66), 
	.B1(\ram[14][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n466));
   AO22CHD U2238 (.O(n813), 
	.B2(n66), 
	.B1(\ram[14][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n466));
   AO22CHD U2239 (.O(n814), 
	.B2(n66), 
	.B1(\ram[14][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n466));
   AO22CHD U2240 (.O(n815), 
	.B2(n66), 
	.B1(\ram[14][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n466));
   AO22CHD U2241 (.O(n816), 
	.B2(n66), 
	.B1(\ram[14][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n466));
   AO22CHD U2242 (.O(n817), 
	.B2(n66), 
	.B1(\ram[14][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n466));
   AO22CHD U2243 (.O(n818), 
	.B2(n66), 
	.B1(\ram[14][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n466));
   AO22CHD U2244 (.O(n819), 
	.B2(n66), 
	.B1(\ram[14][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n466));
   AO22CHD U2245 (.O(n820), 
	.B2(n66), 
	.B1(\ram[14][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n466));
   AO22CHD U2246 (.O(n821), 
	.B2(n66), 
	.B1(\ram[14][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n466));
   AO22CHD U2247 (.O(n822), 
	.B2(n69), 
	.B1(\ram[15][0] ), 
	.A2(n6), 
	.A1(n468));
   AO22CHD U2248 (.O(n823), 
	.B2(n69), 
	.B1(\ram[15][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n468));
   AO22CHD U2249 (.O(n824), 
	.B2(n69), 
	.B1(\ram[15][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n468));
   AO22CHD U2250 (.O(n825), 
	.B2(n69), 
	.B1(\ram[15][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n468));
   AO22CHD U2251 (.O(n826), 
	.B2(n69), 
	.B1(\ram[15][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n468));
   AO22CHD U2252 (.O(n827), 
	.B2(n69), 
	.B1(\ram[15][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n468));
   AO22CHD U2253 (.O(n828), 
	.B2(n69), 
	.B1(\ram[15][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n468));
   AO22CHD U2254 (.O(n829), 
	.B2(n69), 
	.B1(\ram[15][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n468));
   AO22CHD U2255 (.O(n830), 
	.B2(n69), 
	.B1(\ram[15][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n468));
   AO22CHD U2256 (.O(n831), 
	.B2(n69), 
	.B1(\ram[15][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n468));
   AO22CHD U2257 (.O(n832), 
	.B2(n69), 
	.B1(\ram[15][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n468));
   AO22CHD U2258 (.O(n833), 
	.B2(n69), 
	.B1(\ram[15][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n468));
   AO22CHD U2259 (.O(n834), 
	.B2(n69), 
	.B1(\ram[15][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n468));
   AO22CHD U2260 (.O(n835), 
	.B2(n69), 
	.B1(\ram[15][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n468));
   AO22CHD U2261 (.O(n836), 
	.B2(n69), 
	.B1(\ram[15][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n468));
   AO22CHD U2262 (.O(n837), 
	.B2(n69), 
	.B1(\ram[15][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n468));
   AO22CHD U2263 (.O(n838), 
	.B2(n74), 
	.B1(\ram[16][0] ), 
	.A2(n6), 
	.A1(n470));
   AO22CHD U2264 (.O(n839), 
	.B2(n74), 
	.B1(\ram[16][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n470));
   AO22CHD U2265 (.O(n840), 
	.B2(n74), 
	.B1(\ram[16][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n470));
   AO22CHD U2266 (.O(n841), 
	.B2(n74), 
	.B1(\ram[16][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n470));
   AO22CHD U2267 (.O(n842), 
	.B2(n74), 
	.B1(\ram[16][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n470));
   AO22CHD U2268 (.O(n843), 
	.B2(n74), 
	.B1(\ram[16][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n470));
   AO22CHD U2269 (.O(n844), 
	.B2(n74), 
	.B1(\ram[16][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n470));
   AO22CHD U2270 (.O(n845), 
	.B2(n74), 
	.B1(\ram[16][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n470));
   AO22CHD U2271 (.O(n846), 
	.B2(n74), 
	.B1(\ram[16][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n470));
   AO22CHD U2272 (.O(n847), 
	.B2(n74), 
	.B1(\ram[16][9] ), 
	.A2(n17), 
	.A1(n470));
   AO22CHD U2273 (.O(n848), 
	.B2(n74), 
	.B1(\ram[16][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n470));
   AO22CHD U2274 (.O(n849), 
	.B2(n74), 
	.B1(\ram[16][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n470));
   AO22CHD U2275 (.O(n850), 
	.B2(n74), 
	.B1(\ram[16][12] ), 
	.A2(n20), 
	.A1(n470));
   AO22CHD U2276 (.O(n851), 
	.B2(n74), 
	.B1(\ram[16][13] ), 
	.A2(n21), 
	.A1(n470));
   AO22CHD U2277 (.O(n852), 
	.B2(n74), 
	.B1(\ram[16][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n470));
   AO22CHD U2278 (.O(n853), 
	.B2(n74), 
	.B1(\ram[16][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n470));
   AO22CHD U2279 (.O(n854), 
	.B2(n77), 
	.B1(\ram[17][0] ), 
	.A2(n6), 
	.A1(n472));
   AO22CHD U2280 (.O(n855), 
	.B2(n77), 
	.B1(\ram[17][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n472));
   AO22CHD U2281 (.O(n856), 
	.B2(n77), 
	.B1(\ram[17][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n472));
   AO22CHD U2282 (.O(n857), 
	.B2(n77), 
	.B1(\ram[17][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n472));
   AO22CHD U2283 (.O(n858), 
	.B2(n77), 
	.B1(\ram[17][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n472));
   AO22CHD U2284 (.O(n859), 
	.B2(n77), 
	.B1(\ram[17][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n472));
   AO22CHD U2285 (.O(n860), 
	.B2(n77), 
	.B1(\ram[17][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n472));
   AO22CHD U2286 (.O(n861), 
	.B2(n77), 
	.B1(\ram[17][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n472));
   AO22CHD U2287 (.O(n862), 
	.B2(n77), 
	.B1(\ram[17][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n472));
   AO22CHD U2288 (.O(n863), 
	.B2(n77), 
	.B1(\ram[17][9] ), 
	.A2(n17), 
	.A1(n472));
   AO22CHD U2289 (.O(n864), 
	.B2(n77), 
	.B1(\ram[17][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n472));
   AO22CHD U2290 (.O(n865), 
	.B2(n77), 
	.B1(\ram[17][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n472));
   AO22CHD U2291 (.O(n866), 
	.B2(n77), 
	.B1(\ram[17][12] ), 
	.A2(n20), 
	.A1(n472));
   AO22CHD U2292 (.O(n867), 
	.B2(n77), 
	.B1(\ram[17][13] ), 
	.A2(n21), 
	.A1(n472));
   AO22CHD U2293 (.O(n868), 
	.B2(n77), 
	.B1(\ram[17][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n472));
   AO22CHD U2294 (.O(n869), 
	.B2(n77), 
	.B1(\ram[17][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n472));
   AO22CHD U2295 (.O(n870), 
	.B2(n79), 
	.B1(\ram[18][0] ), 
	.A2(n6), 
	.A1(n475));
   AO22CHD U2296 (.O(n871), 
	.B2(n79), 
	.B1(\ram[18][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n475));
   AO22CHD U2297 (.O(n872), 
	.B2(n79), 
	.B1(\ram[18][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n475));
   AO22CHD U2298 (.O(n873), 
	.B2(n79), 
	.B1(\ram[18][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n475));
   AO22CHD U2299 (.O(n874), 
	.B2(n79), 
	.B1(\ram[18][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n475));
   AO22CHD U2300 (.O(n875), 
	.B2(n79), 
	.B1(\ram[18][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n475));
   AO22CHD U2301 (.O(n876), 
	.B2(n79), 
	.B1(\ram[18][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n475));
   AO22CHD U2302 (.O(n877), 
	.B2(n79), 
	.B1(\ram[18][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n475));
   AO22CHD U2303 (.O(n878), 
	.B2(n79), 
	.B1(\ram[18][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n475));
   AO22CHD U2304 (.O(n879), 
	.B2(n79), 
	.B1(\ram[18][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n475));
   AO22CHD U2305 (.O(n880), 
	.B2(n79), 
	.B1(\ram[18][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n475));
   AO22CHD U2306 (.O(n881), 
	.B2(n79), 
	.B1(\ram[18][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n475));
   AO22CHD U2307 (.O(n882), 
	.B2(n79), 
	.B1(\ram[18][12] ), 
	.A2(n20), 
	.A1(n475));
   AO22CHD U2308 (.O(n883), 
	.B2(n79), 
	.B1(\ram[18][13] ), 
	.A2(n21), 
	.A1(n475));
   AO22CHD U2309 (.O(n884), 
	.B2(n79), 
	.B1(\ram[18][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n475));
   AO22CHD U2310 (.O(n885), 
	.B2(n79), 
	.B1(\ram[18][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n475));
   AO22CHD U2311 (.O(n886), 
	.B2(n81), 
	.B1(\ram[19][0] ), 
	.A2(n6), 
	.A1(n477));
   AO22CHD U2312 (.O(n887), 
	.B2(n81), 
	.B1(\ram[19][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n477));
   AO22CHD U2313 (.O(n888), 
	.B2(n81), 
	.B1(\ram[19][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n477));
   AO22CHD U2314 (.O(n889), 
	.B2(n81), 
	.B1(\ram[19][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n477));
   AO22CHD U2315 (.O(n890), 
	.B2(n81), 
	.B1(\ram[19][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n477));
   AO22CHD U2316 (.O(n891), 
	.B2(n81), 
	.B1(\ram[19][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n477));
   AO22CHD U2317 (.O(n892), 
	.B2(n81), 
	.B1(\ram[19][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n477));
   AO22CHD U2318 (.O(n893), 
	.B2(n81), 
	.B1(\ram[19][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n477));
   AO22CHD U2319 (.O(n894), 
	.B2(n81), 
	.B1(\ram[19][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n477));
   AO22CHD U2320 (.O(n895), 
	.B2(n81), 
	.B1(\ram[19][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n477));
   AO22CHD U2321 (.O(n896), 
	.B2(n81), 
	.B1(\ram[19][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n477));
   AO22CHD U2322 (.O(n897), 
	.B2(n81), 
	.B1(\ram[19][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n477));
   AO22CHD U2323 (.O(n898), 
	.B2(n81), 
	.B1(\ram[19][12] ), 
	.A2(n20), 
	.A1(n477));
   AO22CHD U2324 (.O(n899), 
	.B2(n81), 
	.B1(\ram[19][13] ), 
	.A2(n21), 
	.A1(n477));
   AO22CHD U2325 (.O(n900), 
	.B2(n81), 
	.B1(\ram[19][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n477));
   AO22CHD U2326 (.O(n901), 
	.B2(n81), 
	.B1(\ram[19][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n477));
   AO22CHD U2327 (.O(n902), 
	.B2(n83), 
	.B1(\ram[20][0] ), 
	.A2(n6), 
	.A1(n478));
   AO22CHD U2328 (.O(n903), 
	.B2(n83), 
	.B1(\ram[20][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n478));
   AO22CHD U2329 (.O(n904), 
	.B2(n83), 
	.B1(\ram[20][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n478));
   AO22CHD U2330 (.O(n905), 
	.B2(n83), 
	.B1(\ram[20][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n478));
   AO22CHD U2331 (.O(n906), 
	.B2(n83), 
	.B1(\ram[20][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n478));
   AO22CHD U2332 (.O(n907), 
	.B2(n83), 
	.B1(\ram[20][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n478));
   AO22CHD U2333 (.O(n908), 
	.B2(n83), 
	.B1(\ram[20][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n478));
   AO22CHD U2334 (.O(n909), 
	.B2(n83), 
	.B1(\ram[20][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n478));
   AO22CHD U2335 (.O(n910), 
	.B2(n83), 
	.B1(\ram[20][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n478));
   AO22CHD U2336 (.O(n911), 
	.B2(n83), 
	.B1(\ram[20][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n478));
   AO22CHD U2337 (.O(n912), 
	.B2(n83), 
	.B1(\ram[20][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n478));
   AO22CHD U2338 (.O(n913), 
	.B2(n83), 
	.B1(\ram[20][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n478));
   AO22CHD U2339 (.O(n914), 
	.B2(n83), 
	.B1(\ram[20][12] ), 
	.A2(n20), 
	.A1(n478));
   AO22CHD U2340 (.O(n915), 
	.B2(n83), 
	.B1(\ram[20][13] ), 
	.A2(n21), 
	.A1(n478));
   AO22CHD U2341 (.O(n916), 
	.B2(n83), 
	.B1(\ram[20][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n478));
   AO22CHD U2342 (.O(n917), 
	.B2(n83), 
	.B1(\ram[20][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n478));
   AO22CHD U2343 (.O(n918), 
	.B2(n85), 
	.B1(\ram[21][0] ), 
	.A2(n6), 
	.A1(n480));
   AO22CHD U2344 (.O(n919), 
	.B2(n85), 
	.B1(\ram[21][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n480));
   AO22CHD U2345 (.O(n920), 
	.B2(n85), 
	.B1(\ram[21][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n480));
   AO22CHD U2346 (.O(n921), 
	.B2(n85), 
	.B1(\ram[21][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n480));
   AO22CHD U2347 (.O(n922), 
	.B2(n85), 
	.B1(\ram[21][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n480));
   AO22CHD U2348 (.O(n923), 
	.B2(n85), 
	.B1(\ram[21][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n480));
   AO22CHD U2349 (.O(n924), 
	.B2(n85), 
	.B1(\ram[21][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n480));
   AO22CHD U2350 (.O(n925), 
	.B2(n85), 
	.B1(\ram[21][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n480));
   AO22CHD U2351 (.O(n926), 
	.B2(n85), 
	.B1(\ram[21][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n480));
   AO22CHD U2352 (.O(n927), 
	.B2(n85), 
	.B1(\ram[21][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n480));
   AO22CHD U2353 (.O(n928), 
	.B2(n85), 
	.B1(\ram[21][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n480));
   AO22CHD U2354 (.O(n929), 
	.B2(n85), 
	.B1(\ram[21][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n480));
   AO22CHD U2355 (.O(n930), 
	.B2(n85), 
	.B1(\ram[21][12] ), 
	.A2(n20), 
	.A1(n480));
   AO22CHD U2356 (.O(n931), 
	.B2(n85), 
	.B1(\ram[21][13] ), 
	.A2(n21), 
	.A1(n480));
   AO22CHD U2357 (.O(n932), 
	.B2(n85), 
	.B1(\ram[21][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n480));
   AO22CHD U2358 (.O(n933), 
	.B2(n85), 
	.B1(\ram[21][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n480));
   AO22CHD U2359 (.O(n934), 
	.B2(n87), 
	.B1(\ram[22][0] ), 
	.A2(n6), 
	.A1(n482));
   AO22CHD U2360 (.O(n935), 
	.B2(n87), 
	.B1(\ram[22][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n482));
   AO22CHD U2361 (.O(n936), 
	.B2(n87), 
	.B1(\ram[22][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n482));
   AO22CHD U2362 (.O(n937), 
	.B2(n87), 
	.B1(\ram[22][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n482));
   AO22CHD U2363 (.O(n938), 
	.B2(n87), 
	.B1(\ram[22][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n482));
   AO22CHD U2364 (.O(n939), 
	.B2(n87), 
	.B1(\ram[22][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n482));
   AO22CHD U2365 (.O(n940), 
	.B2(n87), 
	.B1(\ram[22][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n482));
   AO22CHD U2366 (.O(n941), 
	.B2(n87), 
	.B1(\ram[22][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n482));
   AO22CHD U2367 (.O(n942), 
	.B2(n87), 
	.B1(\ram[22][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n482));
   AO22CHD U2368 (.O(n943), 
	.B2(n87), 
	.B1(\ram[22][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n482));
   AO22CHD U2369 (.O(n944), 
	.B2(n87), 
	.B1(\ram[22][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n482));
   AO22CHD U2370 (.O(n945), 
	.B2(n87), 
	.B1(\ram[22][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n482));
   AO22CHD U2371 (.O(n946), 
	.B2(n87), 
	.B1(\ram[22][12] ), 
	.A2(n20), 
	.A1(n482));
   AO22CHD U2372 (.O(n947), 
	.B2(n87), 
	.B1(\ram[22][13] ), 
	.A2(n21), 
	.A1(n482));
   AO22CHD U2373 (.O(n948), 
	.B2(n87), 
	.B1(\ram[22][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n482));
   AO22CHD U2374 (.O(n949), 
	.B2(n87), 
	.B1(\ram[22][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n482));
   AO22CHD U2375 (.O(n950), 
	.B2(n89), 
	.B1(\ram[23][0] ), 
	.A2(n6), 
	.A1(n484));
   AO22CHD U2376 (.O(n951), 
	.B2(n89), 
	.B1(\ram[23][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n484));
   AO22CHD U2377 (.O(n952), 
	.B2(n89), 
	.B1(\ram[23][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n484));
   AO22CHD U2378 (.O(n953), 
	.B2(n89), 
	.B1(\ram[23][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n484));
   AO22CHD U2379 (.O(n954), 
	.B2(n89), 
	.B1(\ram[23][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n484));
   AO22CHD U2380 (.O(n955), 
	.B2(n89), 
	.B1(\ram[23][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n484));
   AO22CHD U2381 (.O(n956), 
	.B2(n89), 
	.B1(\ram[23][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n484));
   AO22CHD U2382 (.O(n957), 
	.B2(n89), 
	.B1(\ram[23][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n484));
   AO22CHD U2383 (.O(n958), 
	.B2(n89), 
	.B1(\ram[23][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n484));
   AO22CHD U2384 (.O(n959), 
	.B2(n89), 
	.B1(\ram[23][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n484));
   AO22CHD U2385 (.O(n960), 
	.B2(n89), 
	.B1(\ram[23][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n484));
   AO22CHD U2386 (.O(n961), 
	.B2(n89), 
	.B1(\ram[23][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n484));
   AO22CHD U2387 (.O(n962), 
	.B2(n89), 
	.B1(\ram[23][12] ), 
	.A2(n20), 
	.A1(n484));
   AO22CHD U2388 (.O(n963), 
	.B2(n89), 
	.B1(\ram[23][13] ), 
	.A2(n21), 
	.A1(n484));
   AO22CHD U2389 (.O(n964), 
	.B2(n89), 
	.B1(\ram[23][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n484));
   AO22CHD U2390 (.O(n965), 
	.B2(n89), 
	.B1(\ram[23][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n484));
   AO22CHD U2391 (.O(n966), 
	.B2(n91), 
	.B1(\ram[24][0] ), 
	.A2(n6), 
	.A1(n486));
   AO22CHD U2392 (.O(n967), 
	.B2(n91), 
	.B1(\ram[24][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n486));
   AO22CHD U2393 (.O(n968), 
	.B2(n91), 
	.B1(\ram[24][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n486));
   AO22CHD U2394 (.O(n969), 
	.B2(n91), 
	.B1(\ram[24][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n486));
   AO22CHD U2395 (.O(n970), 
	.B2(n91), 
	.B1(\ram[24][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n486));
   AO22CHD U2396 (.O(n971), 
	.B2(n91), 
	.B1(\ram[24][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n486));
   AO22CHD U2397 (.O(n972), 
	.B2(n91), 
	.B1(\ram[24][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n486));
   AO22CHD U2398 (.O(n973), 
	.B2(n91), 
	.B1(\ram[24][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n486));
   AO22CHD U2399 (.O(n974), 
	.B2(n91), 
	.B1(\ram[24][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n486));
   AO22CHD U2400 (.O(n975), 
	.B2(n91), 
	.B1(\ram[24][9] ), 
	.A2(n17), 
	.A1(n486));
   AO22CHD U2401 (.O(n976), 
	.B2(n91), 
	.B1(\ram[24][10] ), 
	.A2(n18), 
	.A1(n486));
   AO22CHD U2402 (.O(n977), 
	.B2(n91), 
	.B1(\ram[24][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n486));
   AO22CHD U2403 (.O(n978), 
	.B2(n91), 
	.B1(\ram[24][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n486));
   AO22CHD U2404 (.O(n979), 
	.B2(n91), 
	.B1(\ram[24][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n486));
   AO22CHD U2405 (.O(n980), 
	.B2(n91), 
	.B1(\ram[24][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n486));
   AO22CHD U2406 (.O(n981), 
	.B2(n91), 
	.B1(\ram[24][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n486));
   AO22CHD U2407 (.O(n982), 
	.B2(n93), 
	.B1(\ram[25][0] ), 
	.A2(n6), 
	.A1(n488));
   AO22CHD U2408 (.O(n983), 
	.B2(n93), 
	.B1(\ram[25][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n488));
   AO22CHD U2409 (.O(n984), 
	.B2(n93), 
	.B1(\ram[25][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n488));
   AO22CHD U2410 (.O(n985), 
	.B2(n93), 
	.B1(\ram[25][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n488));
   AO22CHD U2411 (.O(n986), 
	.B2(n93), 
	.B1(\ram[25][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n488));
   AO22CHD U2412 (.O(n987), 
	.B2(n93), 
	.B1(\ram[25][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n488));
   AO22CHD U2413 (.O(n988), 
	.B2(n93), 
	.B1(\ram[25][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n488));
   AO22CHD U2414 (.O(n989), 
	.B2(n93), 
	.B1(\ram[25][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n488));
   AO22CHD U2415 (.O(n990), 
	.B2(n93), 
	.B1(\ram[25][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n488));
   AO22CHD U2416 (.O(n991), 
	.B2(n93), 
	.B1(\ram[25][9] ), 
	.A2(n17), 
	.A1(n488));
   AO22CHD U2417 (.O(n992), 
	.B2(n93), 
	.B1(\ram[25][10] ), 
	.A2(n18), 
	.A1(n488));
   AO22CHD U2418 (.O(n993), 
	.B2(n93), 
	.B1(\ram[25][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n488));
   AO22CHD U2419 (.O(n994), 
	.B2(n93), 
	.B1(\ram[25][12] ), 
	.A2(n20), 
	.A1(n488));
   AO22CHD U2420 (.O(n995), 
	.B2(n93), 
	.B1(\ram[25][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n488));
   AO22CHD U2421 (.O(n996), 
	.B2(n93), 
	.B1(\ram[25][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n488));
   AO22CHD U2422 (.O(n997), 
	.B2(n93), 
	.B1(\ram[25][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n488));
   AO22CHD U2423 (.O(n998), 
	.B2(n95), 
	.B1(\ram[26][0] ), 
	.A2(n6), 
	.A1(n490));
   AO22CHD U2424 (.O(n999), 
	.B2(n95), 
	.B1(\ram[26][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n490));
   AO22CHD U2425 (.O(n1000), 
	.B2(n95), 
	.B1(\ram[26][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n490));
   AO22CHD U2426 (.O(n1001), 
	.B2(n95), 
	.B1(\ram[26][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n490));
   AO22CHD U2427 (.O(n1002), 
	.B2(n95), 
	.B1(\ram[26][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n490));
   AO22CHD U2428 (.O(n1003), 
	.B2(n95), 
	.B1(\ram[26][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n490));
   AO22CHD U2429 (.O(n1004), 
	.B2(n95), 
	.B1(\ram[26][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n490));
   AO22CHD U2430 (.O(n1005), 
	.B2(n95), 
	.B1(\ram[26][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n490));
   AO22CHD U2431 (.O(n1006), 
	.B2(n95), 
	.B1(\ram[26][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n490));
   AO22CHD U2432 (.O(n1007), 
	.B2(n95), 
	.B1(\ram[26][9] ), 
	.A2(n17), 
	.A1(n490));
   AO22CHD U2433 (.O(n1008), 
	.B2(n95), 
	.B1(\ram[26][10] ), 
	.A2(n18), 
	.A1(n490));
   AO22CHD U2434 (.O(n1009), 
	.B2(n95), 
	.B1(\ram[26][11] ), 
	.A2(n19), 
	.A1(n490));
   AO22CHD U2435 (.O(n1010), 
	.B2(n95), 
	.B1(\ram[26][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n490));
   AO22CHD U2436 (.O(n1011), 
	.B2(n95), 
	.B1(\ram[26][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n490));
   AO22CHD U2437 (.O(n1012), 
	.B2(n95), 
	.B1(\ram[26][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n490));
   AO22CHD U2438 (.O(n1013), 
	.B2(n95), 
	.B1(\ram[26][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n490));
   AO22CHD U2439 (.O(n1014), 
	.B2(n97), 
	.B1(\ram[27][0] ), 
	.A2(n6), 
	.A1(n492));
   AO22CHD U2440 (.O(n1015), 
	.B2(n97), 
	.B1(\ram[27][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n492));
   AO22CHD U2441 (.O(n1016), 
	.B2(n97), 
	.B1(\ram[27][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n492));
   AO22CHD U2442 (.O(n1017), 
	.B2(n97), 
	.B1(\ram[27][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n492));
   AO22CHD U2443 (.O(n1018), 
	.B2(n97), 
	.B1(\ram[27][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n492));
   AO22CHD U2444 (.O(n1019), 
	.B2(n97), 
	.B1(\ram[27][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n492));
   AO22CHD U2445 (.O(n1020), 
	.B2(n97), 
	.B1(\ram[27][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n492));
   AO22CHD U2446 (.O(n1021), 
	.B2(n97), 
	.B1(\ram[27][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n492));
   AO22CHD U2447 (.O(n1022), 
	.B2(n97), 
	.B1(\ram[27][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n492));
   AO22CHD U2448 (.O(n1023), 
	.B2(n97), 
	.B1(\ram[27][9] ), 
	.A2(n17), 
	.A1(n492));
   AO22CHD U2449 (.O(n1024), 
	.B2(n97), 
	.B1(\ram[27][10] ), 
	.A2(n18), 
	.A1(n492));
   AO22CHD U2450 (.O(n1025), 
	.B2(n97), 
	.B1(\ram[27][11] ), 
	.A2(n19), 
	.A1(n492));
   AO22CHD U2451 (.O(n1026), 
	.B2(n97), 
	.B1(\ram[27][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n492));
   AO22CHD U2452 (.O(n1027), 
	.B2(n97), 
	.B1(\ram[27][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n492));
   AO22CHD U2453 (.O(n1028), 
	.B2(n97), 
	.B1(\ram[27][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n492));
   AO22CHD U2454 (.O(n1029), 
	.B2(n97), 
	.B1(\ram[27][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n492));
   AO22CHD U2455 (.O(n1030), 
	.B2(n99), 
	.B1(\ram[28][0] ), 
	.A2(n6), 
	.A1(n494));
   AO22CHD U2456 (.O(n1031), 
	.B2(n99), 
	.B1(\ram[28][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n494));
   AO22CHD U2457 (.O(n1032), 
	.B2(n99), 
	.B1(\ram[28][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n494));
   AO22CHD U2458 (.O(n1033), 
	.B2(n99), 
	.B1(\ram[28][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n494));
   AO22CHD U2459 (.O(n1034), 
	.B2(n99), 
	.B1(\ram[28][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n494));
   AO22CHD U2460 (.O(n1035), 
	.B2(n99), 
	.B1(\ram[28][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n494));
   AO22CHD U2461 (.O(n1036), 
	.B2(n99), 
	.B1(\ram[28][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n494));
   AO22CHD U2462 (.O(n1037), 
	.B2(n99), 
	.B1(\ram[28][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n494));
   AO22CHD U2463 (.O(n1038), 
	.B2(n99), 
	.B1(\ram[28][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n494));
   AO22CHD U2464 (.O(n1039), 
	.B2(n99), 
	.B1(\ram[28][9] ), 
	.A2(n17), 
	.A1(n494));
   AO22CHD U2465 (.O(n1040), 
	.B2(n99), 
	.B1(\ram[28][10] ), 
	.A2(n18), 
	.A1(n494));
   AO22CHD U2466 (.O(n1041), 
	.B2(n99), 
	.B1(\ram[28][11] ), 
	.A2(n19), 
	.A1(n494));
   AO22CHD U2467 (.O(n1042), 
	.B2(n99), 
	.B1(\ram[28][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n494));
   AO22CHD U2468 (.O(n1043), 
	.B2(n99), 
	.B1(\ram[28][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n494));
   AO22CHD U2469 (.O(n1044), 
	.B2(n99), 
	.B1(\ram[28][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n494));
   AO22CHD U2470 (.O(n1045), 
	.B2(n99), 
	.B1(\ram[28][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n494));
   AO22CHD U2471 (.O(n1046), 
	.B2(n101), 
	.B1(\ram[29][0] ), 
	.A2(n6), 
	.A1(n496));
   AO22CHD U2472 (.O(n1047), 
	.B2(n101), 
	.B1(\ram[29][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n496));
   AO22CHD U2473 (.O(n1048), 
	.B2(n101), 
	.B1(\ram[29][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n496));
   AO22CHD U2474 (.O(n1049), 
	.B2(n101), 
	.B1(\ram[29][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n496));
   AO22CHD U2475 (.O(n1050), 
	.B2(n101), 
	.B1(\ram[29][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n496));
   AO22CHD U2476 (.O(n1051), 
	.B2(n101), 
	.B1(\ram[29][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n496));
   AO22CHD U2477 (.O(n1052), 
	.B2(n101), 
	.B1(\ram[29][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n496));
   AO22CHD U2478 (.O(n1053), 
	.B2(n101), 
	.B1(\ram[29][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n496));
   AO22CHD U2479 (.O(n1054), 
	.B2(n101), 
	.B1(\ram[29][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n496));
   AO22CHD U2480 (.O(n1055), 
	.B2(n101), 
	.B1(\ram[29][9] ), 
	.A2(n17), 
	.A1(n496));
   AO22CHD U2481 (.O(n1056), 
	.B2(n101), 
	.B1(\ram[29][10] ), 
	.A2(n18), 
	.A1(n496));
   AO22CHD U2482 (.O(n1057), 
	.B2(n101), 
	.B1(\ram[29][11] ), 
	.A2(n19), 
	.A1(n496));
   AO22CHD U2483 (.O(n1058), 
	.B2(n101), 
	.B1(\ram[29][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n496));
   AO22CHD U2484 (.O(n1059), 
	.B2(n101), 
	.B1(\ram[29][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n496));
   AO22CHD U2485 (.O(n1060), 
	.B2(n101), 
	.B1(\ram[29][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n496));
   AO22CHD U2486 (.O(n1061), 
	.B2(n101), 
	.B1(\ram[29][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n496));
   AO22CHD U2487 (.O(n1062), 
	.B2(n103), 
	.B1(\ram[30][0] ), 
	.A2(n6), 
	.A1(n498));
   AO22CHD U2488 (.O(n1063), 
	.B2(n103), 
	.B1(\ram[30][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n498));
   AO22CHD U2489 (.O(n1064), 
	.B2(n103), 
	.B1(\ram[30][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n498));
   AO22CHD U2490 (.O(n1065), 
	.B2(n103), 
	.B1(\ram[30][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n498));
   AO22CHD U2491 (.O(n1066), 
	.B2(n103), 
	.B1(\ram[30][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n498));
   AO22CHD U2492 (.O(n1067), 
	.B2(n103), 
	.B1(\ram[30][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n498));
   AO22CHD U2493 (.O(n1068), 
	.B2(n103), 
	.B1(\ram[30][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n498));
   AO22CHD U2494 (.O(n1069), 
	.B2(n103), 
	.B1(\ram[30][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n498));
   AO22CHD U2495 (.O(n1070), 
	.B2(n103), 
	.B1(\ram[30][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n498));
   AO22CHD U2496 (.O(n1071), 
	.B2(n103), 
	.B1(\ram[30][9] ), 
	.A2(n17), 
	.A1(n498));
   AO22CHD U2497 (.O(n1072), 
	.B2(n103), 
	.B1(\ram[30][10] ), 
	.A2(n18), 
	.A1(n498));
   AO22CHD U2498 (.O(n1073), 
	.B2(n103), 
	.B1(\ram[30][11] ), 
	.A2(n19), 
	.A1(n498));
   AO22CHD U2499 (.O(n1074), 
	.B2(n103), 
	.B1(\ram[30][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n498));
   AO22CHD U2500 (.O(n1075), 
	.B2(n103), 
	.B1(\ram[30][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n498));
   AO22CHD U2501 (.O(n1076), 
	.B2(n103), 
	.B1(\ram[30][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n498));
   AO22CHD U2502 (.O(n1077), 
	.B2(n103), 
	.B1(\ram[30][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n498));
   AO22CHD U2503 (.O(n1078), 
	.B2(n105), 
	.B1(\ram[31][0] ), 
	.A2(n6), 
	.A1(n500));
   AO22CHD U2504 (.O(n1079), 
	.B2(n105), 
	.B1(\ram[31][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n500));
   AO22CHD U2505 (.O(n1080), 
	.B2(n105), 
	.B1(\ram[31][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n500));
   AO22CHD U2506 (.O(n1081), 
	.B2(n105), 
	.B1(\ram[31][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n500));
   AO22CHD U2507 (.O(n1082), 
	.B2(n105), 
	.B1(\ram[31][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n500));
   AO22CHD U2508 (.O(n1083), 
	.B2(n105), 
	.B1(\ram[31][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n500));
   AO22CHD U2509 (.O(n1084), 
	.B2(n105), 
	.B1(\ram[31][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n500));
   AO22CHD U2510 (.O(n1085), 
	.B2(n105), 
	.B1(\ram[31][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n500));
   AO22CHD U2511 (.O(n1086), 
	.B2(n105), 
	.B1(\ram[31][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n500));
   AO22CHD U2512 (.O(n1087), 
	.B2(n105), 
	.B1(\ram[31][9] ), 
	.A2(n17), 
	.A1(n500));
   AO22CHD U2513 (.O(n1088), 
	.B2(n105), 
	.B1(\ram[31][10] ), 
	.A2(n18), 
	.A1(n500));
   AO22CHD U2514 (.O(n1089), 
	.B2(n105), 
	.B1(\ram[31][11] ), 
	.A2(n19), 
	.A1(n500));
   AO22CHD U2515 (.O(n1090), 
	.B2(n105), 
	.B1(\ram[31][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n500));
   AO22CHD U2516 (.O(n1091), 
	.B2(n105), 
	.B1(\ram[31][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n500));
   AO22CHD U2517 (.O(n1092), 
	.B2(n105), 
	.B1(\ram[31][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n500));
   AO22CHD U2518 (.O(n1093), 
	.B2(n105), 
	.B1(\ram[31][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n500));
   AO22CHD U2519 (.O(n1094), 
	.B2(n108), 
	.B1(\ram[32][0] ), 
	.A2(n6), 
	.A1(n502));
   AO22CHD U2520 (.O(n1095), 
	.B2(n108), 
	.B1(\ram[32][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n502));
   AO22CHD U2521 (.O(n1096), 
	.B2(n108), 
	.B1(\ram[32][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n502));
   AO22CHD U2522 (.O(n1097), 
	.B2(n108), 
	.B1(\ram[32][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n502));
   AO22CHD U2523 (.O(n1098), 
	.B2(n108), 
	.B1(\ram[32][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n502));
   AO22CHD U2524 (.O(n1099), 
	.B2(n108), 
	.B1(\ram[32][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n502));
   AO22CHD U2525 (.O(n1100), 
	.B2(n108), 
	.B1(\ram[32][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n502));
   AO22CHD U2526 (.O(n1101), 
	.B2(n108), 
	.B1(\ram[32][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n502));
   AO22CHD U2527 (.O(n1102), 
	.B2(n108), 
	.B1(\ram[32][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n502));
   AO22CHD U2528 (.O(n1103), 
	.B2(n108), 
	.B1(\ram[32][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n502));
   AO22CHD U2529 (.O(n1104), 
	.B2(n108), 
	.B1(\ram[32][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n502));
   AO22CHD U2530 (.O(n1105), 
	.B2(n108), 
	.B1(\ram[32][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n502));
   AO22CHD U2531 (.O(n1106), 
	.B2(n108), 
	.B1(\ram[32][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n502));
   AO22CHD U2532 (.O(n1107), 
	.B2(n108), 
	.B1(\ram[32][13] ), 
	.A2(n21), 
	.A1(n502));
   AO22CHD U2533 (.O(n1108), 
	.B2(n108), 
	.B1(\ram[32][14] ), 
	.A2(n22), 
	.A1(n502));
   AO22CHD U2534 (.O(n1109), 
	.B2(n108), 
	.B1(\ram[32][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n502));
   AO22CHD U2535 (.O(n1110), 
	.B2(n111), 
	.B1(\ram[33][0] ), 
	.A2(n6), 
	.A1(n504));
   AO22CHD U2536 (.O(n1111), 
	.B2(n111), 
	.B1(\ram[33][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n504));
   AO22CHD U2537 (.O(n1112), 
	.B2(n111), 
	.B1(\ram[33][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n504));
   AO22CHD U2538 (.O(n1113), 
	.B2(n111), 
	.B1(\ram[33][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n504));
   AO22CHD U2539 (.O(n1114), 
	.B2(n111), 
	.B1(\ram[33][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n504));
   AO22CHD U2540 (.O(n1115), 
	.B2(n111), 
	.B1(\ram[33][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n504));
   AO22CHD U2541 (.O(n1116), 
	.B2(n111), 
	.B1(\ram[33][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n504));
   AO22CHD U2542 (.O(n1117), 
	.B2(n111), 
	.B1(\ram[33][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n504));
   AO22CHD U2543 (.O(n1118), 
	.B2(n111), 
	.B1(\ram[33][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n504));
   AO22CHD U2544 (.O(n1119), 
	.B2(n111), 
	.B1(\ram[33][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n504));
   AO22CHD U2545 (.O(n1120), 
	.B2(n111), 
	.B1(\ram[33][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n504));
   AO22CHD U2546 (.O(n1121), 
	.B2(n111), 
	.B1(\ram[33][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n504));
   AO22CHD U2547 (.O(n1122), 
	.B2(n111), 
	.B1(\ram[33][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n504));
   AO22CHD U2548 (.O(n1123), 
	.B2(n111), 
	.B1(\ram[33][13] ), 
	.A2(n21), 
	.A1(n504));
   AO22CHD U2549 (.O(n1124), 
	.B2(n111), 
	.B1(\ram[33][14] ), 
	.A2(n22), 
	.A1(n504));
   AO22CHD U2550 (.O(n1125), 
	.B2(n111), 
	.B1(\ram[33][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n504));
   AO22CHD U2551 (.O(n1126), 
	.B2(n113), 
	.B1(\ram[34][0] ), 
	.A2(n6), 
	.A1(n506));
   AO22CHD U2552 (.O(n1127), 
	.B2(n113), 
	.B1(\ram[34][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n506));
   AO22CHD U2553 (.O(n1128), 
	.B2(n113), 
	.B1(\ram[34][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n506));
   AO22CHD U2554 (.O(n1129), 
	.B2(n113), 
	.B1(\ram[34][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n506));
   AO22CHD U2555 (.O(n1130), 
	.B2(n113), 
	.B1(\ram[34][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n506));
   AO22CHD U2556 (.O(n1131), 
	.B2(n113), 
	.B1(\ram[34][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n506));
   AO22CHD U2557 (.O(n1132), 
	.B2(n113), 
	.B1(\ram[34][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n506));
   AO22CHD U2558 (.O(n1133), 
	.B2(n113), 
	.B1(\ram[34][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n506));
   AO22CHD U2559 (.O(n1134), 
	.B2(n113), 
	.B1(\ram[34][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n506));
   AO22CHD U2560 (.O(n1135), 
	.B2(n113), 
	.B1(\ram[34][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n506));
   AO22CHD U2561 (.O(n1136), 
	.B2(n113), 
	.B1(\ram[34][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n506));
   AO22CHD U2562 (.O(n1137), 
	.B2(n113), 
	.B1(\ram[34][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n506));
   AO22CHD U2563 (.O(n1138), 
	.B2(n113), 
	.B1(\ram[34][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n506));
   AO22CHD U2564 (.O(n1139), 
	.B2(n113), 
	.B1(\ram[34][13] ), 
	.A2(n21), 
	.A1(n506));
   AO22CHD U2565 (.O(n1140), 
	.B2(n113), 
	.B1(\ram[34][14] ), 
	.A2(n22), 
	.A1(n506));
   AO22CHD U2566 (.O(n1141), 
	.B2(n113), 
	.B1(\ram[34][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n506));
   AO22CHD U2567 (.O(n1142), 
	.B2(n115), 
	.B1(\ram[35][0] ), 
	.A2(n6), 
	.A1(n508));
   AO22CHD U2568 (.O(n1143), 
	.B2(n115), 
	.B1(\ram[35][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n508));
   AO22CHD U2569 (.O(n1144), 
	.B2(n115), 
	.B1(\ram[35][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n508));
   AO22CHD U2570 (.O(n1145), 
	.B2(n115), 
	.B1(\ram[35][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n508));
   AO22CHD U2571 (.O(n1146), 
	.B2(n115), 
	.B1(\ram[35][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n508));
   AO22CHD U2572 (.O(n1147), 
	.B2(n115), 
	.B1(\ram[35][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n508));
   AO22CHD U2573 (.O(n1148), 
	.B2(n115), 
	.B1(\ram[35][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n508));
   AO22CHD U2574 (.O(n1149), 
	.B2(n115), 
	.B1(\ram[35][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n508));
   AO22CHD U2575 (.O(n1150), 
	.B2(n115), 
	.B1(\ram[35][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n508));
   AO22CHD U2576 (.O(n1151), 
	.B2(n115), 
	.B1(\ram[35][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n508));
   AO22CHD U2577 (.O(n1152), 
	.B2(n115), 
	.B1(\ram[35][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n508));
   AO22CHD U2578 (.O(n1153), 
	.B2(n115), 
	.B1(\ram[35][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n508));
   AO22CHD U2579 (.O(n1154), 
	.B2(n115), 
	.B1(\ram[35][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n508));
   AO22CHD U2580 (.O(n1155), 
	.B2(n115), 
	.B1(\ram[35][13] ), 
	.A2(n21), 
	.A1(n508));
   AO22CHD U2581 (.O(n1156), 
	.B2(n115), 
	.B1(\ram[35][14] ), 
	.A2(n22), 
	.A1(n508));
   AO22CHD U2582 (.O(n1157), 
	.B2(n115), 
	.B1(\ram[35][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n508));
   AO22CHD U2583 (.O(n1158), 
	.B2(n117), 
	.B1(\ram[36][0] ), 
	.A2(n6), 
	.A1(n510));
   AO22CHD U2584 (.O(n1159), 
	.B2(n117), 
	.B1(\ram[36][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n510));
   AO22CHD U2585 (.O(n1160), 
	.B2(n117), 
	.B1(\ram[36][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n510));
   AO22CHD U2586 (.O(n1161), 
	.B2(n117), 
	.B1(\ram[36][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n510));
   AO22CHD U2587 (.O(n1162), 
	.B2(n117), 
	.B1(\ram[36][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n510));
   AO22CHD U2588 (.O(n1163), 
	.B2(n117), 
	.B1(\ram[36][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n510));
   AO22CHD U2589 (.O(n1164), 
	.B2(n117), 
	.B1(\ram[36][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n510));
   AO22CHD U2590 (.O(n1165), 
	.B2(n117), 
	.B1(\ram[36][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n510));
   AO22CHD U2591 (.O(n1166), 
	.B2(n117), 
	.B1(\ram[36][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n510));
   AO22CHD U2592 (.O(n1167), 
	.B2(n117), 
	.B1(\ram[36][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n510));
   AO22CHD U2593 (.O(n1168), 
	.B2(n117), 
	.B1(\ram[36][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n510));
   AO22CHD U2594 (.O(n1169), 
	.B2(n117), 
	.B1(\ram[36][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n510));
   AO22CHD U2595 (.O(n1170), 
	.B2(n117), 
	.B1(\ram[36][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n510));
   AO22CHD U2596 (.O(n1171), 
	.B2(n117), 
	.B1(\ram[36][13] ), 
	.A2(n21), 
	.A1(n510));
   AO22CHD U2597 (.O(n1172), 
	.B2(n117), 
	.B1(\ram[36][14] ), 
	.A2(n22), 
	.A1(n510));
   AO22CHD U2598 (.O(n1173), 
	.B2(n117), 
	.B1(\ram[36][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n510));
   AO22CHD U2599 (.O(n1174), 
	.B2(n119), 
	.B1(\ram[37][0] ), 
	.A2(n6), 
	.A1(n511));
   AO22CHD U2600 (.O(n1175), 
	.B2(n119), 
	.B1(\ram[37][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n511));
   AO22CHD U2601 (.O(n1176), 
	.B2(n119), 
	.B1(\ram[37][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n511));
   AO22CHD U2602 (.O(n1177), 
	.B2(n119), 
	.B1(\ram[37][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n511));
   AO22CHD U2603 (.O(n1178), 
	.B2(n119), 
	.B1(\ram[37][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n511));
   AO22CHD U2604 (.O(n1179), 
	.B2(n119), 
	.B1(\ram[37][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n511));
   AO22CHD U2605 (.O(n1180), 
	.B2(n119), 
	.B1(\ram[37][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n511));
   AO22CHD U2606 (.O(n1181), 
	.B2(n119), 
	.B1(\ram[37][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n511));
   AO22CHD U2607 (.O(n1182), 
	.B2(n119), 
	.B1(\ram[37][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n511));
   AO22CHD U2608 (.O(n1183), 
	.B2(n119), 
	.B1(\ram[37][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n511));
   AO22CHD U2609 (.O(n1184), 
	.B2(n119), 
	.B1(\ram[37][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n511));
   AO22CHD U2610 (.O(n1185), 
	.B2(n119), 
	.B1(\ram[37][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n511));
   AO22CHD U2611 (.O(n1186), 
	.B2(n119), 
	.B1(\ram[37][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n511));
   AO22CHD U2612 (.O(n1187), 
	.B2(n119), 
	.B1(\ram[37][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n511));
   AO22CHD U2613 (.O(n1188), 
	.B2(n119), 
	.B1(\ram[37][14] ), 
	.A2(n22), 
	.A1(n511));
   AO22CHD U2614 (.O(n1189), 
	.B2(n119), 
	.B1(\ram[37][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n511));
   AO22CHD U2615 (.O(n1190), 
	.B2(n121), 
	.B1(\ram[38][0] ), 
	.A2(n6), 
	.A1(n513));
   AO22CHD U2616 (.O(n1191), 
	.B2(n121), 
	.B1(\ram[38][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n513));
   AO22CHD U2617 (.O(n1192), 
	.B2(n121), 
	.B1(\ram[38][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n513));
   AO22CHD U2618 (.O(n1193), 
	.B2(n121), 
	.B1(\ram[38][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n513));
   AO22CHD U2619 (.O(n1194), 
	.B2(n121), 
	.B1(\ram[38][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n513));
   AO22CHD U2620 (.O(n1195), 
	.B2(n121), 
	.B1(\ram[38][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n513));
   AO22CHD U2621 (.O(n1196), 
	.B2(n121), 
	.B1(\ram[38][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n513));
   AO22CHD U2622 (.O(n1197), 
	.B2(n121), 
	.B1(\ram[38][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n513));
   AO22CHD U2623 (.O(n1198), 
	.B2(n121), 
	.B1(\ram[38][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n513));
   AO22CHD U2624 (.O(n1199), 
	.B2(n121), 
	.B1(\ram[38][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n513));
   AO22CHD U2625 (.O(n1200), 
	.B2(n121), 
	.B1(\ram[38][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n513));
   AO22CHD U2626 (.O(n1201), 
	.B2(n121), 
	.B1(\ram[38][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n513));
   AO22CHD U2627 (.O(n1202), 
	.B2(n121), 
	.B1(\ram[38][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n513));
   AO22CHD U2628 (.O(n1203), 
	.B2(n121), 
	.B1(\ram[38][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n513));
   AO22CHD U2629 (.O(n1204), 
	.B2(n121), 
	.B1(\ram[38][14] ), 
	.A2(n22), 
	.A1(n513));
   AO22CHD U2630 (.O(n1205), 
	.B2(n121), 
	.B1(\ram[38][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n513));
   AO22CHD U2631 (.O(n1206), 
	.B2(n123), 
	.B1(\ram[39][0] ), 
	.A2(n6), 
	.A1(n515));
   AO22CHD U2632 (.O(n1207), 
	.B2(n123), 
	.B1(\ram[39][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n515));
   AO22CHD U2633 (.O(n1208), 
	.B2(n123), 
	.B1(\ram[39][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n515));
   AO22CHD U2634 (.O(n1209), 
	.B2(n123), 
	.B1(\ram[39][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n515));
   AO22CHD U2635 (.O(n1210), 
	.B2(n123), 
	.B1(\ram[39][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n515));
   AO22CHD U2636 (.O(n1211), 
	.B2(n123), 
	.B1(\ram[39][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n515));
   AO22CHD U2637 (.O(n1212), 
	.B2(n123), 
	.B1(\ram[39][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n515));
   AO22CHD U2638 (.O(n1213), 
	.B2(n123), 
	.B1(\ram[39][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n515));
   AO22CHD U2639 (.O(n1214), 
	.B2(n123), 
	.B1(\ram[39][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n515));
   AO22CHD U2640 (.O(n1215), 
	.B2(n123), 
	.B1(\ram[39][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n515));
   AO22CHD U2641 (.O(n1216), 
	.B2(n123), 
	.B1(\ram[39][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n515));
   AO22CHD U2642 (.O(n1217), 
	.B2(n123), 
	.B1(\ram[39][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n515));
   AO22CHD U2643 (.O(n1218), 
	.B2(n123), 
	.B1(\ram[39][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n515));
   AO22CHD U2644 (.O(n1219), 
	.B2(n123), 
	.B1(\ram[39][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n515));
   AO22CHD U2645 (.O(n1220), 
	.B2(n123), 
	.B1(\ram[39][14] ), 
	.A2(n22), 
	.A1(n515));
   AO22CHD U2646 (.O(n1221), 
	.B2(n123), 
	.B1(\ram[39][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n515));
   AO22CHD U2647 (.O(n1222), 
	.B2(n125), 
	.B1(\ram[40][0] ), 
	.A2(n6), 
	.A1(n517));
   AO22CHD U2648 (.O(n1223), 
	.B2(n125), 
	.B1(\ram[40][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n517));
   AO22CHD U2649 (.O(n1224), 
	.B2(n125), 
	.B1(\ram[40][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n517));
   AO22CHD U2650 (.O(n1225), 
	.B2(n125), 
	.B1(\ram[40][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n517));
   AO22CHD U2651 (.O(n1226), 
	.B2(n125), 
	.B1(\ram[40][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n517));
   AO22CHD U2652 (.O(n1227), 
	.B2(n125), 
	.B1(\ram[40][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n517));
   AO22CHD U2653 (.O(n1228), 
	.B2(n125), 
	.B1(\ram[40][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n517));
   AO22CHD U2654 (.O(n1229), 
	.B2(n125), 
	.B1(\ram[40][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n517));
   AO22CHD U2655 (.O(n1230), 
	.B2(n125), 
	.B1(\ram[40][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n517));
   AO22CHD U2656 (.O(n1231), 
	.B2(n125), 
	.B1(\ram[40][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n517));
   AO22CHD U2657 (.O(n1232), 
	.B2(n125), 
	.B1(\ram[40][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n517));
   AO22CHD U2658 (.O(n1233), 
	.B2(n125), 
	.B1(\ram[40][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n517));
   AO22CHD U2659 (.O(n1234), 
	.B2(n125), 
	.B1(\ram[40][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n517));
   AO22CHD U2660 (.O(n1235), 
	.B2(n125), 
	.B1(\ram[40][13] ), 
	.A2(n21), 
	.A1(n517));
   AO22CHD U2661 (.O(n1236), 
	.B2(n125), 
	.B1(\ram[40][14] ), 
	.A2(n22), 
	.A1(n517));
   AO22CHD U2662 (.O(n1237), 
	.B2(n125), 
	.B1(\ram[40][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n517));
   AO22CHD U2663 (.O(n1238), 
	.B2(n127), 
	.B1(\ram[41][0] ), 
	.A2(n6), 
	.A1(n519));
   AO22CHD U2664 (.O(n1239), 
	.B2(n127), 
	.B1(\ram[41][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n519));
   AO22CHD U2665 (.O(n1240), 
	.B2(n127), 
	.B1(\ram[41][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n519));
   AO22CHD U2666 (.O(n1241), 
	.B2(n127), 
	.B1(\ram[41][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n519));
   AO22CHD U2667 (.O(n1242), 
	.B2(n127), 
	.B1(\ram[41][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n519));
   AO22CHD U2668 (.O(n1243), 
	.B2(n127), 
	.B1(\ram[41][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n519));
   AO22CHD U2669 (.O(n1244), 
	.B2(n127), 
	.B1(\ram[41][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n519));
   AO22CHD U2670 (.O(n1245), 
	.B2(n127), 
	.B1(\ram[41][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n519));
   AO22CHD U2671 (.O(n1246), 
	.B2(n127), 
	.B1(\ram[41][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n519));
   AO22CHD U2672 (.O(n1247), 
	.B2(n127), 
	.B1(\ram[41][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n519));
   AO22CHD U2673 (.O(n1248), 
	.B2(n127), 
	.B1(\ram[41][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n519));
   AO22CHD U2674 (.O(n1249), 
	.B2(n127), 
	.B1(\ram[41][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n519));
   AO22CHD U2675 (.O(n1250), 
	.B2(n127), 
	.B1(\ram[41][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n519));
   AO22CHD U2676 (.O(n1251), 
	.B2(n127), 
	.B1(\ram[41][13] ), 
	.A2(n21), 
	.A1(n519));
   AO22CHD U2677 (.O(n1252), 
	.B2(n127), 
	.B1(\ram[41][14] ), 
	.A2(n22), 
	.A1(n519));
   AO22CHD U2678 (.O(n1253), 
	.B2(n127), 
	.B1(\ram[41][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n519));
   AO22CHD U2679 (.O(n1254), 
	.B2(n129), 
	.B1(\ram[42][0] ), 
	.A2(n6), 
	.A1(n521));
   AO22CHD U2680 (.O(n1255), 
	.B2(n129), 
	.B1(\ram[42][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n521));
   AO22CHD U2681 (.O(n1256), 
	.B2(n129), 
	.B1(\ram[42][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n521));
   AO22CHD U2682 (.O(n1257), 
	.B2(n129), 
	.B1(\ram[42][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n521));
   AO22CHD U2683 (.O(n1258), 
	.B2(n129), 
	.B1(\ram[42][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n521));
   AO22CHD U2684 (.O(n1259), 
	.B2(n129), 
	.B1(\ram[42][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n521));
   AO22CHD U2685 (.O(n1260), 
	.B2(n129), 
	.B1(\ram[42][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n521));
   AO22CHD U2686 (.O(n1261), 
	.B2(n129), 
	.B1(\ram[42][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n521));
   AO22CHD U2687 (.O(n1262), 
	.B2(n129), 
	.B1(\ram[42][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n521));
   AO22CHD U2688 (.O(n1263), 
	.B2(n129), 
	.B1(\ram[42][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n521));
   AO22CHD U2689 (.O(n1264), 
	.B2(n129), 
	.B1(\ram[42][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n521));
   AO22CHD U2690 (.O(n1265), 
	.B2(n129), 
	.B1(\ram[42][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n521));
   AO22CHD U2691 (.O(n1266), 
	.B2(n129), 
	.B1(\ram[42][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n521));
   AO22CHD U2692 (.O(n1267), 
	.B2(n129), 
	.B1(\ram[42][13] ), 
	.A2(n21), 
	.A1(n521));
   AO22CHD U2693 (.O(n1268), 
	.B2(n129), 
	.B1(\ram[42][14] ), 
	.A2(n22), 
	.A1(n521));
   AO22CHD U2694 (.O(n1269), 
	.B2(n129), 
	.B1(\ram[42][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n521));
   AO22CHD U2695 (.O(n1270), 
	.B2(n131), 
	.B1(\ram[43][0] ), 
	.A2(n6), 
	.A1(n523));
   AO22CHD U2696 (.O(n1271), 
	.B2(n131), 
	.B1(\ram[43][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n523));
   AO22CHD U2697 (.O(n1272), 
	.B2(n131), 
	.B1(\ram[43][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n523));
   AO22CHD U2698 (.O(n1273), 
	.B2(n131), 
	.B1(\ram[43][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n523));
   AO22CHD U2699 (.O(n1274), 
	.B2(n131), 
	.B1(\ram[43][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n523));
   AO22CHD U2700 (.O(n1275), 
	.B2(n131), 
	.B1(\ram[43][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n523));
   AO22CHD U2701 (.O(n1276), 
	.B2(n131), 
	.B1(\ram[43][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n523));
   AO22CHD U2702 (.O(n1277), 
	.B2(n131), 
	.B1(\ram[43][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n523));
   AO22CHD U2703 (.O(n1278), 
	.B2(n131), 
	.B1(\ram[43][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n523));
   AO22CHD U2704 (.O(n1279), 
	.B2(n131), 
	.B1(\ram[43][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n523));
   AO22CHD U2705 (.O(n1280), 
	.B2(n131), 
	.B1(\ram[43][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n523));
   AO22CHD U2706 (.O(n1281), 
	.B2(n131), 
	.B1(\ram[43][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n523));
   AO22CHD U2707 (.O(n1282), 
	.B2(n131), 
	.B1(\ram[43][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n523));
   AO22CHD U2708 (.O(n1283), 
	.B2(n131), 
	.B1(\ram[43][13] ), 
	.A2(n21), 
	.A1(n523));
   AO22CHD U2709 (.O(n1284), 
	.B2(n131), 
	.B1(\ram[43][14] ), 
	.A2(n22), 
	.A1(n523));
   AO22CHD U2710 (.O(n1285), 
	.B2(n131), 
	.B1(\ram[43][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n523));
   AO22CHD U2711 (.O(n1286), 
	.B2(n133), 
	.B1(\ram[44][0] ), 
	.A2(n6), 
	.A1(n525));
   AO22CHD U2712 (.O(n1287), 
	.B2(n133), 
	.B1(\ram[44][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n525));
   AO22CHD U2713 (.O(n1288), 
	.B2(n133), 
	.B1(\ram[44][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n525));
   AO22CHD U2714 (.O(n1289), 
	.B2(n133), 
	.B1(\ram[44][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n525));
   AO22CHD U2715 (.O(n1290), 
	.B2(n133), 
	.B1(\ram[44][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n525));
   AO22CHD U2716 (.O(n1291), 
	.B2(n133), 
	.B1(\ram[44][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n525));
   AO22CHD U2717 (.O(n1292), 
	.B2(n133), 
	.B1(\ram[44][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n525));
   AO22CHD U2718 (.O(n1293), 
	.B2(n133), 
	.B1(\ram[44][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n525));
   AO22CHD U2719 (.O(n1294), 
	.B2(n133), 
	.B1(\ram[44][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n525));
   AO22CHD U2720 (.O(n1295), 
	.B2(n133), 
	.B1(\ram[44][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n525));
   AO22CHD U2721 (.O(n1296), 
	.B2(n133), 
	.B1(\ram[44][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n525));
   AO22CHD U2722 (.O(n1297), 
	.B2(n133), 
	.B1(\ram[44][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n525));
   AO22CHD U2723 (.O(n1298), 
	.B2(n133), 
	.B1(\ram[44][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n525));
   AO22CHD U2724 (.O(n1299), 
	.B2(n133), 
	.B1(\ram[44][13] ), 
	.A2(n21), 
	.A1(n525));
   AO22CHD U2725 (.O(n1300), 
	.B2(n133), 
	.B1(\ram[44][14] ), 
	.A2(n22), 
	.A1(n525));
   AO22CHD U2726 (.O(n1301), 
	.B2(n133), 
	.B1(\ram[44][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n525));
   AO22CHD U2727 (.O(n1302), 
	.B2(n135), 
	.B1(\ram[45][0] ), 
	.A2(n6), 
	.A1(n527));
   AO22CHD U2728 (.O(n1303), 
	.B2(n135), 
	.B1(\ram[45][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n527));
   AO22CHD U2729 (.O(n1304), 
	.B2(n135), 
	.B1(\ram[45][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n527));
   AO22CHD U2730 (.O(n1305), 
	.B2(n135), 
	.B1(\ram[45][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n527));
   AO22CHD U2731 (.O(n1306), 
	.B2(n135), 
	.B1(\ram[45][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n527));
   AO22CHD U2732 (.O(n1307), 
	.B2(n135), 
	.B1(\ram[45][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n527));
   AO22CHD U2733 (.O(n1308), 
	.B2(n135), 
	.B1(\ram[45][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n527));
   AO22CHD U2734 (.O(n1309), 
	.B2(n135), 
	.B1(\ram[45][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n527));
   AO22CHD U2735 (.O(n1310), 
	.B2(n135), 
	.B1(\ram[45][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n527));
   AO22CHD U2736 (.O(n1311), 
	.B2(n135), 
	.B1(\ram[45][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n527));
   AO22CHD U2737 (.O(n1312), 
	.B2(n135), 
	.B1(\ram[45][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n527));
   AO22CHD U2738 (.O(n1313), 
	.B2(n135), 
	.B1(\ram[45][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n527));
   AO22CHD U2739 (.O(n1314), 
	.B2(n135), 
	.B1(\ram[45][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n527));
   AO22CHD U2740 (.O(n1315), 
	.B2(n135), 
	.B1(\ram[45][13] ), 
	.A2(n21), 
	.A1(n527));
   AO22CHD U2741 (.O(n1316), 
	.B2(n135), 
	.B1(\ram[45][14] ), 
	.A2(n22), 
	.A1(n527));
   AO22CHD U2742 (.O(n1317), 
	.B2(n135), 
	.B1(\ram[45][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n527));
   AO22CHD U2743 (.O(n1318), 
	.B2(n137), 
	.B1(\ram[46][0] ), 
	.A2(n6), 
	.A1(n529));
   AO22CHD U2744 (.O(n1319), 
	.B2(n137), 
	.B1(\ram[46][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n529));
   AO22CHD U2745 (.O(n1320), 
	.B2(n137), 
	.B1(\ram[46][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n529));
   AO22CHD U2746 (.O(n1321), 
	.B2(n137), 
	.B1(\ram[46][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n529));
   AO22CHD U2747 (.O(n1322), 
	.B2(n137), 
	.B1(\ram[46][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n529));
   AO22CHD U2748 (.O(n1323), 
	.B2(n137), 
	.B1(\ram[46][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n529));
   AO22CHD U2749 (.O(n1324), 
	.B2(n137), 
	.B1(\ram[46][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n529));
   AO22CHD U2750 (.O(n1325), 
	.B2(n137), 
	.B1(\ram[46][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n529));
   AO22CHD U2751 (.O(n1326), 
	.B2(n137), 
	.B1(\ram[46][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n529));
   AO22CHD U2752 (.O(n1327), 
	.B2(n137), 
	.B1(\ram[46][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n529));
   AO22CHD U2753 (.O(n1328), 
	.B2(n137), 
	.B1(\ram[46][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n529));
   AO22CHD U2754 (.O(n1329), 
	.B2(n137), 
	.B1(\ram[46][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n529));
   AO22CHD U2755 (.O(n1330), 
	.B2(n137), 
	.B1(\ram[46][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n529));
   AO22CHD U2756 (.O(n1331), 
	.B2(n137), 
	.B1(\ram[46][13] ), 
	.A2(n21), 
	.A1(n529));
   AO22CHD U2757 (.O(n1332), 
	.B2(n137), 
	.B1(\ram[46][14] ), 
	.A2(n22), 
	.A1(n529));
   AO22CHD U2758 (.O(n1333), 
	.B2(n137), 
	.B1(\ram[46][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n529));
   AO22CHD U2759 (.O(n1334), 
	.B2(n139), 
	.B1(\ram[47][0] ), 
	.A2(n6), 
	.A1(n531));
   AO22CHD U2760 (.O(n1335), 
	.B2(n139), 
	.B1(\ram[47][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n531));
   AO22CHD U2761 (.O(n1336), 
	.B2(n139), 
	.B1(\ram[47][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n531));
   AO22CHD U2762 (.O(n1337), 
	.B2(n139), 
	.B1(\ram[47][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n531));
   AO22CHD U2763 (.O(n1338), 
	.B2(n139), 
	.B1(\ram[47][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n531));
   AO22CHD U2764 (.O(n1339), 
	.B2(n139), 
	.B1(\ram[47][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n531));
   AO22CHD U2765 (.O(n1340), 
	.B2(n139), 
	.B1(\ram[47][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n531));
   AO22CHD U2766 (.O(n1341), 
	.B2(n139), 
	.B1(\ram[47][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n531));
   AO22CHD U2767 (.O(n1342), 
	.B2(n139), 
	.B1(\ram[47][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n531));
   AO22CHD U2768 (.O(n1343), 
	.B2(n139), 
	.B1(\ram[47][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n531));
   AO22CHD U2769 (.O(n1344), 
	.B2(n139), 
	.B1(\ram[47][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n531));
   AO22CHD U2770 (.O(n1345), 
	.B2(n139), 
	.B1(\ram[47][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n531));
   AO22CHD U2771 (.O(n1346), 
	.B2(n139), 
	.B1(\ram[47][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n531));
   AO22CHD U2772 (.O(n1347), 
	.B2(n139), 
	.B1(\ram[47][13] ), 
	.A2(n21), 
	.A1(n531));
   AO22CHD U2773 (.O(n1348), 
	.B2(n139), 
	.B1(\ram[47][14] ), 
	.A2(n22), 
	.A1(n531));
   AO22CHD U2774 (.O(n1349), 
	.B2(n139), 
	.B1(\ram[47][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n531));
   AO22CHD U2775 (.O(n1350), 
	.B2(n142), 
	.B1(\ram[48][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n533));
   AO22CHD U2776 (.O(n1351), 
	.B2(n142), 
	.B1(\ram[48][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n533));
   AO22CHD U2777 (.O(n1352), 
	.B2(n142), 
	.B1(\ram[48][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n533));
   AO22CHD U2778 (.O(n1353), 
	.B2(n142), 
	.B1(\ram[48][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n533));
   AO22CHD U2779 (.O(n1354), 
	.B2(n142), 
	.B1(\ram[48][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n533));
   AO22CHD U2780 (.O(n1355), 
	.B2(n142), 
	.B1(\ram[48][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n533));
   AO22CHD U2781 (.O(n1356), 
	.B2(n142), 
	.B1(\ram[48][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n533));
   AO22CHD U2782 (.O(n1357), 
	.B2(n142), 
	.B1(\ram[48][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n533));
   AO22CHD U2783 (.O(n1358), 
	.B2(n142), 
	.B1(\ram[48][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n533));
   AO22CHD U2784 (.O(n1359), 
	.B2(n142), 
	.B1(\ram[48][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n533));
   AO22CHD U2785 (.O(n1360), 
	.B2(n142), 
	.B1(\ram[48][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n533));
   AO22CHD U2786 (.O(n1361), 
	.B2(n142), 
	.B1(\ram[48][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n533));
   AO22CHD U2787 (.O(n1362), 
	.B2(n142), 
	.B1(\ram[48][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n533));
   AO22CHD U2788 (.O(n1363), 
	.B2(n142), 
	.B1(\ram[48][13] ), 
	.A2(n21), 
	.A1(n533));
   AO22CHD U2789 (.O(n1364), 
	.B2(n142), 
	.B1(\ram[48][14] ), 
	.A2(n22), 
	.A1(n533));
   AO22CHD U2790 (.O(n1365), 
	.B2(n142), 
	.B1(\ram[48][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n533));
   AO22CHD U2791 (.O(n1366), 
	.B2(n145), 
	.B1(\ram[49][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n535));
   AO22CHD U2792 (.O(n1367), 
	.B2(n145), 
	.B1(\ram[49][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n535));
   AO22CHD U2793 (.O(n1368), 
	.B2(n145), 
	.B1(\ram[49][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n535));
   AO22CHD U2794 (.O(n1369), 
	.B2(n145), 
	.B1(\ram[49][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n535));
   AO22CHD U2795 (.O(n1370), 
	.B2(n145), 
	.B1(\ram[49][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n535));
   AO22CHD U2796 (.O(n1371), 
	.B2(n145), 
	.B1(\ram[49][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n535));
   AO22CHD U2797 (.O(n1372), 
	.B2(n145), 
	.B1(\ram[49][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n535));
   AO22CHD U2798 (.O(n1373), 
	.B2(n145), 
	.B1(\ram[49][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n535));
   AO22CHD U2799 (.O(n1374), 
	.B2(n145), 
	.B1(\ram[49][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n535));
   AO22CHD U2800 (.O(n1375), 
	.B2(n145), 
	.B1(\ram[49][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n535));
   AO22CHD U2801 (.O(n1376), 
	.B2(n145), 
	.B1(\ram[49][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n535));
   AO22CHD U2802 (.O(n1377), 
	.B2(n145), 
	.B1(\ram[49][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n535));
   AO22CHD U2803 (.O(n1378), 
	.B2(n145), 
	.B1(\ram[49][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n535));
   AO22CHD U2804 (.O(n1379), 
	.B2(n145), 
	.B1(\ram[49][13] ), 
	.A2(n21), 
	.A1(n535));
   AO22CHD U2805 (.O(n1380), 
	.B2(n145), 
	.B1(\ram[49][14] ), 
	.A2(n22), 
	.A1(n535));
   AO22CHD U2806 (.O(n1381), 
	.B2(n145), 
	.B1(\ram[49][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n535));
   AO22CHD U2807 (.O(n1382), 
	.B2(n147), 
	.B1(\ram[50][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n537));
   AO22CHD U2808 (.O(n1383), 
	.B2(n147), 
	.B1(\ram[50][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n537));
   AO22CHD U2809 (.O(n1384), 
	.B2(n147), 
	.B1(\ram[50][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n537));
   AO22CHD U2810 (.O(n1385), 
	.B2(n147), 
	.B1(\ram[50][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n537));
   AO22CHD U2811 (.O(n1386), 
	.B2(n147), 
	.B1(\ram[50][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n537));
   AO22CHD U2812 (.O(n1387), 
	.B2(n147), 
	.B1(\ram[50][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n537));
   AO22CHD U2813 (.O(n1388), 
	.B2(n147), 
	.B1(\ram[50][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n537));
   AO22CHD U2814 (.O(n1389), 
	.B2(n147), 
	.B1(\ram[50][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n537));
   AO22CHD U2815 (.O(n1390), 
	.B2(n147), 
	.B1(\ram[50][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n537));
   AO22CHD U2816 (.O(n1391), 
	.B2(n147), 
	.B1(\ram[50][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n537));
   AO22CHD U2817 (.O(n1392), 
	.B2(n147), 
	.B1(\ram[50][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n537));
   AO22CHD U2818 (.O(n1393), 
	.B2(n147), 
	.B1(\ram[50][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n537));
   AO22CHD U2819 (.O(n1394), 
	.B2(n147), 
	.B1(\ram[50][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n537));
   AO22CHD U2820 (.O(n1395), 
	.B2(n147), 
	.B1(\ram[50][13] ), 
	.A2(n21), 
	.A1(n537));
   AO22CHD U2821 (.O(n1396), 
	.B2(n147), 
	.B1(\ram[50][14] ), 
	.A2(n22), 
	.A1(n537));
   AO22CHD U2822 (.O(n1397), 
	.B2(n147), 
	.B1(\ram[50][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n537));
   AO22CHD U2823 (.O(n1398), 
	.B2(n149), 
	.B1(\ram[51][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n539));
   AO22CHD U2824 (.O(n1399), 
	.B2(n149), 
	.B1(\ram[51][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n539));
   AO22CHD U2825 (.O(n1400), 
	.B2(n149), 
	.B1(\ram[51][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n539));
   AO22CHD U2826 (.O(n1401), 
	.B2(n149), 
	.B1(\ram[51][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n539));
   AO22CHD U2827 (.O(n1402), 
	.B2(n149), 
	.B1(\ram[51][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n539));
   AO22CHD U2828 (.O(n1403), 
	.B2(n149), 
	.B1(\ram[51][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n539));
   AO22CHD U2829 (.O(n1404), 
	.B2(n149), 
	.B1(\ram[51][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n539));
   AO22CHD U2830 (.O(n1405), 
	.B2(n149), 
	.B1(\ram[51][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n539));
   AO22CHD U2831 (.O(n1406), 
	.B2(n149), 
	.B1(\ram[51][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n539));
   AO22CHD U2832 (.O(n1407), 
	.B2(n149), 
	.B1(\ram[51][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n539));
   AO22CHD U2833 (.O(n1408), 
	.B2(n149), 
	.B1(\ram[51][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n539));
   AO22CHD U2834 (.O(n1409), 
	.B2(n149), 
	.B1(\ram[51][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n539));
   AO22CHD U2835 (.O(n1410), 
	.B2(n149), 
	.B1(\ram[51][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n539));
   AO22CHD U2836 (.O(n1411), 
	.B2(n149), 
	.B1(\ram[51][13] ), 
	.A2(n21), 
	.A1(n539));
   AO22CHD U2837 (.O(n1412), 
	.B2(n149), 
	.B1(\ram[51][14] ), 
	.A2(n22), 
	.A1(n539));
   AO22CHD U2838 (.O(n1413), 
	.B2(n149), 
	.B1(\ram[51][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n539));
   AO22CHD U2839 (.O(n1414), 
	.B2(n151), 
	.B1(\ram[52][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n541));
   AO22CHD U2840 (.O(n1415), 
	.B2(n151), 
	.B1(\ram[52][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n541));
   AO22CHD U2841 (.O(n1416), 
	.B2(n151), 
	.B1(\ram[52][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n541));
   AO22CHD U2842 (.O(n1417), 
	.B2(n151), 
	.B1(\ram[52][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n541));
   AO22CHD U2843 (.O(n1418), 
	.B2(n151), 
	.B1(\ram[52][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n541));
   AO22CHD U2844 (.O(n1419), 
	.B2(n151), 
	.B1(\ram[52][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n541));
   AO22CHD U2845 (.O(n1420), 
	.B2(n151), 
	.B1(\ram[52][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n541));
   AO22CHD U2846 (.O(n1421), 
	.B2(n151), 
	.B1(\ram[52][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n541));
   AO22CHD U2847 (.O(n1422), 
	.B2(n151), 
	.B1(\ram[52][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n541));
   AO22CHD U2848 (.O(n1423), 
	.B2(n151), 
	.B1(\ram[52][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n541));
   AO22CHD U2849 (.O(n1424), 
	.B2(n151), 
	.B1(\ram[52][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n541));
   AO22CHD U2850 (.O(n1425), 
	.B2(n151), 
	.B1(\ram[52][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n541));
   AO22CHD U2851 (.O(n1426), 
	.B2(n151), 
	.B1(\ram[52][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n541));
   AO22CHD U2852 (.O(n1427), 
	.B2(n151), 
	.B1(\ram[52][13] ), 
	.A2(n21), 
	.A1(n541));
   AO22CHD U2853 (.O(n1428), 
	.B2(n151), 
	.B1(\ram[52][14] ), 
	.A2(n22), 
	.A1(n541));
   AO22CHD U2854 (.O(n1429), 
	.B2(n151), 
	.B1(\ram[52][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n541));
   AO22CHD U2855 (.O(n1430), 
	.B2(n153), 
	.B1(\ram[53][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n543));
   AO22CHD U2856 (.O(n1431), 
	.B2(n153), 
	.B1(\ram[53][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n543));
   AO22CHD U2857 (.O(n1432), 
	.B2(n153), 
	.B1(\ram[53][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n543));
   AO22CHD U2858 (.O(n1433), 
	.B2(n153), 
	.B1(\ram[53][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n543));
   AO22CHD U2859 (.O(n1434), 
	.B2(n153), 
	.B1(\ram[53][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n543));
   AO22CHD U2860 (.O(n1435), 
	.B2(n153), 
	.B1(\ram[53][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n543));
   AO22CHD U2861 (.O(n1436), 
	.B2(n153), 
	.B1(\ram[53][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n543));
   AO22CHD U2862 (.O(n1437), 
	.B2(n153), 
	.B1(\ram[53][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n543));
   AO22CHD U2863 (.O(n1438), 
	.B2(n153), 
	.B1(\ram[53][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n543));
   AO22CHD U2864 (.O(n1439), 
	.B2(n153), 
	.B1(\ram[53][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n543));
   AO22CHD U2865 (.O(n1440), 
	.B2(n153), 
	.B1(\ram[53][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n543));
   AO22CHD U2866 (.O(n1441), 
	.B2(n153), 
	.B1(\ram[53][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n543));
   AO22CHD U2867 (.O(n1442), 
	.B2(n153), 
	.B1(\ram[53][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n543));
   AO22CHD U2868 (.O(n1443), 
	.B2(n153), 
	.B1(\ram[53][13] ), 
	.A2(n21), 
	.A1(n543));
   AO22CHD U2869 (.O(n1444), 
	.B2(n153), 
	.B1(\ram[53][14] ), 
	.A2(n22), 
	.A1(n543));
   AO22CHD U2870 (.O(n1445), 
	.B2(n153), 
	.B1(\ram[53][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n543));
   AO22CHD U2871 (.O(n1446), 
	.B2(n155), 
	.B1(\ram[54][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n546));
   AO22CHD U2872 (.O(n1447), 
	.B2(n155), 
	.B1(\ram[54][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n546));
   AO22CHD U2873 (.O(n1448), 
	.B2(n155), 
	.B1(\ram[54][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n546));
   AO22CHD U2874 (.O(n1449), 
	.B2(n155), 
	.B1(\ram[54][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n546));
   AO22CHD U2875 (.O(n1450), 
	.B2(n155), 
	.B1(\ram[54][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n546));
   AO22CHD U2876 (.O(n1451), 
	.B2(n155), 
	.B1(\ram[54][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n546));
   AO22CHD U2877 (.O(n1452), 
	.B2(n155), 
	.B1(\ram[54][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n546));
   AO22CHD U2878 (.O(n1453), 
	.B2(n155), 
	.B1(\ram[54][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n546));
   AO22CHD U2879 (.O(n1454), 
	.B2(n155), 
	.B1(\ram[54][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n546));
   AO22CHD U2880 (.O(n1455), 
	.B2(n155), 
	.B1(\ram[54][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n546));
   AO22CHD U2881 (.O(n1456), 
	.B2(n155), 
	.B1(\ram[54][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n546));
   AO22CHD U2882 (.O(n1457), 
	.B2(n155), 
	.B1(\ram[54][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n546));
   AO22CHD U2883 (.O(n1458), 
	.B2(n155), 
	.B1(\ram[54][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n546));
   AO22CHD U2884 (.O(n1459), 
	.B2(n155), 
	.B1(\ram[54][13] ), 
	.A2(n21), 
	.A1(n546));
   AO22CHD U2885 (.O(n1460), 
	.B2(n155), 
	.B1(\ram[54][14] ), 
	.A2(n22), 
	.A1(n546));
   AO22CHD U2886 (.O(n1461), 
	.B2(n155), 
	.B1(\ram[54][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n546));
   AO22CHD U2887 (.O(n1462), 
	.B2(n157), 
	.B1(\ram[55][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n549));
   AO22CHD U2888 (.O(n1463), 
	.B2(n157), 
	.B1(\ram[55][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n549));
   AO22CHD U2889 (.O(n1464), 
	.B2(n157), 
	.B1(\ram[55][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n549));
   AO22CHD U2890 (.O(n1465), 
	.B2(n157), 
	.B1(\ram[55][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n549));
   AO22CHD U2891 (.O(n1466), 
	.B2(n157), 
	.B1(\ram[55][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n549));
   AO22CHD U2892 (.O(n1467), 
	.B2(n157), 
	.B1(\ram[55][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n549));
   AO22CHD U2893 (.O(n1468), 
	.B2(n157), 
	.B1(\ram[55][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n549));
   AO22CHD U2894 (.O(n1469), 
	.B2(n157), 
	.B1(\ram[55][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n549));
   AO22CHD U2895 (.O(n1470), 
	.B2(n157), 
	.B1(\ram[55][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n549));
   AO22CHD U2896 (.O(n1471), 
	.B2(n157), 
	.B1(\ram[55][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n549));
   AO22CHD U2897 (.O(n1472), 
	.B2(n157), 
	.B1(\ram[55][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n549));
   AO22CHD U2898 (.O(n1473), 
	.B2(n157), 
	.B1(\ram[55][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n549));
   AO22CHD U2899 (.O(n1474), 
	.B2(n157), 
	.B1(\ram[55][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n549));
   AO22CHD U2900 (.O(n1475), 
	.B2(n157), 
	.B1(\ram[55][13] ), 
	.A2(n21), 
	.A1(n549));
   AO22CHD U2901 (.O(n1476), 
	.B2(n157), 
	.B1(\ram[55][14] ), 
	.A2(n22), 
	.A1(n549));
   AO22CHD U2902 (.O(n1477), 
	.B2(n157), 
	.B1(\ram[55][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n549));
   AO22CHD U2903 (.O(n1478), 
	.B2(n159), 
	.B1(\ram[56][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n552));
   AO22CHD U2904 (.O(n1479), 
	.B2(n159), 
	.B1(\ram[56][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n552));
   AO22CHD U2905 (.O(n1480), 
	.B2(n159), 
	.B1(\ram[56][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n552));
   AO22CHD U2906 (.O(n1481), 
	.B2(n159), 
	.B1(\ram[56][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n552));
   AO22CHD U2907 (.O(n1482), 
	.B2(n159), 
	.B1(\ram[56][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n552));
   AO22CHD U2908 (.O(n1483), 
	.B2(n159), 
	.B1(\ram[56][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n552));
   AO22CHD U2909 (.O(n1484), 
	.B2(n159), 
	.B1(\ram[56][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n552));
   AO22CHD U2910 (.O(n1485), 
	.B2(n159), 
	.B1(\ram[56][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n552));
   AO22CHD U2911 (.O(n1486), 
	.B2(n159), 
	.B1(\ram[56][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n552));
   AO22CHD U2912 (.O(n1487), 
	.B2(n159), 
	.B1(\ram[56][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n552));
   AO22CHD U2913 (.O(n1488), 
	.B2(n159), 
	.B1(\ram[56][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n552));
   AO22CHD U2914 (.O(n1489), 
	.B2(n159), 
	.B1(\ram[56][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n552));
   AO22CHD U2915 (.O(n1490), 
	.B2(n159), 
	.B1(\ram[56][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n552));
   AO22CHD U2916 (.O(n1491), 
	.B2(n159), 
	.B1(\ram[56][13] ), 
	.A2(n21), 
	.A1(n552));
   AO22CHD U2917 (.O(n1492), 
	.B2(n159), 
	.B1(\ram[56][14] ), 
	.A2(n22), 
	.A1(n552));
   AO22CHD U2918 (.O(n1493), 
	.B2(n159), 
	.B1(\ram[56][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n552));
   AO22CHD U2919 (.O(n1494), 
	.B2(n161), 
	.B1(\ram[57][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n555));
   AO22CHD U2920 (.O(n1495), 
	.B2(n161), 
	.B1(\ram[57][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n555));
   AO22CHD U2921 (.O(n1496), 
	.B2(n161), 
	.B1(\ram[57][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n555));
   AO22CHD U2922 (.O(n1497), 
	.B2(n161), 
	.B1(\ram[57][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n555));
   AO22CHD U2923 (.O(n1498), 
	.B2(n161), 
	.B1(\ram[57][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n555));
   AO22CHD U2924 (.O(n1499), 
	.B2(n161), 
	.B1(\ram[57][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n555));
   AO22CHD U2925 (.O(n1500), 
	.B2(n161), 
	.B1(\ram[57][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n555));
   AO22CHD U2926 (.O(n1501), 
	.B2(n161), 
	.B1(\ram[57][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n555));
   AO22CHD U2927 (.O(n1502), 
	.B2(n161), 
	.B1(\ram[57][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n555));
   AO22CHD U2928 (.O(n1503), 
	.B2(n161), 
	.B1(\ram[57][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n555));
   AO22CHD U2929 (.O(n1504), 
	.B2(n161), 
	.B1(\ram[57][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n555));
   AO22CHD U2930 (.O(n1505), 
	.B2(n161), 
	.B1(\ram[57][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n555));
   AO22CHD U2931 (.O(n1506), 
	.B2(n161), 
	.B1(\ram[57][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n555));
   AO22CHD U2932 (.O(n1507), 
	.B2(n161), 
	.B1(\ram[57][13] ), 
	.A2(n21), 
	.A1(n555));
   AO22CHD U2933 (.O(n1508), 
	.B2(n161), 
	.B1(\ram[57][14] ), 
	.A2(n22), 
	.A1(n555));
   AO22CHD U2934 (.O(n1509), 
	.B2(n161), 
	.B1(\ram[57][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n555));
   AO22CHD U2935 (.O(n1510), 
	.B2(n163), 
	.B1(\ram[58][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n558));
   AO22CHD U2936 (.O(n1511), 
	.B2(n163), 
	.B1(\ram[58][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n558));
   AO22CHD U2937 (.O(n1512), 
	.B2(n163), 
	.B1(\ram[58][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n558));
   AO22CHD U2938 (.O(n1513), 
	.B2(n163), 
	.B1(\ram[58][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n558));
   AO22CHD U2939 (.O(n1514), 
	.B2(n163), 
	.B1(\ram[58][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n558));
   AO22CHD U2940 (.O(n1515), 
	.B2(n163), 
	.B1(\ram[58][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n558));
   AO22CHD U2941 (.O(n1516), 
	.B2(n163), 
	.B1(\ram[58][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n558));
   AO22CHD U2942 (.O(n1517), 
	.B2(n163), 
	.B1(\ram[58][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n558));
   AO22CHD U2943 (.O(n1518), 
	.B2(n163), 
	.B1(\ram[58][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n558));
   AO22CHD U2944 (.O(n1519), 
	.B2(n163), 
	.B1(\ram[58][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n558));
   AO22CHD U2945 (.O(n1520), 
	.B2(n163), 
	.B1(\ram[58][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n558));
   AO22CHD U2946 (.O(n1521), 
	.B2(n163), 
	.B1(\ram[58][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n558));
   AO22CHD U2947 (.O(n1522), 
	.B2(n163), 
	.B1(\ram[58][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n558));
   AO22CHD U2948 (.O(n1523), 
	.B2(n163), 
	.B1(\ram[58][13] ), 
	.A2(n21), 
	.A1(n558));
   AO22CHD U2949 (.O(n1524), 
	.B2(n163), 
	.B1(\ram[58][14] ), 
	.A2(n22), 
	.A1(n558));
   AO22CHD U2950 (.O(n1525), 
	.B2(n163), 
	.B1(\ram[58][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n558));
   AO22CHD U2951 (.O(n1526), 
	.B2(n165), 
	.B1(\ram[59][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n560));
   AO22CHD U2952 (.O(n1527), 
	.B2(n165), 
	.B1(\ram[59][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n560));
   AO22CHD U2953 (.O(n1528), 
	.B2(n165), 
	.B1(\ram[59][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n560));
   AO22CHD U2954 (.O(n1529), 
	.B2(n165), 
	.B1(\ram[59][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n560));
   AO22CHD U2955 (.O(n1530), 
	.B2(n165), 
	.B1(\ram[59][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n560));
   AO22CHD U2956 (.O(n1531), 
	.B2(n165), 
	.B1(\ram[59][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n560));
   AO22CHD U2957 (.O(n1532), 
	.B2(n165), 
	.B1(\ram[59][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n560));
   AO22CHD U2958 (.O(n1533), 
	.B2(n165), 
	.B1(\ram[59][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n560));
   AO22CHD U2959 (.O(n1534), 
	.B2(n165), 
	.B1(\ram[59][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n560));
   AO22CHD U2960 (.O(n1535), 
	.B2(n165), 
	.B1(\ram[59][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n560));
   AO22CHD U2961 (.O(n1536), 
	.B2(n165), 
	.B1(\ram[59][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n560));
   AO22CHD U2962 (.O(n1537), 
	.B2(n165), 
	.B1(\ram[59][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n560));
   AO22CHD U2963 (.O(n1538), 
	.B2(n165), 
	.B1(\ram[59][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n560));
   AO22CHD U2964 (.O(n1539), 
	.B2(n165), 
	.B1(\ram[59][13] ), 
	.A2(n21), 
	.A1(n560));
   AO22CHD U2965 (.O(n1540), 
	.B2(n165), 
	.B1(\ram[59][14] ), 
	.A2(n22), 
	.A1(n560));
   AO22CHD U2966 (.O(n1541), 
	.B2(n165), 
	.B1(\ram[59][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n560));
   AO22CHD U2967 (.O(n1542), 
	.B2(n167), 
	.B1(\ram[60][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n562));
   AO22CHD U2968 (.O(n1543), 
	.B2(n167), 
	.B1(\ram[60][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n562));
   AO22CHD U2969 (.O(n1544), 
	.B2(n167), 
	.B1(\ram[60][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n562));
   AO22CHD U2970 (.O(n1545), 
	.B2(n167), 
	.B1(\ram[60][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n562));
   AO22CHD U2971 (.O(n1546), 
	.B2(n167), 
	.B1(\ram[60][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n562));
   AO22CHD U2972 (.O(n1547), 
	.B2(n167), 
	.B1(\ram[60][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n562));
   AO22CHD U2973 (.O(n1548), 
	.B2(n167), 
	.B1(\ram[60][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n562));
   AO22CHD U2974 (.O(n1549), 
	.B2(n167), 
	.B1(\ram[60][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n562));
   AO22CHD U2975 (.O(n1550), 
	.B2(n167), 
	.B1(\ram[60][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n562));
   AO22CHD U2976 (.O(n1551), 
	.B2(n167), 
	.B1(\ram[60][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n562));
   AO22CHD U2977 (.O(n1552), 
	.B2(n167), 
	.B1(\ram[60][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n562));
   AO22CHD U2978 (.O(n1553), 
	.B2(n167), 
	.B1(\ram[60][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n562));
   AO22CHD U2979 (.O(n1554), 
	.B2(n167), 
	.B1(\ram[60][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n562));
   AO22CHD U2980 (.O(n1555), 
	.B2(n167), 
	.B1(\ram[60][13] ), 
	.A2(n21), 
	.A1(n562));
   AO22CHD U2981 (.O(n1556), 
	.B2(n167), 
	.B1(\ram[60][14] ), 
	.A2(n22), 
	.A1(n562));
   AO22CHD U2982 (.O(n1557), 
	.B2(n167), 
	.B1(\ram[60][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n562));
   AO22CHD U2983 (.O(n1558), 
	.B2(n169), 
	.B1(\ram[61][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n564));
   AO22CHD U2984 (.O(n1559), 
	.B2(n169), 
	.B1(\ram[61][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n564));
   AO22CHD U2985 (.O(n1560), 
	.B2(n169), 
	.B1(\ram[61][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n564));
   AO22CHD U2986 (.O(n1561), 
	.B2(n169), 
	.B1(\ram[61][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n564));
   AO22CHD U2987 (.O(n1562), 
	.B2(n169), 
	.B1(\ram[61][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n564));
   AO22CHD U2988 (.O(n1563), 
	.B2(n169), 
	.B1(\ram[61][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n564));
   AO22CHD U2989 (.O(n1564), 
	.B2(n169), 
	.B1(\ram[61][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n564));
   AO22CHD U2990 (.O(n1565), 
	.B2(n169), 
	.B1(\ram[61][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n564));
   AO22CHD U2991 (.O(n1566), 
	.B2(n169), 
	.B1(\ram[61][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n564));
   AO22CHD U2992 (.O(n1567), 
	.B2(n169), 
	.B1(\ram[61][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n564));
   AO22CHD U2993 (.O(n1568), 
	.B2(n169), 
	.B1(\ram[61][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n564));
   AO22CHD U2994 (.O(n1569), 
	.B2(n169), 
	.B1(\ram[61][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n564));
   AO22CHD U2995 (.O(n1570), 
	.B2(n169), 
	.B1(\ram[61][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n564));
   AO22CHD U2996 (.O(n1571), 
	.B2(n169), 
	.B1(\ram[61][13] ), 
	.A2(n21), 
	.A1(n564));
   AO22CHD U2997 (.O(n1572), 
	.B2(n169), 
	.B1(\ram[61][14] ), 
	.A2(n22), 
	.A1(n564));
   AO22CHD U2998 (.O(n1573), 
	.B2(n169), 
	.B1(\ram[61][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n564));
   AO22CHD U2999 (.O(n1574), 
	.B2(n171), 
	.B1(\ram[62][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n567));
   AO22CHD U3000 (.O(n1575), 
	.B2(n171), 
	.B1(\ram[62][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n567));
   AO22CHD U3001 (.O(n1576), 
	.B2(n171), 
	.B1(\ram[62][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n567));
   AO22CHD U3002 (.O(n1577), 
	.B2(n171), 
	.B1(\ram[62][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n567));
   AO22CHD U3003 (.O(n1578), 
	.B2(n171), 
	.B1(\ram[62][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n567));
   AO22CHD U3004 (.O(n1579), 
	.B2(n171), 
	.B1(\ram[62][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n567));
   AO22CHD U3005 (.O(n1580), 
	.B2(n171), 
	.B1(\ram[62][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n567));
   AO22CHD U3006 (.O(n1581), 
	.B2(n171), 
	.B1(\ram[62][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n567));
   AO22CHD U3007 (.O(n1582), 
	.B2(n171), 
	.B1(\ram[62][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n567));
   AO22CHD U3008 (.O(n1583), 
	.B2(n171), 
	.B1(\ram[62][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n567));
   AO22CHD U3009 (.O(n1584), 
	.B2(n171), 
	.B1(\ram[62][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n567));
   AO22CHD U3010 (.O(n1585), 
	.B2(n171), 
	.B1(\ram[62][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n567));
   AO22CHD U3011 (.O(n1586), 
	.B2(n171), 
	.B1(\ram[62][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n567));
   AO22CHD U3012 (.O(n1587), 
	.B2(n171), 
	.B1(\ram[62][13] ), 
	.A2(n21), 
	.A1(n567));
   AO22CHD U3013 (.O(n1588), 
	.B2(n171), 
	.B1(\ram[62][14] ), 
	.A2(n22), 
	.A1(n567));
   AO22CHD U3014 (.O(n1589), 
	.B2(n171), 
	.B1(\ram[62][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n567));
   AO22CHD U3015 (.O(n1590), 
	.B2(n173), 
	.B1(\ram[63][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n569));
   AO22CHD U3016 (.O(n1591), 
	.B2(n173), 
	.B1(\ram[63][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n569));
   AO22CHD U3017 (.O(n1592), 
	.B2(n173), 
	.B1(\ram[63][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n569));
   AO22CHD U3018 (.O(n1593), 
	.B2(n173), 
	.B1(\ram[63][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n569));
   AO22CHD U3019 (.O(n1594), 
	.B2(n173), 
	.B1(\ram[63][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n569));
   AO22CHD U3020 (.O(n1595), 
	.B2(n173), 
	.B1(\ram[63][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n569));
   AO22CHD U3021 (.O(n1596), 
	.B2(n173), 
	.B1(\ram[63][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n569));
   AO22CHD U3022 (.O(n1597), 
	.B2(n173), 
	.B1(\ram[63][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n569));
   AO22CHD U3023 (.O(n1598), 
	.B2(n173), 
	.B1(\ram[63][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n569));
   AO22CHD U3024 (.O(n1599), 
	.B2(n173), 
	.B1(\ram[63][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n569));
   AO22CHD U3025 (.O(n1600), 
	.B2(n173), 
	.B1(\ram[63][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n569));
   AO22CHD U3026 (.O(n1601), 
	.B2(n173), 
	.B1(\ram[63][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n569));
   AO22CHD U3027 (.O(n1602), 
	.B2(n173), 
	.B1(\ram[63][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n569));
   AO22CHD U3028 (.O(n1603), 
	.B2(n173), 
	.B1(\ram[63][13] ), 
	.A2(n21), 
	.A1(n569));
   AO22CHD U3029 (.O(n1604), 
	.B2(n173), 
	.B1(\ram[63][14] ), 
	.A2(n22), 
	.A1(n569));
   AO22CHD U3030 (.O(n1605), 
	.B2(n173), 
	.B1(\ram[63][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n569));
   AO22CHD U3031 (.O(n1606), 
	.B2(n176), 
	.B1(\ram[64][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n56));
   AO22CHD U3032 (.O(n1607), 
	.B2(n176), 
	.B1(\ram[64][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n56));
   AO22CHD U3033 (.O(n1608), 
	.B2(n176), 
	.B1(\ram[64][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n56));
   AO22CHD U3034 (.O(n1609), 
	.B2(n176), 
	.B1(\ram[64][3] ), 
	.A2(n11), 
	.A1(n56));
   AO22CHD U3035 (.O(n1610), 
	.B2(n176), 
	.B1(\ram[64][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n56));
   AO22CHD U3036 (.O(n1611), 
	.B2(n176), 
	.B1(\ram[64][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n56));
   AO22CHD U3037 (.O(n1612), 
	.B2(n176), 
	.B1(\ram[64][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n56));
   AO22CHD U3038 (.O(n1613), 
	.B2(n176), 
	.B1(\ram[64][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n56));
   AO22CHD U3039 (.O(n1614), 
	.B2(n176), 
	.B1(\ram[64][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n56));
   AO22CHD U3040 (.O(n1615), 
	.B2(n176), 
	.B1(\ram[64][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n56));
   AO22CHD U3041 (.O(n1616), 
	.B2(n176), 
	.B1(\ram[64][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n56));
   AO22CHD U3042 (.O(n1617), 
	.B2(n176), 
	.B1(\ram[64][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n56));
   AO22CHD U3043 (.O(n1618), 
	.B2(n176), 
	.B1(\ram[64][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n56));
   AO22CHD U3044 (.O(n1619), 
	.B2(n176), 
	.B1(\ram[64][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n56));
   AO22CHD U3045 (.O(n1620), 
	.B2(n176), 
	.B1(\ram[64][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n56));
   AO22CHD U3046 (.O(n1621), 
	.B2(n176), 
	.B1(\ram[64][15] ), 
	.A2(n23), 
	.A1(n56));
   AO22CHD U3047 (.O(n1622), 
	.B2(n179), 
	.B1(\ram[65][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n58));
   AO22CHD U3048 (.O(n1623), 
	.B2(n179), 
	.B1(\ram[65][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n58));
   AO22CHD U3049 (.O(n1624), 
	.B2(n179), 
	.B1(\ram[65][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n58));
   AO22CHD U3050 (.O(n1625), 
	.B2(n179), 
	.B1(\ram[65][3] ), 
	.A2(n11), 
	.A1(n58));
   AO22CHD U3051 (.O(n1626), 
	.B2(n179), 
	.B1(\ram[65][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n58));
   AO22CHD U3052 (.O(n1627), 
	.B2(n179), 
	.B1(\ram[65][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n58));
   AO22CHD U3053 (.O(n1628), 
	.B2(n179), 
	.B1(\ram[65][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n58));
   AO22CHD U3054 (.O(n1629), 
	.B2(n179), 
	.B1(\ram[65][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n58));
   AO22CHD U3055 (.O(n1630), 
	.B2(n179), 
	.B1(\ram[65][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n58));
   AO22CHD U3056 (.O(n1631), 
	.B2(n179), 
	.B1(\ram[65][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n58));
   AO22CHD U3057 (.O(n1632), 
	.B2(n179), 
	.B1(\ram[65][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n58));
   AO22CHD U3058 (.O(n1633), 
	.B2(n179), 
	.B1(\ram[65][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n58));
   AO22CHD U3059 (.O(n1634), 
	.B2(n179), 
	.B1(\ram[65][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n58));
   AO22CHD U3060 (.O(n1635), 
	.B2(n179), 
	.B1(\ram[65][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n58));
   AO22CHD U3061 (.O(n1636), 
	.B2(n179), 
	.B1(\ram[65][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n58));
   AO22CHD U3062 (.O(n1637), 
	.B2(n179), 
	.B1(\ram[65][15] ), 
	.A2(n23), 
	.A1(n58));
   AO22CHD U3063 (.O(n1638), 
	.B2(n181), 
	.B1(\ram[66][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n59));
   AO22CHD U3064 (.O(n1639), 
	.B2(n181), 
	.B1(\ram[66][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n59));
   AO22CHD U3065 (.O(n1640), 
	.B2(n181), 
	.B1(\ram[66][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n59));
   AO22CHD U3066 (.O(n1641), 
	.B2(n181), 
	.B1(\ram[66][3] ), 
	.A2(n11), 
	.A1(n59));
   AO22CHD U3067 (.O(n1642), 
	.B2(n181), 
	.B1(\ram[66][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n59));
   AO22CHD U3068 (.O(n1643), 
	.B2(n181), 
	.B1(\ram[66][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n59));
   AO22CHD U3069 (.O(n1644), 
	.B2(n181), 
	.B1(\ram[66][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n59));
   AO22CHD U3070 (.O(n1645), 
	.B2(n181), 
	.B1(\ram[66][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n59));
   AO22CHD U3071 (.O(n1646), 
	.B2(n181), 
	.B1(\ram[66][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n59));
   AO22CHD U3072 (.O(n1647), 
	.B2(n181), 
	.B1(\ram[66][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n59));
   AO22CHD U3073 (.O(n1648), 
	.B2(n181), 
	.B1(\ram[66][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n59));
   AO22CHD U3074 (.O(n1649), 
	.B2(n181), 
	.B1(\ram[66][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n59));
   AO22CHD U3075 (.O(n1650), 
	.B2(n181), 
	.B1(\ram[66][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n59));
   AO22CHD U3076 (.O(n1651), 
	.B2(n181), 
	.B1(\ram[66][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n59));
   AO22CHD U3077 (.O(n1652), 
	.B2(n181), 
	.B1(\ram[66][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n59));
   AO22CHD U3078 (.O(n1653), 
	.B2(n181), 
	.B1(\ram[66][15] ), 
	.A2(n23), 
	.A1(n59));
   AO22CHD U3079 (.O(n1654), 
	.B2(n183), 
	.B1(\ram[67][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n61));
   AO22CHD U3080 (.O(n1655), 
	.B2(n183), 
	.B1(\ram[67][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n61));
   AO22CHD U3081 (.O(n1656), 
	.B2(n183), 
	.B1(\ram[67][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n61));
   AO22CHD U3082 (.O(n1657), 
	.B2(n183), 
	.B1(\ram[67][3] ), 
	.A2(n11), 
	.A1(n61));
   AO22CHD U3083 (.O(n1658), 
	.B2(n183), 
	.B1(\ram[67][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n61));
   AO22CHD U3084 (.O(n1659), 
	.B2(n183), 
	.B1(\ram[67][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n61));
   AO22CHD U3085 (.O(n1660), 
	.B2(n183), 
	.B1(\ram[67][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n61));
   AO22CHD U3086 (.O(n1661), 
	.B2(n183), 
	.B1(\ram[67][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n61));
   AO22CHD U3087 (.O(n1662), 
	.B2(n183), 
	.B1(\ram[67][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n61));
   AO22CHD U3088 (.O(n1663), 
	.B2(n183), 
	.B1(\ram[67][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n61));
   AO22CHD U3089 (.O(n1664), 
	.B2(n183), 
	.B1(\ram[67][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n61));
   AO22CHD U3090 (.O(n1665), 
	.B2(n183), 
	.B1(\ram[67][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n61));
   AO22CHD U3091 (.O(n1666), 
	.B2(n183), 
	.B1(\ram[67][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n61));
   AO22CHD U3092 (.O(n1667), 
	.B2(n183), 
	.B1(\ram[67][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n61));
   AO22CHD U3093 (.O(n1668), 
	.B2(n183), 
	.B1(\ram[67][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n61));
   AO22CHD U3094 (.O(n1669), 
	.B2(n183), 
	.B1(\ram[67][15] ), 
	.A2(n23), 
	.A1(n61));
   AO22CHD U3095 (.O(n1670), 
	.B2(n185), 
	.B1(\ram[68][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n62));
   AO22CHD U3096 (.O(n1671), 
	.B2(n185), 
	.B1(\ram[68][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n62));
   AO22CHD U3097 (.O(n1672), 
	.B2(n185), 
	.B1(\ram[68][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n62));
   AO22CHD U3098 (.O(n1673), 
	.B2(n185), 
	.B1(\ram[68][3] ), 
	.A2(n11), 
	.A1(n62));
   AO22CHD U3099 (.O(n1674), 
	.B2(n185), 
	.B1(\ram[68][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n62));
   AO22CHD U3100 (.O(n1675), 
	.B2(n185), 
	.B1(\ram[68][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n62));
   AO22CHD U3101 (.O(n1676), 
	.B2(n185), 
	.B1(\ram[68][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n62));
   AO22CHD U3102 (.O(n1677), 
	.B2(n185), 
	.B1(\ram[68][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n62));
   AO22CHD U3103 (.O(n1678), 
	.B2(n185), 
	.B1(\ram[68][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n62));
   AO22CHD U3104 (.O(n1679), 
	.B2(n185), 
	.B1(\ram[68][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n62));
   AO22CHD U3105 (.O(n1680), 
	.B2(n185), 
	.B1(\ram[68][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n62));
   AO22CHD U3106 (.O(n1681), 
	.B2(n185), 
	.B1(\ram[68][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n62));
   AO22CHD U3107 (.O(n1682), 
	.B2(n185), 
	.B1(\ram[68][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n62));
   AO22CHD U3108 (.O(n1683), 
	.B2(n185), 
	.B1(\ram[68][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n62));
   AO22CHD U3109 (.O(n1684), 
	.B2(n185), 
	.B1(\ram[68][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n62));
   AO22CHD U3110 (.O(n1685), 
	.B2(n185), 
	.B1(\ram[68][15] ), 
	.A2(n23), 
	.A1(n62));
   AO22CHD U3111 (.O(n1686), 
	.B2(n187), 
	.B1(\ram[69][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n64));
   AO22CHD U3112 (.O(n1687), 
	.B2(n187), 
	.B1(\ram[69][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n64));
   AO22CHD U3113 (.O(n1688), 
	.B2(n187), 
	.B1(\ram[69][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n64));
   AO22CHD U3114 (.O(n1689), 
	.B2(n187), 
	.B1(\ram[69][3] ), 
	.A2(n11), 
	.A1(n64));
   AO22CHD U3115 (.O(n1690), 
	.B2(n187), 
	.B1(\ram[69][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n64));
   AO22CHD U3116 (.O(n1691), 
	.B2(n187), 
	.B1(\ram[69][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n64));
   AO22CHD U3117 (.O(n1692), 
	.B2(n187), 
	.B1(\ram[69][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n64));
   AO22CHD U3118 (.O(n1693), 
	.B2(n187), 
	.B1(\ram[69][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n64));
   AO22CHD U3119 (.O(n1694), 
	.B2(n187), 
	.B1(\ram[69][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n64));
   AO22CHD U3120 (.O(n1695), 
	.B2(n187), 
	.B1(\ram[69][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n64));
   AO22CHD U3121 (.O(n1696), 
	.B2(n187), 
	.B1(\ram[69][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n64));
   AO22CHD U3122 (.O(n1697), 
	.B2(n187), 
	.B1(\ram[69][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n64));
   AO22CHD U3123 (.O(n1698), 
	.B2(n187), 
	.B1(\ram[69][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n64));
   AO22CHD U3124 (.O(n1699), 
	.B2(n187), 
	.B1(\ram[69][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n64));
   AO22CHD U3125 (.O(n1700), 
	.B2(n187), 
	.B1(\ram[69][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n64));
   AO22CHD U3126 (.O(n1701), 
	.B2(n187), 
	.B1(\ram[69][15] ), 
	.A2(n23), 
	.A1(n64));
   AO22CHD U3127 (.O(n1702), 
	.B2(n189), 
	.B1(\ram[70][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n65));
   AO22CHD U3128 (.O(n1703), 
	.B2(n189), 
	.B1(\ram[70][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n65));
   AO22CHD U3129 (.O(n1704), 
	.B2(n189), 
	.B1(\ram[70][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n65));
   AO22CHD U3130 (.O(n1705), 
	.B2(n189), 
	.B1(\ram[70][3] ), 
	.A2(n11), 
	.A1(n65));
   AO22CHD U3131 (.O(n1706), 
	.B2(n189), 
	.B1(\ram[70][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n65));
   AO22CHD U3132 (.O(n1707), 
	.B2(n189), 
	.B1(\ram[70][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n65));
   AO22CHD U3133 (.O(n1708), 
	.B2(n189), 
	.B1(\ram[70][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n65));
   AO22CHD U3134 (.O(n1709), 
	.B2(n189), 
	.B1(\ram[70][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n65));
   AO22CHD U3135 (.O(n1710), 
	.B2(n189), 
	.B1(\ram[70][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n65));
   AO22CHD U3136 (.O(n1711), 
	.B2(n189), 
	.B1(\ram[70][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n65));
   AO22CHD U3137 (.O(n1712), 
	.B2(n189), 
	.B1(\ram[70][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n65));
   AO22CHD U3138 (.O(n1713), 
	.B2(n189), 
	.B1(\ram[70][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n65));
   AO22CHD U3139 (.O(n1714), 
	.B2(n189), 
	.B1(\ram[70][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n65));
   AO22CHD U3140 (.O(n1715), 
	.B2(n189), 
	.B1(\ram[70][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n65));
   AO22CHD U3141 (.O(n1716), 
	.B2(n189), 
	.B1(\ram[70][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n65));
   AO22CHD U3142 (.O(n1717), 
	.B2(n189), 
	.B1(\ram[70][15] ), 
	.A2(n23), 
	.A1(n65));
   AO22CHD U3143 (.O(n1718), 
	.B2(n191), 
	.B1(\ram[71][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n67));
   AO22CHD U3144 (.O(n1719), 
	.B2(n191), 
	.B1(\ram[71][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n67));
   AO22CHD U3145 (.O(n1720), 
	.B2(n191), 
	.B1(\ram[71][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n67));
   AO22CHD U3146 (.O(n1721), 
	.B2(n191), 
	.B1(\ram[71][3] ), 
	.A2(n11), 
	.A1(n67));
   AO22CHD U3147 (.O(n1722), 
	.B2(n191), 
	.B1(\ram[71][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n67));
   AO22CHD U3148 (.O(n1723), 
	.B2(n191), 
	.B1(\ram[71][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n67));
   AO22CHD U3149 (.O(n1724), 
	.B2(n191), 
	.B1(\ram[71][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n67));
   AO22CHD U3150 (.O(n1725), 
	.B2(n191), 
	.B1(\ram[71][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n67));
   AO22CHD U3151 (.O(n1726), 
	.B2(n191), 
	.B1(\ram[71][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n67));
   AO22CHD U3152 (.O(n1727), 
	.B2(n191), 
	.B1(\ram[71][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n67));
   AO22CHD U3153 (.O(n1728), 
	.B2(n191), 
	.B1(\ram[71][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n67));
   AO22CHD U3154 (.O(n1729), 
	.B2(n191), 
	.B1(\ram[71][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n67));
   AO22CHD U3155 (.O(n1730), 
	.B2(n191), 
	.B1(\ram[71][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n67));
   AO22CHD U3156 (.O(n1731), 
	.B2(n191), 
	.B1(\ram[71][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n67));
   AO22CHD U3157 (.O(n1732), 
	.B2(n191), 
	.B1(\ram[71][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n67));
   AO22CHD U3158 (.O(n1733), 
	.B2(n191), 
	.B1(\ram[71][15] ), 
	.A2(n23), 
	.A1(n67));
   AO22CHD U3159 (.O(n1734), 
	.B2(n193), 
	.B1(\ram[72][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n68));
   AO22CHD U3160 (.O(n1735), 
	.B2(n193), 
	.B1(\ram[72][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n68));
   AO22CHD U3161 (.O(n1736), 
	.B2(n193), 
	.B1(\ram[72][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n68));
   AO22CHD U3162 (.O(n1737), 
	.B2(n193), 
	.B1(\ram[72][3] ), 
	.A2(n11), 
	.A1(n68));
   AO22CHD U3163 (.O(n1738), 
	.B2(n193), 
	.B1(\ram[72][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n68));
   AO22CHD U3164 (.O(n1739), 
	.B2(n193), 
	.B1(\ram[72][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n68));
   AO22CHD U3165 (.O(n1740), 
	.B2(n193), 
	.B1(\ram[72][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n68));
   AO22CHD U3166 (.O(n1741), 
	.B2(n193), 
	.B1(\ram[72][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n68));
   AO22CHD U3167 (.O(n1742), 
	.B2(n193), 
	.B1(\ram[72][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n68));
   AO22CHD U3168 (.O(n1743), 
	.B2(n193), 
	.B1(\ram[72][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n68));
   AO22CHD U3169 (.O(n1744), 
	.B2(n193), 
	.B1(\ram[72][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n68));
   AO22CHD U3170 (.O(n1745), 
	.B2(n193), 
	.B1(\ram[72][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n68));
   AO22CHD U3171 (.O(n1746), 
	.B2(n193), 
	.B1(\ram[72][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n68));
   AO22CHD U3172 (.O(n1747), 
	.B2(n193), 
	.B1(\ram[72][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n68));
   AO22CHD U3173 (.O(n1748), 
	.B2(n193), 
	.B1(\ram[72][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n68));
   AO22CHD U3174 (.O(n1749), 
	.B2(n193), 
	.B1(\ram[72][15] ), 
	.A2(n23), 
	.A1(n68));
   AO22CHD U3175 (.O(n1750), 
	.B2(n195), 
	.B1(\ram[73][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n70));
   AO22CHD U3176 (.O(n1751), 
	.B2(n195), 
	.B1(\ram[73][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n70));
   AO22CHD U3177 (.O(n1752), 
	.B2(n195), 
	.B1(\ram[73][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n70));
   AO22CHD U3178 (.O(n1753), 
	.B2(n195), 
	.B1(\ram[73][3] ), 
	.A2(n11), 
	.A1(n70));
   AO22CHD U3179 (.O(n1754), 
	.B2(n195), 
	.B1(\ram[73][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n70));
   AO22CHD U3180 (.O(n1755), 
	.B2(n195), 
	.B1(\ram[73][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n70));
   AO22CHD U3181 (.O(n1756), 
	.B2(n195), 
	.B1(\ram[73][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n70));
   AO22CHD U3182 (.O(n1757), 
	.B2(n195), 
	.B1(\ram[73][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n70));
   AO22CHD U3183 (.O(n1758), 
	.B2(n195), 
	.B1(\ram[73][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n70));
   AO22CHD U3184 (.O(n1759), 
	.B2(n195), 
	.B1(\ram[73][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n70));
   AO22CHD U3185 (.O(n1760), 
	.B2(n195), 
	.B1(\ram[73][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n70));
   AO22CHD U3186 (.O(n1761), 
	.B2(n195), 
	.B1(\ram[73][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n70));
   AO22CHD U3187 (.O(n1762), 
	.B2(n195), 
	.B1(\ram[73][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n70));
   AO22CHD U3188 (.O(n1763), 
	.B2(n195), 
	.B1(\ram[73][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n70));
   AO22CHD U3189 (.O(n1764), 
	.B2(n195), 
	.B1(\ram[73][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n70));
   AO22CHD U3190 (.O(n1765), 
	.B2(n195), 
	.B1(\ram[73][15] ), 
	.A2(n23), 
	.A1(n70));
   AO22CHD U3191 (.O(n1766), 
	.B2(n197), 
	.B1(\ram[74][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n73));
   AO22CHD U3192 (.O(n1767), 
	.B2(n197), 
	.B1(\ram[74][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n73));
   AO22CHD U3193 (.O(n1768), 
	.B2(n197), 
	.B1(\ram[74][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n73));
   AO22CHD U3194 (.O(n1769), 
	.B2(n197), 
	.B1(\ram[74][3] ), 
	.A2(n11), 
	.A1(n73));
   AO22CHD U3195 (.O(n1770), 
	.B2(n197), 
	.B1(\ram[74][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n73));
   AO22CHD U3196 (.O(n1771), 
	.B2(n197), 
	.B1(\ram[74][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n73));
   AO22CHD U3197 (.O(n1772), 
	.B2(n197), 
	.B1(\ram[74][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n73));
   AO22CHD U3198 (.O(n1773), 
	.B2(n197), 
	.B1(\ram[74][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n73));
   AO22CHD U3199 (.O(n1774), 
	.B2(n197), 
	.B1(\ram[74][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n73));
   AO22CHD U3200 (.O(n1775), 
	.B2(n197), 
	.B1(\ram[74][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n73));
   AO22CHD U3201 (.O(n1776), 
	.B2(n197), 
	.B1(\ram[74][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n73));
   AO22CHD U3202 (.O(n1777), 
	.B2(n197), 
	.B1(\ram[74][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n73));
   AO22CHD U3203 (.O(n1778), 
	.B2(n197), 
	.B1(\ram[74][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n73));
   AO22CHD U3204 (.O(n1779), 
	.B2(n197), 
	.B1(\ram[74][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n73));
   AO22CHD U3205 (.O(n1780), 
	.B2(n197), 
	.B1(\ram[74][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n73));
   AO22CHD U3206 (.O(n1781), 
	.B2(n197), 
	.B1(\ram[74][15] ), 
	.A2(n23), 
	.A1(n73));
   AO22CHD U3207 (.O(n1782), 
	.B2(n199), 
	.B1(\ram[75][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n75));
   AO22CHD U3208 (.O(n1783), 
	.B2(n199), 
	.B1(\ram[75][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n75));
   AO22CHD U3209 (.O(n1784), 
	.B2(n199), 
	.B1(\ram[75][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n75));
   AO22CHD U3210 (.O(n1785), 
	.B2(n199), 
	.B1(\ram[75][3] ), 
	.A2(n11), 
	.A1(n75));
   AO22CHD U3211 (.O(n1786), 
	.B2(n199), 
	.B1(\ram[75][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n75));
   AO22CHD U3212 (.O(n1787), 
	.B2(n199), 
	.B1(\ram[75][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n75));
   AO22CHD U3213 (.O(n1788), 
	.B2(n199), 
	.B1(\ram[75][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n75));
   AO22CHD U3214 (.O(n1789), 
	.B2(n199), 
	.B1(\ram[75][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n75));
   AO22CHD U3215 (.O(n1790), 
	.B2(n199), 
	.B1(\ram[75][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n75));
   AO22CHD U3216 (.O(n1791), 
	.B2(n199), 
	.B1(\ram[75][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n75));
   AO22CHD U3217 (.O(n1792), 
	.B2(n199), 
	.B1(\ram[75][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n75));
   AO22CHD U3218 (.O(n1793), 
	.B2(n199), 
	.B1(\ram[75][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n75));
   AO22CHD U3219 (.O(n1794), 
	.B2(n199), 
	.B1(\ram[75][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n75));
   AO22CHD U3220 (.O(n1795), 
	.B2(n199), 
	.B1(\ram[75][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n75));
   AO22CHD U3221 (.O(n1796), 
	.B2(n199), 
	.B1(\ram[75][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n75));
   AO22CHD U3222 (.O(n1797), 
	.B2(n199), 
	.B1(\ram[75][15] ), 
	.A2(n23), 
	.A1(n75));
   AO22CHD U3223 (.O(n1798), 
	.B2(n201), 
	.B1(\ram[76][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n76));
   AO22CHD U3224 (.O(n1799), 
	.B2(n201), 
	.B1(\ram[76][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n76));
   AO22CHD U3225 (.O(n1800), 
	.B2(n201), 
	.B1(\ram[76][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n76));
   AO22CHD U3226 (.O(n1801), 
	.B2(n201), 
	.B1(\ram[76][3] ), 
	.A2(n11), 
	.A1(n76));
   AO22CHD U3227 (.O(n1802), 
	.B2(n201), 
	.B1(\ram[76][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n76));
   AO22CHD U3228 (.O(n1803), 
	.B2(n201), 
	.B1(\ram[76][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n76));
   AO22CHD U3229 (.O(n1804), 
	.B2(n201), 
	.B1(\ram[76][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n76));
   AO22CHD U3230 (.O(n1805), 
	.B2(n201), 
	.B1(\ram[76][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n76));
   AO22CHD U3231 (.O(n1806), 
	.B2(n201), 
	.B1(\ram[76][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n76));
   AO22CHD U3232 (.O(n1807), 
	.B2(n201), 
	.B1(\ram[76][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n76));
   AO22CHD U3233 (.O(n1808), 
	.B2(n201), 
	.B1(\ram[76][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n76));
   AO22CHD U3234 (.O(n1809), 
	.B2(n201), 
	.B1(\ram[76][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n76));
   AO22CHD U3235 (.O(n1810), 
	.B2(n201), 
	.B1(\ram[76][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n76));
   AO22CHD U3236 (.O(n1811), 
	.B2(n201), 
	.B1(\ram[76][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n76));
   AO22CHD U3237 (.O(n1812), 
	.B2(n201), 
	.B1(\ram[76][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n76));
   AO22CHD U3238 (.O(n1813), 
	.B2(n201), 
	.B1(\ram[76][15] ), 
	.A2(n23), 
	.A1(n76));
   AO22CHD U3239 (.O(n1814), 
	.B2(n203), 
	.B1(\ram[77][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n78));
   AO22CHD U3240 (.O(n1815), 
	.B2(n203), 
	.B1(\ram[77][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n78));
   AO22CHD U3241 (.O(n1816), 
	.B2(n203), 
	.B1(\ram[77][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n78));
   AO22CHD U3242 (.O(n1817), 
	.B2(n203), 
	.B1(\ram[77][3] ), 
	.A2(n11), 
	.A1(n78));
   AO22CHD U3243 (.O(n1818), 
	.B2(n203), 
	.B1(\ram[77][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n78));
   AO22CHD U3244 (.O(n1819), 
	.B2(n203), 
	.B1(\ram[77][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n78));
   AO22CHD U3245 (.O(n1820), 
	.B2(n203), 
	.B1(\ram[77][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n78));
   AO22CHD U3246 (.O(n1821), 
	.B2(n203), 
	.B1(\ram[77][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n78));
   AO22CHD U3247 (.O(n1822), 
	.B2(n203), 
	.B1(\ram[77][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n78));
   AO22CHD U3248 (.O(n1823), 
	.B2(n203), 
	.B1(\ram[77][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n78));
   AO22CHD U3249 (.O(n1824), 
	.B2(n203), 
	.B1(\ram[77][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n78));
   AO22CHD U3250 (.O(n1825), 
	.B2(n203), 
	.B1(\ram[77][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n78));
   AO22CHD U3251 (.O(n1826), 
	.B2(n203), 
	.B1(\ram[77][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n78));
   AO22CHD U3252 (.O(n1827), 
	.B2(n203), 
	.B1(\ram[77][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n78));
   AO22CHD U3253 (.O(n1828), 
	.B2(n203), 
	.B1(\ram[77][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n78));
   AO22CHD U3254 (.O(n1829), 
	.B2(n203), 
	.B1(\ram[77][15] ), 
	.A2(n23), 
	.A1(n78));
   AO22CHD U3255 (.O(n1830), 
	.B2(n205), 
	.B1(\ram[78][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n80));
   AO22CHD U3256 (.O(n1831), 
	.B2(n205), 
	.B1(\ram[78][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n80));
   AO22CHD U3257 (.O(n1832), 
	.B2(n205), 
	.B1(\ram[78][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n80));
   AO22CHD U3258 (.O(n1833), 
	.B2(n205), 
	.B1(\ram[78][3] ), 
	.A2(n11), 
	.A1(n80));
   AO22CHD U3259 (.O(n1834), 
	.B2(n205), 
	.B1(\ram[78][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n80));
   AO22CHD U3260 (.O(n1835), 
	.B2(n205), 
	.B1(\ram[78][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n80));
   AO22CHD U3261 (.O(n1836), 
	.B2(n205), 
	.B1(\ram[78][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n80));
   AO22CHD U3262 (.O(n1837), 
	.B2(n205), 
	.B1(\ram[78][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n80));
   AO22CHD U3263 (.O(n1838), 
	.B2(n205), 
	.B1(\ram[78][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n80));
   AO22CHD U3264 (.O(n1839), 
	.B2(n205), 
	.B1(\ram[78][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n80));
   AO22CHD U3265 (.O(n1840), 
	.B2(n205), 
	.B1(\ram[78][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n80));
   AO22CHD U3266 (.O(n1841), 
	.B2(n205), 
	.B1(\ram[78][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n80));
   AO22CHD U3267 (.O(n1842), 
	.B2(n205), 
	.B1(\ram[78][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n80));
   AO22CHD U3268 (.O(n1843), 
	.B2(n205), 
	.B1(\ram[78][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n80));
   AO22CHD U3269 (.O(n1844), 
	.B2(n205), 
	.B1(\ram[78][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n80));
   AO22CHD U3270 (.O(n1845), 
	.B2(n205), 
	.B1(\ram[78][15] ), 
	.A2(n23), 
	.A1(n80));
   AO22CHD U3271 (.O(n1846), 
	.B2(n207), 
	.B1(\ram[79][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n82));
   AO22CHD U3272 (.O(n1847), 
	.B2(n207), 
	.B1(\ram[79][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n82));
   AO22CHD U3273 (.O(n1848), 
	.B2(n207), 
	.B1(\ram[79][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n82));
   AO22CHD U3274 (.O(n1849), 
	.B2(n207), 
	.B1(\ram[79][3] ), 
	.A2(n11), 
	.A1(n82));
   AO22CHD U3275 (.O(n1850), 
	.B2(n207), 
	.B1(\ram[79][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n82));
   AO22CHD U3276 (.O(n1851), 
	.B2(n207), 
	.B1(\ram[79][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n82));
   AO22CHD U3277 (.O(n1852), 
	.B2(n207), 
	.B1(\ram[79][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n82));
   AO22CHD U3278 (.O(n1853), 
	.B2(n207), 
	.B1(\ram[79][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n82));
   AO22CHD U3279 (.O(n1854), 
	.B2(n207), 
	.B1(\ram[79][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n82));
   AO22CHD U3280 (.O(n1855), 
	.B2(n207), 
	.B1(\ram[79][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n82));
   AO22CHD U3281 (.O(n1856), 
	.B2(n207), 
	.B1(\ram[79][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n82));
   AO22CHD U3282 (.O(n1857), 
	.B2(n207), 
	.B1(\ram[79][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n82));
   AO22CHD U3283 (.O(n1858), 
	.B2(n207), 
	.B1(\ram[79][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n82));
   AO22CHD U3284 (.O(n1859), 
	.B2(n207), 
	.B1(\ram[79][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n82));
   AO22CHD U3285 (.O(n1860), 
	.B2(n207), 
	.B1(\ram[79][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n82));
   AO22CHD U3286 (.O(n1861), 
	.B2(n207), 
	.B1(\ram[79][15] ), 
	.A2(n23), 
	.A1(n82));
   AO22CHD U3287 (.O(n1862), 
	.B2(n210), 
	.B1(\ram[80][0] ), 
	.A2(n6), 
	.A1(n84));
   AO22CHD U3288 (.O(n1863), 
	.B2(n210), 
	.B1(\ram[80][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n84));
   AO22CHD U3289 (.O(n1864), 
	.B2(n210), 
	.B1(\ram[80][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n84));
   AO22CHD U3290 (.O(n1865), 
	.B2(n210), 
	.B1(\ram[80][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n84));
   AO22CHD U3291 (.O(n1866), 
	.B2(n210), 
	.B1(\ram[80][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n84));
   AO22CHD U3292 (.O(n1867), 
	.B2(n210), 
	.B1(\ram[80][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n84));
   AO22CHD U3293 (.O(n1868), 
	.B2(n210), 
	.B1(\ram[80][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n84));
   AO22CHD U3294 (.O(n1869), 
	.B2(n210), 
	.B1(\ram[80][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n84));
   AO22CHD U3295 (.O(n1870), 
	.B2(n210), 
	.B1(\ram[80][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n84));
   AO22CHD U3296 (.O(n1871), 
	.B2(n210), 
	.B1(\ram[80][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n84));
   AO22CHD U3297 (.O(n1872), 
	.B2(n210), 
	.B1(\ram[80][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n84));
   AO22CHD U3298 (.O(n1873), 
	.B2(n210), 
	.B1(\ram[80][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n84));
   AO22CHD U3299 (.O(n1874), 
	.B2(n210), 
	.B1(\ram[80][12] ), 
	.A2(n20), 
	.A1(n84));
   AO22CHD U3300 (.O(n1875), 
	.B2(n210), 
	.B1(\ram[80][13] ), 
	.A2(n21), 
	.A1(n84));
   AO22CHD U3301 (.O(n1876), 
	.B2(n210), 
	.B1(\ram[80][14] ), 
	.A2(n22), 
	.A1(n84));
   AO22CHD U3302 (.O(n1877), 
	.B2(n210), 
	.B1(\ram[80][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n84));
   AO22CHD U3303 (.O(n1878), 
	.B2(n213), 
	.B1(\ram[81][0] ), 
	.A2(n6), 
	.A1(n86));
   AO22CHD U3304 (.O(n1879), 
	.B2(n213), 
	.B1(\ram[81][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n86));
   AO22CHD U3305 (.O(n1880), 
	.B2(n213), 
	.B1(\ram[81][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n86));
   AO22CHD U3306 (.O(n1881), 
	.B2(n213), 
	.B1(\ram[81][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n86));
   AO22CHD U3307 (.O(n1882), 
	.B2(n213), 
	.B1(\ram[81][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n86));
   AO22CHD U3308 (.O(n1883), 
	.B2(n213), 
	.B1(\ram[81][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n86));
   AO22CHD U3309 (.O(n1884), 
	.B2(n213), 
	.B1(\ram[81][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n86));
   AO22CHD U3310 (.O(n1885), 
	.B2(n213), 
	.B1(\ram[81][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n86));
   AO22CHD U3311 (.O(n1886), 
	.B2(n213), 
	.B1(\ram[81][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n86));
   AO22CHD U3312 (.O(n1887), 
	.B2(n213), 
	.B1(\ram[81][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n86));
   AO22CHD U3313 (.O(n1888), 
	.B2(n213), 
	.B1(\ram[81][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n86));
   AO22CHD U3314 (.O(n1889), 
	.B2(n213), 
	.B1(\ram[81][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n86));
   AO22CHD U3315 (.O(n1890), 
	.B2(n213), 
	.B1(\ram[81][12] ), 
	.A2(n20), 
	.A1(n86));
   AO22CHD U3316 (.O(n1891), 
	.B2(n213), 
	.B1(\ram[81][13] ), 
	.A2(n21), 
	.A1(n86));
   AO22CHD U3317 (.O(n1892), 
	.B2(n213), 
	.B1(\ram[81][14] ), 
	.A2(n22), 
	.A1(n86));
   AO22CHD U3318 (.O(n1893), 
	.B2(n213), 
	.B1(\ram[81][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n86));
   AO22CHD U3319 (.O(n1894), 
	.B2(n215), 
	.B1(\ram[82][0] ), 
	.A2(n6), 
	.A1(n88));
   AO22CHD U3320 (.O(n1895), 
	.B2(n215), 
	.B1(\ram[82][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n88));
   AO22CHD U3321 (.O(n1896), 
	.B2(n215), 
	.B1(\ram[82][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n88));
   AO22CHD U3322 (.O(n1897), 
	.B2(n215), 
	.B1(\ram[82][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n88));
   AO22CHD U3323 (.O(n1898), 
	.B2(n215), 
	.B1(\ram[82][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n88));
   AO22CHD U3324 (.O(n1899), 
	.B2(n215), 
	.B1(\ram[82][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n88));
   AO22CHD U3325 (.O(n1900), 
	.B2(n215), 
	.B1(\ram[82][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n88));
   AO22CHD U3326 (.O(n1901), 
	.B2(n215), 
	.B1(\ram[82][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n88));
   AO22CHD U3327 (.O(n1902), 
	.B2(n215), 
	.B1(\ram[82][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n88));
   AO22CHD U3328 (.O(n1903), 
	.B2(n215), 
	.B1(\ram[82][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n88));
   AO22CHD U3329 (.O(n1904), 
	.B2(n215), 
	.B1(\ram[82][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n88));
   AO22CHD U3330 (.O(n1905), 
	.B2(n215), 
	.B1(\ram[82][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n88));
   AO22CHD U3331 (.O(n1906), 
	.B2(n215), 
	.B1(\ram[82][12] ), 
	.A2(n20), 
	.A1(n88));
   AO22CHD U3332 (.O(n1907), 
	.B2(n215), 
	.B1(\ram[82][13] ), 
	.A2(n21), 
	.A1(n88));
   AO22CHD U3333 (.O(n1908), 
	.B2(n215), 
	.B1(\ram[82][14] ), 
	.A2(n22), 
	.A1(n88));
   AO22CHD U3334 (.O(n1909), 
	.B2(n215), 
	.B1(\ram[82][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n88));
   AO22CHD U3335 (.O(n1910), 
	.B2(n217), 
	.B1(\ram[83][0] ), 
	.A2(n6), 
	.A1(n90));
   AO22CHD U3336 (.O(n1911), 
	.B2(n217), 
	.B1(\ram[83][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n90));
   AO22CHD U3337 (.O(n1912), 
	.B2(n217), 
	.B1(\ram[83][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n90));
   AO22CHD U3338 (.O(n1913), 
	.B2(n217), 
	.B1(\ram[83][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n90));
   AO22CHD U3339 (.O(n1914), 
	.B2(n217), 
	.B1(\ram[83][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n90));
   AO22CHD U3340 (.O(n1915), 
	.B2(n217), 
	.B1(\ram[83][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n90));
   AO22CHD U3341 (.O(n1916), 
	.B2(n217), 
	.B1(\ram[83][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n90));
   AO22CHD U3342 (.O(n1917), 
	.B2(n217), 
	.B1(\ram[83][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n90));
   AO22CHD U3343 (.O(n1918), 
	.B2(n217), 
	.B1(\ram[83][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n90));
   AO22CHD U3344 (.O(n1919), 
	.B2(n217), 
	.B1(\ram[83][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n90));
   AO22CHD U3345 (.O(n1920), 
	.B2(n217), 
	.B1(\ram[83][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n90));
   AO22CHD U3346 (.O(n1921), 
	.B2(n217), 
	.B1(\ram[83][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n90));
   AO22CHD U3347 (.O(n1922), 
	.B2(n217), 
	.B1(\ram[83][12] ), 
	.A2(n20), 
	.A1(n90));
   AO22CHD U3348 (.O(n1923), 
	.B2(n217), 
	.B1(\ram[83][13] ), 
	.A2(n21), 
	.A1(n90));
   AO22CHD U3349 (.O(n1924), 
	.B2(n217), 
	.B1(\ram[83][14] ), 
	.A2(n22), 
	.A1(n90));
   AO22CHD U3350 (.O(n1925), 
	.B2(n217), 
	.B1(\ram[83][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n90));
   AO22CHD U3351 (.O(n1926), 
	.B2(n219), 
	.B1(\ram[84][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n92));
   AO22CHD U3352 (.O(n1927), 
	.B2(n219), 
	.B1(\ram[84][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n92));
   AO22CHD U3353 (.O(n1928), 
	.B2(n219), 
	.B1(\ram[84][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n92));
   AO22CHD U3354 (.O(n1929), 
	.B2(n219), 
	.B1(\ram[84][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n92));
   AO22CHD U3355 (.O(n1930), 
	.B2(n219), 
	.B1(\ram[84][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n92));
   AO22CHD U3356 (.O(n1931), 
	.B2(n219), 
	.B1(\ram[84][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n92));
   AO22CHD U3357 (.O(n1932), 
	.B2(n219), 
	.B1(\ram[84][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n92));
   AO22CHD U3358 (.O(n1933), 
	.B2(n219), 
	.B1(\ram[84][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n92));
   AO22CHD U3359 (.O(n1934), 
	.B2(n219), 
	.B1(\ram[84][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n92));
   AO22CHD U3360 (.O(n1935), 
	.B2(n219), 
	.B1(\ram[84][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n92));
   AO22CHD U3361 (.O(n1936), 
	.B2(n219), 
	.B1(\ram[84][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n92));
   AO22CHD U3362 (.O(n1937), 
	.B2(n219), 
	.B1(\ram[84][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n92));
   AO22CHD U3363 (.O(n1938), 
	.B2(n219), 
	.B1(\ram[84][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n92));
   AO22CHD U3364 (.O(n1939), 
	.B2(n219), 
	.B1(\ram[84][13] ), 
	.A2(n21), 
	.A1(n92));
   AO22CHD U3365 (.O(n1940), 
	.B2(n219), 
	.B1(\ram[84][14] ), 
	.A2(n22), 
	.A1(n92));
   AO22CHD U3366 (.O(n1941), 
	.B2(n219), 
	.B1(\ram[84][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n92));
   AO22CHD U3367 (.O(n1942), 
	.B2(n221), 
	.B1(\ram[85][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n94));
   AO22CHD U3368 (.O(n1943), 
	.B2(n221), 
	.B1(\ram[85][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n94));
   AO22CHD U3369 (.O(n1944), 
	.B2(n221), 
	.B1(\ram[85][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n94));
   AO22CHD U3370 (.O(n1945), 
	.B2(n221), 
	.B1(\ram[85][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n94));
   AO22CHD U3371 (.O(n1946), 
	.B2(n221), 
	.B1(\ram[85][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n94));
   AO22CHD U3372 (.O(n1947), 
	.B2(n221), 
	.B1(\ram[85][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n94));
   AO22CHD U3373 (.O(n1948), 
	.B2(n221), 
	.B1(\ram[85][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n94));
   AO22CHD U3374 (.O(n1949), 
	.B2(n221), 
	.B1(\ram[85][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n94));
   AO22CHD U3375 (.O(n1950), 
	.B2(n221), 
	.B1(\ram[85][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n94));
   AO22CHD U3376 (.O(n1951), 
	.B2(n221), 
	.B1(\ram[85][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n94));
   AO22CHD U3377 (.O(n1952), 
	.B2(n221), 
	.B1(\ram[85][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n94));
   AO22CHD U3378 (.O(n1953), 
	.B2(n221), 
	.B1(\ram[85][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n94));
   AO22CHD U3379 (.O(n1954), 
	.B2(n221), 
	.B1(\ram[85][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n94));
   AO22CHD U3380 (.O(n1955), 
	.B2(n221), 
	.B1(\ram[85][13] ), 
	.A2(n21), 
	.A1(n94));
   AO22CHD U3381 (.O(n1956), 
	.B2(n221), 
	.B1(\ram[85][14] ), 
	.A2(n22), 
	.A1(n94));
   AO22CHD U3382 (.O(n1957), 
	.B2(n221), 
	.B1(\ram[85][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n94));
   AO22CHD U3383 (.O(n1958), 
	.B2(n223), 
	.B1(\ram[86][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n96));
   AO22CHD U3384 (.O(n1959), 
	.B2(n223), 
	.B1(\ram[86][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n96));
   AO22CHD U3385 (.O(n1960), 
	.B2(n223), 
	.B1(\ram[86][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n96));
   AO22CHD U3386 (.O(n1961), 
	.B2(n223), 
	.B1(\ram[86][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n96));
   AO22CHD U3387 (.O(n1962), 
	.B2(n223), 
	.B1(\ram[86][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n96));
   AO22CHD U3388 (.O(n1963), 
	.B2(n223), 
	.B1(\ram[86][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n96));
   AO22CHD U3389 (.O(n1964), 
	.B2(n223), 
	.B1(\ram[86][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n96));
   AO22CHD U3390 (.O(n1965), 
	.B2(n223), 
	.B1(\ram[86][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n96));
   AO22CHD U3391 (.O(n1966), 
	.B2(n223), 
	.B1(\ram[86][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n96));
   AO22CHD U3392 (.O(n1967), 
	.B2(n223), 
	.B1(\ram[86][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n96));
   AO22CHD U3393 (.O(n1968), 
	.B2(n223), 
	.B1(\ram[86][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n96));
   AO22CHD U3394 (.O(n1969), 
	.B2(n223), 
	.B1(\ram[86][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n96));
   AO22CHD U3395 (.O(n1970), 
	.B2(n223), 
	.B1(\ram[86][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n96));
   AO22CHD U3396 (.O(n1971), 
	.B2(n223), 
	.B1(\ram[86][13] ), 
	.A2(n21), 
	.A1(n96));
   AO22CHD U3397 (.O(n1972), 
	.B2(n223), 
	.B1(\ram[86][14] ), 
	.A2(n22), 
	.A1(n96));
   AO22CHD U3398 (.O(n1973), 
	.B2(n223), 
	.B1(\ram[86][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n96));
   AO22CHD U3399 (.O(n1974), 
	.B2(n225), 
	.B1(\ram[87][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n98));
   AO22CHD U3400 (.O(n1975), 
	.B2(n225), 
	.B1(\ram[87][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n98));
   AO22CHD U3401 (.O(n1976), 
	.B2(n225), 
	.B1(\ram[87][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n98));
   AO22CHD U3402 (.O(n1977), 
	.B2(n225), 
	.B1(\ram[87][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n98));
   AO22CHD U3403 (.O(n1978), 
	.B2(n225), 
	.B1(\ram[87][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n98));
   AO22CHD U3404 (.O(n1979), 
	.B2(n225), 
	.B1(\ram[87][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n98));
   AO22CHD U3405 (.O(n1980), 
	.B2(n225), 
	.B1(\ram[87][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n98));
   AO22CHD U3406 (.O(n1981), 
	.B2(n225), 
	.B1(\ram[87][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n98));
   AO22CHD U3407 (.O(n1982), 
	.B2(n225), 
	.B1(\ram[87][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n98));
   AO22CHD U3408 (.O(n1983), 
	.B2(n225), 
	.B1(\ram[87][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n98));
   AO22CHD U3409 (.O(n1984), 
	.B2(n225), 
	.B1(\ram[87][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n98));
   AO22CHD U3410 (.O(n1985), 
	.B2(n225), 
	.B1(\ram[87][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n98));
   AO22CHD U3411 (.O(n1986), 
	.B2(n225), 
	.B1(\ram[87][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n98));
   AO22CHD U3412 (.O(n1987), 
	.B2(n225), 
	.B1(\ram[87][13] ), 
	.A2(n21), 
	.A1(n98));
   AO22CHD U3413 (.O(n1988), 
	.B2(n225), 
	.B1(\ram[87][14] ), 
	.A2(n22), 
	.A1(n98));
   AO22CHD U3414 (.O(n1989), 
	.B2(n225), 
	.B1(\ram[87][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n98));
   AO22CHD U3415 (.O(n1990), 
	.B2(n227), 
	.B1(\ram[88][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n100));
   AO22CHD U3416 (.O(n1991), 
	.B2(n227), 
	.B1(\ram[88][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n100));
   AO22CHD U3417 (.O(n1992), 
	.B2(n227), 
	.B1(\ram[88][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n100));
   AO22CHD U3418 (.O(n1993), 
	.B2(n227), 
	.B1(\ram[88][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n100));
   AO22CHD U3419 (.O(n1994), 
	.B2(n227), 
	.B1(\ram[88][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n100));
   AO22CHD U3420 (.O(n1995), 
	.B2(n227), 
	.B1(\ram[88][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n100));
   AO22CHD U3421 (.O(n1996), 
	.B2(n227), 
	.B1(\ram[88][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n100));
   AO22CHD U3422 (.O(n1997), 
	.B2(n227), 
	.B1(\ram[88][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n100));
   AO22CHD U3423 (.O(n1998), 
	.B2(n227), 
	.B1(\ram[88][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n100));
   AO22CHD U3424 (.O(n1999), 
	.B2(n227), 
	.B1(\ram[88][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n100));
   AO22CHD U3425 (.O(n2000), 
	.B2(n227), 
	.B1(\ram[88][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n100));
   AO22CHD U3426 (.O(n2001), 
	.B2(n227), 
	.B1(\ram[88][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n100));
   AO22CHD U3427 (.O(n2002), 
	.B2(n227), 
	.B1(\ram[88][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n100));
   AO22CHD U3428 (.O(n2003), 
	.B2(n227), 
	.B1(\ram[88][13] ), 
	.A2(n21), 
	.A1(n100));
   AO22CHD U3429 (.O(n2004), 
	.B2(n227), 
	.B1(\ram[88][14] ), 
	.A2(n22), 
	.A1(n100));
   AO22CHD U3430 (.O(n2005), 
	.B2(n227), 
	.B1(\ram[88][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n100));
   AO22CHD U3431 (.O(n2006), 
	.B2(n229), 
	.B1(\ram[89][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n102));
   AO22CHD U3432 (.O(n2007), 
	.B2(n229), 
	.B1(\ram[89][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n102));
   AO22CHD U3433 (.O(n2008), 
	.B2(n229), 
	.B1(\ram[89][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n102));
   AO22CHD U3434 (.O(n2009), 
	.B2(n229), 
	.B1(\ram[89][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n102));
   AO22CHD U3435 (.O(n2010), 
	.B2(n229), 
	.B1(\ram[89][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n102));
   AO22CHD U3436 (.O(n2011), 
	.B2(n229), 
	.B1(\ram[89][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n102));
   AO22CHD U3437 (.O(n2012), 
	.B2(n229), 
	.B1(\ram[89][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n102));
   AO22CHD U3438 (.O(n2013), 
	.B2(n229), 
	.B1(\ram[89][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n102));
   AO22CHD U3439 (.O(n2014), 
	.B2(n229), 
	.B1(\ram[89][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n102));
   AO22CHD U3440 (.O(n2015), 
	.B2(n229), 
	.B1(\ram[89][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n102));
   AO22CHD U3441 (.O(n2016), 
	.B2(n229), 
	.B1(\ram[89][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n102));
   AO22CHD U3442 (.O(n2017), 
	.B2(n229), 
	.B1(\ram[89][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n102));
   AO22CHD U3443 (.O(n2018), 
	.B2(n229), 
	.B1(\ram[89][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n102));
   AO22CHD U3444 (.O(n2019), 
	.B2(n229), 
	.B1(\ram[89][13] ), 
	.A2(n21), 
	.A1(n102));
   AO22CHD U3445 (.O(n2020), 
	.B2(n229), 
	.B1(\ram[89][14] ), 
	.A2(n22), 
	.A1(n102));
   AO22CHD U3446 (.O(n2021), 
	.B2(n229), 
	.B1(\ram[89][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n102));
   AO22CHD U3447 (.O(n2022), 
	.B2(n231), 
	.B1(\ram[90][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n104));
   AO22CHD U3448 (.O(n2023), 
	.B2(n231), 
	.B1(\ram[90][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n104));
   AO22CHD U3449 (.O(n2024), 
	.B2(n231), 
	.B1(\ram[90][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n104));
   AO22CHD U3450 (.O(n2025), 
	.B2(n231), 
	.B1(\ram[90][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n104));
   AO22CHD U3451 (.O(n2026), 
	.B2(n231), 
	.B1(\ram[90][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n104));
   AO22CHD U3452 (.O(n2027), 
	.B2(n231), 
	.B1(\ram[90][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n104));
   AO22CHD U3453 (.O(n2028), 
	.B2(n231), 
	.B1(\ram[90][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n104));
   AO22CHD U3454 (.O(n2029), 
	.B2(n231), 
	.B1(\ram[90][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n104));
   AO22CHD U3455 (.O(n2030), 
	.B2(n231), 
	.B1(\ram[90][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n104));
   AO22CHD U3456 (.O(n2031), 
	.B2(n231), 
	.B1(\ram[90][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n104));
   AO22CHD U3457 (.O(n2032), 
	.B2(n231), 
	.B1(\ram[90][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n104));
   AO22CHD U3458 (.O(n2033), 
	.B2(n231), 
	.B1(\ram[90][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n104));
   AO22CHD U3459 (.O(n2034), 
	.B2(n231), 
	.B1(\ram[90][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n104));
   AO22CHD U3460 (.O(n2035), 
	.B2(n231), 
	.B1(\ram[90][13] ), 
	.A2(n21), 
	.A1(n104));
   AO22CHD U3461 (.O(n2036), 
	.B2(n231), 
	.B1(\ram[90][14] ), 
	.A2(n22), 
	.A1(n104));
   AO22CHD U3462 (.O(n2037), 
	.B2(n231), 
	.B1(\ram[90][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n104));
   AO22CHD U3463 (.O(n2038), 
	.B2(n233), 
	.B1(\ram[91][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n107));
   AO22CHD U3464 (.O(n2039), 
	.B2(n233), 
	.B1(\ram[91][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n107));
   AO22CHD U3465 (.O(n2040), 
	.B2(n233), 
	.B1(\ram[91][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n107));
   AO22CHD U3466 (.O(n2041), 
	.B2(n233), 
	.B1(\ram[91][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n107));
   AO22CHD U3467 (.O(n2042), 
	.B2(n233), 
	.B1(\ram[91][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n107));
   AO22CHD U3468 (.O(n2043), 
	.B2(n233), 
	.B1(\ram[91][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n107));
   AO22CHD U3469 (.O(n2044), 
	.B2(n233), 
	.B1(\ram[91][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n107));
   AO22CHD U3470 (.O(n2045), 
	.B2(n233), 
	.B1(\ram[91][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n107));
   AO22CHD U3471 (.O(n2046), 
	.B2(n233), 
	.B1(\ram[91][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n107));
   AO22CHD U3472 (.O(n2047), 
	.B2(n233), 
	.B1(\ram[91][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n107));
   AO22CHD U3473 (.O(n2048), 
	.B2(n233), 
	.B1(\ram[91][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n107));
   AO22CHD U3474 (.O(n2049), 
	.B2(n233), 
	.B1(\ram[91][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n107));
   AO22CHD U3475 (.O(n2050), 
	.B2(n233), 
	.B1(\ram[91][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n107));
   AO22CHD U3476 (.O(n2051), 
	.B2(n233), 
	.B1(\ram[91][13] ), 
	.A2(n21), 
	.A1(n107));
   AO22CHD U3477 (.O(n2052), 
	.B2(n233), 
	.B1(\ram[91][14] ), 
	.A2(n22), 
	.A1(n107));
   AO22CHD U3478 (.O(n2053), 
	.B2(n233), 
	.B1(\ram[91][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n107));
   AO22CHD U3479 (.O(n2054), 
	.B2(n235), 
	.B1(\ram[92][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n109));
   AO22CHD U3480 (.O(n2055), 
	.B2(n235), 
	.B1(\ram[92][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n109));
   AO22CHD U3481 (.O(n2056), 
	.B2(n235), 
	.B1(\ram[92][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n109));
   AO22CHD U3482 (.O(n2057), 
	.B2(n235), 
	.B1(\ram[92][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n109));
   AO22CHD U3483 (.O(n2058), 
	.B2(n235), 
	.B1(\ram[92][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n109));
   AO22CHD U3484 (.O(n2059), 
	.B2(n235), 
	.B1(\ram[92][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n109));
   AO22CHD U3485 (.O(n2060), 
	.B2(n235), 
	.B1(\ram[92][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n109));
   AO22CHD U3486 (.O(n2061), 
	.B2(n235), 
	.B1(\ram[92][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n109));
   AO22CHD U3487 (.O(n2062), 
	.B2(n235), 
	.B1(\ram[92][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n109));
   AO22CHD U3488 (.O(n2063), 
	.B2(n235), 
	.B1(\ram[92][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n109));
   AO22CHD U3489 (.O(n2064), 
	.B2(n235), 
	.B1(\ram[92][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n109));
   AO22CHD U3490 (.O(n2065), 
	.B2(n235), 
	.B1(\ram[92][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n109));
   AO22CHD U3491 (.O(n2066), 
	.B2(n235), 
	.B1(\ram[92][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n109));
   AO22CHD U3492 (.O(n2067), 
	.B2(n235), 
	.B1(\ram[92][13] ), 
	.A2(n21), 
	.A1(n109));
   AO22CHD U3493 (.O(n2068), 
	.B2(n235), 
	.B1(\ram[92][14] ), 
	.A2(n22), 
	.A1(n109));
   AO22CHD U3494 (.O(n2069), 
	.B2(n235), 
	.B1(\ram[92][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n109));
   AO22CHD U3495 (.O(n2070), 
	.B2(n237), 
	.B1(\ram[93][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n110));
   AO22CHD U3496 (.O(n2071), 
	.B2(n237), 
	.B1(\ram[93][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n110));
   AO22CHD U3497 (.O(n2072), 
	.B2(n237), 
	.B1(\ram[93][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n110));
   AO22CHD U3498 (.O(n2073), 
	.B2(n237), 
	.B1(\ram[93][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n110));
   AO22CHD U3499 (.O(n2074), 
	.B2(n237), 
	.B1(\ram[93][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n110));
   AO22CHD U3500 (.O(n2075), 
	.B2(n237), 
	.B1(\ram[93][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n110));
   AO22CHD U3501 (.O(n2076), 
	.B2(n237), 
	.B1(\ram[93][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n110));
   AO22CHD U3502 (.O(n2077), 
	.B2(n237), 
	.B1(\ram[93][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n110));
   AO22CHD U3503 (.O(n2078), 
	.B2(n237), 
	.B1(\ram[93][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n110));
   AO22CHD U3504 (.O(n2079), 
	.B2(n237), 
	.B1(\ram[93][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n110));
   AO22CHD U3505 (.O(n2080), 
	.B2(n237), 
	.B1(\ram[93][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n110));
   AO22CHD U3506 (.O(n2081), 
	.B2(n237), 
	.B1(\ram[93][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n110));
   AO22CHD U3507 (.O(n2082), 
	.B2(n237), 
	.B1(\ram[93][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n110));
   AO22CHD U3508 (.O(n2083), 
	.B2(n237), 
	.B1(\ram[93][13] ), 
	.A2(n21), 
	.A1(n110));
   AO22CHD U3509 (.O(n2084), 
	.B2(n237), 
	.B1(\ram[93][14] ), 
	.A2(n22), 
	.A1(n110));
   AO22CHD U3510 (.O(n2085), 
	.B2(n237), 
	.B1(\ram[93][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n110));
   AO22CHD U3511 (.O(n2086), 
	.B2(n239), 
	.B1(\ram[94][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n112));
   AO22CHD U3512 (.O(n2087), 
	.B2(n239), 
	.B1(\ram[94][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n112));
   AO22CHD U3513 (.O(n2088), 
	.B2(n239), 
	.B1(\ram[94][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n112));
   AO22CHD U3514 (.O(n2089), 
	.B2(n239), 
	.B1(\ram[94][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n112));
   AO22CHD U3515 (.O(n2090), 
	.B2(n239), 
	.B1(\ram[94][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n112));
   AO22CHD U3516 (.O(n2091), 
	.B2(n239), 
	.B1(\ram[94][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n112));
   AO22CHD U3517 (.O(n2092), 
	.B2(n239), 
	.B1(\ram[94][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n112));
   AO22CHD U3518 (.O(n2093), 
	.B2(n239), 
	.B1(\ram[94][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n112));
   AO22CHD U3519 (.O(n2094), 
	.B2(n239), 
	.B1(\ram[94][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n112));
   AO22CHD U3520 (.O(n2095), 
	.B2(n239), 
	.B1(\ram[94][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n112));
   AO22CHD U3521 (.O(n2096), 
	.B2(n239), 
	.B1(\ram[94][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n112));
   AO22CHD U3522 (.O(n2097), 
	.B2(n239), 
	.B1(\ram[94][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n112));
   AO22CHD U3523 (.O(n2098), 
	.B2(n239), 
	.B1(\ram[94][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n112));
   AO22CHD U3524 (.O(n2099), 
	.B2(n239), 
	.B1(\ram[94][13] ), 
	.A2(n21), 
	.A1(n112));
   AO22CHD U3525 (.O(n2100), 
	.B2(n239), 
	.B1(\ram[94][14] ), 
	.A2(n22), 
	.A1(n112));
   AO22CHD U3526 (.O(n2101), 
	.B2(n239), 
	.B1(\ram[94][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n112));
   AO22CHD U3527 (.O(n2102), 
	.B2(n241), 
	.B1(\ram[95][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n114));
   AO22CHD U3528 (.O(n2103), 
	.B2(n241), 
	.B1(\ram[95][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n114));
   AO22CHD U3529 (.O(n2104), 
	.B2(n241), 
	.B1(\ram[95][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n114));
   AO22CHD U3530 (.O(n2105), 
	.B2(n241), 
	.B1(\ram[95][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n114));
   AO22CHD U3531 (.O(n2106), 
	.B2(n241), 
	.B1(\ram[95][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n114));
   AO22CHD U3532 (.O(n2107), 
	.B2(n241), 
	.B1(\ram[95][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n114));
   AO22CHD U3533 (.O(n2108), 
	.B2(n241), 
	.B1(\ram[95][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n114));
   AO22CHD U3534 (.O(n2109), 
	.B2(n241), 
	.B1(\ram[95][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n114));
   AO22CHD U3535 (.O(n2110), 
	.B2(n241), 
	.B1(\ram[95][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n114));
   AO22CHD U3536 (.O(n2111), 
	.B2(n241), 
	.B1(\ram[95][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n114));
   AO22CHD U3537 (.O(n2112), 
	.B2(n241), 
	.B1(\ram[95][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n114));
   AO22CHD U3538 (.O(n2113), 
	.B2(n241), 
	.B1(\ram[95][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n114));
   AO22CHD U3539 (.O(n2114), 
	.B2(n241), 
	.B1(\ram[95][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n114));
   AO22CHD U3540 (.O(n2115), 
	.B2(n241), 
	.B1(\ram[95][13] ), 
	.A2(n21), 
	.A1(n114));
   AO22CHD U3541 (.O(n2116), 
	.B2(n241), 
	.B1(\ram[95][14] ), 
	.A2(n22), 
	.A1(n114));
   AO22CHD U3542 (.O(n2117), 
	.B2(n241), 
	.B1(\ram[95][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n114));
   AO22CHD U3543 (.O(n2118), 
	.B2(n243), 
	.B1(\ram[96][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n116));
   AO22CHD U3544 (.O(n2119), 
	.B2(n243), 
	.B1(\ram[96][1] ), 
	.A2(n9), 
	.A1(n116));
   AO22CHD U3545 (.O(n2120), 
	.B2(n243), 
	.B1(\ram[96][2] ), 
	.A2(n10), 
	.A1(n116));
   AO22CHD U3546 (.O(n2121), 
	.B2(n243), 
	.B1(\ram[96][3] ), 
	.A2(n11), 
	.A1(n116));
   AO22CHD U3547 (.O(n2122), 
	.B2(n243), 
	.B1(\ram[96][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n116));
   AO22CHD U3548 (.O(n2123), 
	.B2(n243), 
	.B1(\ram[96][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n116));
   AO22CHD U3549 (.O(n2124), 
	.B2(n243), 
	.B1(\ram[96][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n116));
   AO22CHD U3550 (.O(n2125), 
	.B2(n243), 
	.B1(\ram[96][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n116));
   AO22CHD U3551 (.O(n2126), 
	.B2(n243), 
	.B1(\ram[96][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n116));
   AO22CHD U3552 (.O(n2127), 
	.B2(n243), 
	.B1(\ram[96][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n116));
   AO22CHD U3553 (.O(n2128), 
	.B2(n243), 
	.B1(\ram[96][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n116));
   AO22CHD U3554 (.O(n2129), 
	.B2(n243), 
	.B1(\ram[96][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n116));
   AO22CHD U3555 (.O(n2130), 
	.B2(n243), 
	.B1(\ram[96][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n116));
   AO22CHD U3556 (.O(n2131), 
	.B2(n243), 
	.B1(\ram[96][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n116));
   AO22CHD U3557 (.O(n2132), 
	.B2(n243), 
	.B1(\ram[96][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n116));
   AO22CHD U3558 (.O(n2133), 
	.B2(n243), 
	.B1(\ram[96][15] ), 
	.A2(n23), 
	.A1(n116));
   AO22CHD U3559 (.O(n2134), 
	.B2(n246), 
	.B1(\ram[97][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n118));
   AO22CHD U3560 (.O(n2135), 
	.B2(n246), 
	.B1(\ram[97][1] ), 
	.A2(n9), 
	.A1(n118));
   AO22CHD U3561 (.O(n2136), 
	.B2(n246), 
	.B1(\ram[97][2] ), 
	.A2(n10), 
	.A1(n118));
   AO22CHD U3562 (.O(n2137), 
	.B2(n246), 
	.B1(\ram[97][3] ), 
	.A2(n11), 
	.A1(n118));
   AO22CHD U3563 (.O(n2138), 
	.B2(n246), 
	.B1(\ram[97][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n118));
   AO22CHD U3564 (.O(n2139), 
	.B2(n246), 
	.B1(\ram[97][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n118));
   AO22CHD U3565 (.O(n2140), 
	.B2(n246), 
	.B1(\ram[97][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n118));
   AO22CHD U3566 (.O(n2141), 
	.B2(n246), 
	.B1(\ram[97][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n118));
   AO22CHD U3567 (.O(n2142), 
	.B2(n246), 
	.B1(\ram[97][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n118));
   AO22CHD U3568 (.O(n2143), 
	.B2(n246), 
	.B1(\ram[97][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n118));
   AO22CHD U3569 (.O(n2144), 
	.B2(n246), 
	.B1(\ram[97][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n118));
   AO22CHD U3570 (.O(n2145), 
	.B2(n246), 
	.B1(\ram[97][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n118));
   AO22CHD U3571 (.O(n2146), 
	.B2(n246), 
	.B1(\ram[97][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n118));
   AO22CHD U3572 (.O(n2147), 
	.B2(n246), 
	.B1(\ram[97][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n118));
   AO22CHD U3573 (.O(n2148), 
	.B2(n246), 
	.B1(\ram[97][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n118));
   AO22CHD U3574 (.O(n2149), 
	.B2(n246), 
	.B1(\ram[97][15] ), 
	.A2(n23), 
	.A1(n118));
   AO22CHD U3575 (.O(n2150), 
	.B2(n248), 
	.B1(\ram[98][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n120));
   AO22CHD U3576 (.O(n2151), 
	.B2(n248), 
	.B1(\ram[98][1] ), 
	.A2(n9), 
	.A1(n120));
   AO22CHD U3577 (.O(n2152), 
	.B2(n248), 
	.B1(\ram[98][2] ), 
	.A2(n10), 
	.A1(n120));
   AO22CHD U3578 (.O(n2153), 
	.B2(n248), 
	.B1(\ram[98][3] ), 
	.A2(n11), 
	.A1(n120));
   AO22CHD U3579 (.O(n2154), 
	.B2(n248), 
	.B1(\ram[98][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n120));
   AO22CHD U3580 (.O(n2155), 
	.B2(n248), 
	.B1(\ram[98][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n120));
   AO22CHD U3581 (.O(n2156), 
	.B2(n248), 
	.B1(\ram[98][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n120));
   AO22CHD U3582 (.O(n2157), 
	.B2(n248), 
	.B1(\ram[98][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n120));
   AO22CHD U3583 (.O(n2158), 
	.B2(n248), 
	.B1(\ram[98][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n120));
   AO22CHD U3584 (.O(n2159), 
	.B2(n248), 
	.B1(\ram[98][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n120));
   AO22CHD U3585 (.O(n2160), 
	.B2(n248), 
	.B1(\ram[98][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n120));
   AO22CHD U3586 (.O(n2161), 
	.B2(n248), 
	.B1(\ram[98][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n120));
   AO22CHD U3587 (.O(n2162), 
	.B2(n248), 
	.B1(\ram[98][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n120));
   AO22CHD U3588 (.O(n2163), 
	.B2(n248), 
	.B1(\ram[98][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n120));
   AO22CHD U3589 (.O(n2164), 
	.B2(n248), 
	.B1(\ram[98][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n120));
   AO22CHD U3590 (.O(n2165), 
	.B2(n248), 
	.B1(\ram[98][15] ), 
	.A2(n23), 
	.A1(n120));
   AO22CHD U3591 (.O(n2166), 
	.B2(n250), 
	.B1(\ram[99][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n122));
   AO22CHD U3592 (.O(n2167), 
	.B2(n250), 
	.B1(\ram[99][1] ), 
	.A2(n9), 
	.A1(n122));
   AO22CHD U3593 (.O(n2168), 
	.B2(n250), 
	.B1(\ram[99][2] ), 
	.A2(n10), 
	.A1(n122));
   AO22CHD U3594 (.O(n2169), 
	.B2(n250), 
	.B1(\ram[99][3] ), 
	.A2(n11), 
	.A1(n122));
   AO22CHD U3595 (.O(n2170), 
	.B2(n250), 
	.B1(\ram[99][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n122));
   AO22CHD U3596 (.O(n2171), 
	.B2(n250), 
	.B1(\ram[99][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n122));
   AO22CHD U3597 (.O(n2172), 
	.B2(n250), 
	.B1(\ram[99][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n122));
   AO22CHD U3598 (.O(n2173), 
	.B2(n250), 
	.B1(\ram[99][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n122));
   AO22CHD U3599 (.O(n2174), 
	.B2(n250), 
	.B1(\ram[99][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n122));
   AO22CHD U3600 (.O(n2175), 
	.B2(n250), 
	.B1(\ram[99][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n122));
   AO22CHD U3601 (.O(n2176), 
	.B2(n250), 
	.B1(\ram[99][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n122));
   AO22CHD U3602 (.O(n2177), 
	.B2(n250), 
	.B1(\ram[99][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n122));
   AO22CHD U3603 (.O(n2178), 
	.B2(n250), 
	.B1(\ram[99][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n122));
   AO22CHD U3604 (.O(n2179), 
	.B2(n250), 
	.B1(\ram[99][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n122));
   AO22CHD U3605 (.O(n2180), 
	.B2(n250), 
	.B1(\ram[99][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n122));
   AO22CHD U3606 (.O(n2181), 
	.B2(n250), 
	.B1(\ram[99][15] ), 
	.A2(n23), 
	.A1(n122));
   AO22CHD U3607 (.O(n2182), 
	.B2(n252), 
	.B1(\ram[100][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n124));
   AO22CHD U3608 (.O(n2183), 
	.B2(n252), 
	.B1(\ram[100][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n124));
   AO22CHD U3609 (.O(n2184), 
	.B2(n252), 
	.B1(\ram[100][2] ), 
	.A2(n10), 
	.A1(n124));
   AO22CHD U3610 (.O(n2185), 
	.B2(n252), 
	.B1(\ram[100][3] ), 
	.A2(n11), 
	.A1(n124));
   AO22CHD U3611 (.O(n2186), 
	.B2(n252), 
	.B1(\ram[100][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n124));
   AO22CHD U3612 (.O(n2187), 
	.B2(n252), 
	.B1(\ram[100][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n124));
   AO22CHD U3613 (.O(n2188), 
	.B2(n252), 
	.B1(\ram[100][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n124));
   AO22CHD U3614 (.O(n2189), 
	.B2(n252), 
	.B1(\ram[100][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n124));
   AO22CHD U3615 (.O(n2190), 
	.B2(n252), 
	.B1(\ram[100][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n124));
   AO22CHD U3616 (.O(n2191), 
	.B2(n252), 
	.B1(\ram[100][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n124));
   AO22CHD U3617 (.O(n2192), 
	.B2(n252), 
	.B1(\ram[100][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n124));
   AO22CHD U3618 (.O(n2193), 
	.B2(n252), 
	.B1(\ram[100][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n124));
   AO22CHD U3619 (.O(n2194), 
	.B2(n252), 
	.B1(\ram[100][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n124));
   AO22CHD U3620 (.O(n2195), 
	.B2(n252), 
	.B1(\ram[100][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n124));
   AO22CHD U3621 (.O(n2196), 
	.B2(n252), 
	.B1(\ram[100][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n124));
   AO22CHD U3622 (.O(n2197), 
	.B2(n252), 
	.B1(\ram[100][15] ), 
	.A2(n23), 
	.A1(n124));
   AO22CHD U3623 (.O(n2198), 
	.B2(n254), 
	.B1(\ram[101][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n126));
   AO22CHD U3624 (.O(n2199), 
	.B2(n254), 
	.B1(\ram[101][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n126));
   AO22CHD U3625 (.O(n2200), 
	.B2(n254), 
	.B1(\ram[101][2] ), 
	.A2(n10), 
	.A1(n126));
   AO22CHD U3626 (.O(n2201), 
	.B2(n254), 
	.B1(\ram[101][3] ), 
	.A2(n11), 
	.A1(n126));
   AO22CHD U3627 (.O(n2202), 
	.B2(n254), 
	.B1(\ram[101][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n126));
   AO22CHD U3628 (.O(n2203), 
	.B2(n254), 
	.B1(\ram[101][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n126));
   AO22CHD U3629 (.O(n2204), 
	.B2(n254), 
	.B1(\ram[101][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n126));
   AO22CHD U3630 (.O(n2205), 
	.B2(n254), 
	.B1(\ram[101][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n126));
   AO22CHD U3631 (.O(n2206), 
	.B2(n254), 
	.B1(\ram[101][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n126));
   AO22CHD U3632 (.O(n2207), 
	.B2(n254), 
	.B1(\ram[101][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n126));
   AO22CHD U3633 (.O(n2208), 
	.B2(n254), 
	.B1(\ram[101][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n126));
   AO22CHD U3634 (.O(n2209), 
	.B2(n254), 
	.B1(\ram[101][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n126));
   AO22CHD U3635 (.O(n2210), 
	.B2(n254), 
	.B1(\ram[101][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n126));
   AO22CHD U3636 (.O(n2211), 
	.B2(n254), 
	.B1(\ram[101][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n126));
   AO22CHD U3637 (.O(n2212), 
	.B2(n254), 
	.B1(\ram[101][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n126));
   AO22CHD U3638 (.O(n2213), 
	.B2(n254), 
	.B1(\ram[101][15] ), 
	.A2(n23), 
	.A1(n126));
   AO22CHD U3639 (.O(n2214), 
	.B2(n256), 
	.B1(\ram[102][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n128));
   AO22CHD U3640 (.O(n2215), 
	.B2(n256), 
	.B1(\ram[102][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n128));
   AO22CHD U3641 (.O(n2216), 
	.B2(n256), 
	.B1(\ram[102][2] ), 
	.A2(n10), 
	.A1(n128));
   AO22CHD U3642 (.O(n2217), 
	.B2(n256), 
	.B1(\ram[102][3] ), 
	.A2(n11), 
	.A1(n128));
   AO22CHD U3643 (.O(n2218), 
	.B2(n256), 
	.B1(\ram[102][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n128));
   AO22CHD U3644 (.O(n2219), 
	.B2(n256), 
	.B1(\ram[102][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n128));
   AO22CHD U3645 (.O(n2220), 
	.B2(n256), 
	.B1(\ram[102][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n128));
   AO22CHD U3646 (.O(n2221), 
	.B2(n256), 
	.B1(\ram[102][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n128));
   AO22CHD U3647 (.O(n2222), 
	.B2(n256), 
	.B1(\ram[102][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n128));
   AO22CHD U3648 (.O(n2223), 
	.B2(n256), 
	.B1(\ram[102][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n128));
   AO22CHD U3649 (.O(n2224), 
	.B2(n256), 
	.B1(\ram[102][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n128));
   AO22CHD U3650 (.O(n2225), 
	.B2(n256), 
	.B1(\ram[102][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n128));
   AO22CHD U3651 (.O(n2226), 
	.B2(n256), 
	.B1(\ram[102][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n128));
   AO22CHD U3652 (.O(n2227), 
	.B2(n256), 
	.B1(\ram[102][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n128));
   AO22CHD U3653 (.O(n2228), 
	.B2(n256), 
	.B1(\ram[102][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n128));
   AO22CHD U3654 (.O(n2229), 
	.B2(n256), 
	.B1(\ram[102][15] ), 
	.A2(n23), 
	.A1(n128));
   AO22CHD U3655 (.O(n2230), 
	.B2(n258), 
	.B1(\ram[103][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n130));
   AO22CHD U3656 (.O(n2231), 
	.B2(n258), 
	.B1(\ram[103][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n130));
   AO22CHD U3657 (.O(n2232), 
	.B2(n258), 
	.B1(\ram[103][2] ), 
	.A2(n10), 
	.A1(n130));
   AO22CHD U3658 (.O(n2233), 
	.B2(n258), 
	.B1(\ram[103][3] ), 
	.A2(n11), 
	.A1(n130));
   AO22CHD U3659 (.O(n2234), 
	.B2(n258), 
	.B1(\ram[103][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n130));
   AO22CHD U3660 (.O(n2235), 
	.B2(n258), 
	.B1(\ram[103][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n130));
   AO22CHD U3661 (.O(n2236), 
	.B2(n258), 
	.B1(\ram[103][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n130));
   AO22CHD U3662 (.O(n2237), 
	.B2(n258), 
	.B1(\ram[103][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n130));
   AO22CHD U3663 (.O(n2238), 
	.B2(n258), 
	.B1(\ram[103][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n130));
   AO22CHD U3664 (.O(n2239), 
	.B2(n258), 
	.B1(\ram[103][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n130));
   AO22CHD U3665 (.O(n2240), 
	.B2(n258), 
	.B1(\ram[103][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n130));
   AO22CHD U3666 (.O(n2241), 
	.B2(n258), 
	.B1(\ram[103][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n130));
   AO22CHD U3667 (.O(n2242), 
	.B2(n258), 
	.B1(\ram[103][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n130));
   AO22CHD U3668 (.O(n2243), 
	.B2(n258), 
	.B1(\ram[103][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n130));
   AO22CHD U3669 (.O(n2244), 
	.B2(n258), 
	.B1(\ram[103][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n130));
   AO22CHD U3670 (.O(n2245), 
	.B2(n258), 
	.B1(\ram[103][15] ), 
	.A2(n23), 
	.A1(n130));
   AO22CHD U3671 (.O(n2246), 
	.B2(n260), 
	.B1(\ram[104][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n132));
   AO22CHD U3672 (.O(n2247), 
	.B2(n260), 
	.B1(\ram[104][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n132));
   AO22CHD U3673 (.O(n2248), 
	.B2(n260), 
	.B1(\ram[104][2] ), 
	.A2(n10), 
	.A1(n132));
   AO22CHD U3674 (.O(n2249), 
	.B2(n260), 
	.B1(\ram[104][3] ), 
	.A2(n11), 
	.A1(n132));
   AO22CHD U3675 (.O(n2250), 
	.B2(n260), 
	.B1(\ram[104][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n132));
   AO22CHD U3676 (.O(n2251), 
	.B2(n260), 
	.B1(\ram[104][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n132));
   AO22CHD U3677 (.O(n2252), 
	.B2(n260), 
	.B1(\ram[104][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n132));
   AO22CHD U3678 (.O(n2253), 
	.B2(n260), 
	.B1(\ram[104][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n132));
   AO22CHD U3679 (.O(n2254), 
	.B2(n260), 
	.B1(\ram[104][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n132));
   AO22CHD U3680 (.O(n2255), 
	.B2(n260), 
	.B1(\ram[104][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n132));
   AO22CHD U3681 (.O(n2256), 
	.B2(n260), 
	.B1(\ram[104][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n132));
   AO22CHD U3682 (.O(n2257), 
	.B2(n260), 
	.B1(\ram[104][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n132));
   AO22CHD U3683 (.O(n2258), 
	.B2(n260), 
	.B1(\ram[104][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n132));
   AO22CHD U3684 (.O(n2259), 
	.B2(n260), 
	.B1(\ram[104][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n132));
   AO22CHD U3685 (.O(n2260), 
	.B2(n260), 
	.B1(\ram[104][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n132));
   AO22CHD U3686 (.O(n2261), 
	.B2(n260), 
	.B1(\ram[104][15] ), 
	.A2(n23), 
	.A1(n132));
   AO22CHD U3687 (.O(n2262), 
	.B2(n262), 
	.B1(\ram[105][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n134));
   AO22CHD U3688 (.O(n2263), 
	.B2(n262), 
	.B1(\ram[105][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n134));
   AO22CHD U3689 (.O(n2264), 
	.B2(n262), 
	.B1(\ram[105][2] ), 
	.A2(n10), 
	.A1(n134));
   AO22CHD U3690 (.O(n2265), 
	.B2(n262), 
	.B1(\ram[105][3] ), 
	.A2(n11), 
	.A1(n134));
   AO22CHD U3691 (.O(n2266), 
	.B2(n262), 
	.B1(\ram[105][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n134));
   AO22CHD U3692 (.O(n2267), 
	.B2(n262), 
	.B1(\ram[105][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n134));
   AO22CHD U3693 (.O(n2268), 
	.B2(n262), 
	.B1(\ram[105][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n134));
   AO22CHD U3694 (.O(n2269), 
	.B2(n262), 
	.B1(\ram[105][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n134));
   AO22CHD U3695 (.O(n2270), 
	.B2(n262), 
	.B1(\ram[105][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n134));
   AO22CHD U3696 (.O(n2271), 
	.B2(n262), 
	.B1(\ram[105][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n134));
   AO22CHD U3697 (.O(n2272), 
	.B2(n262), 
	.B1(\ram[105][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n134));
   AO22CHD U3698 (.O(n2273), 
	.B2(n262), 
	.B1(\ram[105][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n134));
   AO22CHD U3699 (.O(n2274), 
	.B2(n262), 
	.B1(\ram[105][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n134));
   AO22CHD U3700 (.O(n2275), 
	.B2(n262), 
	.B1(\ram[105][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n134));
   AO22CHD U3701 (.O(n2276), 
	.B2(n262), 
	.B1(\ram[105][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n134));
   AO22CHD U3702 (.O(n2277), 
	.B2(n262), 
	.B1(\ram[105][15] ), 
	.A2(n23), 
	.A1(n134));
   AO22CHD U3703 (.O(n2278), 
	.B2(n264), 
	.B1(\ram[106][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n136));
   AO22CHD U3704 (.O(n2279), 
	.B2(n264), 
	.B1(\ram[106][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n136));
   AO22CHD U3705 (.O(n2280), 
	.B2(n264), 
	.B1(\ram[106][2] ), 
	.A2(n10), 
	.A1(n136));
   AO22CHD U3706 (.O(n2281), 
	.B2(n264), 
	.B1(\ram[106][3] ), 
	.A2(n11), 
	.A1(n136));
   AO22CHD U3707 (.O(n2282), 
	.B2(n264), 
	.B1(\ram[106][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n136));
   AO22CHD U3708 (.O(n2283), 
	.B2(n264), 
	.B1(\ram[106][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n136));
   AO22CHD U3709 (.O(n2284), 
	.B2(n264), 
	.B1(\ram[106][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n136));
   AO22CHD U3710 (.O(n2285), 
	.B2(n264), 
	.B1(\ram[106][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n136));
   AO22CHD U3711 (.O(n2286), 
	.B2(n264), 
	.B1(\ram[106][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n136));
   AO22CHD U3712 (.O(n2287), 
	.B2(n264), 
	.B1(\ram[106][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n136));
   AO22CHD U3713 (.O(n2288), 
	.B2(n264), 
	.B1(\ram[106][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n136));
   AO22CHD U3714 (.O(n2289), 
	.B2(n264), 
	.B1(\ram[106][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n136));
   AO22CHD U3715 (.O(n2290), 
	.B2(n264), 
	.B1(\ram[106][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n136));
   AO22CHD U3716 (.O(n2291), 
	.B2(n264), 
	.B1(\ram[106][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n136));
   AO22CHD U3717 (.O(n2292), 
	.B2(n264), 
	.B1(\ram[106][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n136));
   AO22CHD U3718 (.O(n2293), 
	.B2(n264), 
	.B1(\ram[106][15] ), 
	.A2(n23), 
	.A1(n136));
   AO22CHD U3719 (.O(n2294), 
	.B2(n266), 
	.B1(\ram[107][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n138));
   AO22CHD U3720 (.O(n2295), 
	.B2(n266), 
	.B1(\ram[107][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n138));
   AO22CHD U3721 (.O(n2296), 
	.B2(n266), 
	.B1(\ram[107][2] ), 
	.A2(n10), 
	.A1(n138));
   AO22CHD U3722 (.O(n2297), 
	.B2(n266), 
	.B1(\ram[107][3] ), 
	.A2(n11), 
	.A1(n138));
   AO22CHD U3723 (.O(n2298), 
	.B2(n266), 
	.B1(\ram[107][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n138));
   AO22CHD U3724 (.O(n2299), 
	.B2(n266), 
	.B1(\ram[107][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n138));
   AO22CHD U3725 (.O(n2300), 
	.B2(n266), 
	.B1(\ram[107][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n138));
   AO22CHD U3726 (.O(n2301), 
	.B2(n266), 
	.B1(\ram[107][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n138));
   AO22CHD U3727 (.O(n2302), 
	.B2(n266), 
	.B1(\ram[107][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n138));
   AO22CHD U3728 (.O(n2303), 
	.B2(n266), 
	.B1(\ram[107][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n138));
   AO22CHD U3729 (.O(n2304), 
	.B2(n266), 
	.B1(\ram[107][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n138));
   AO22CHD U3730 (.O(n2305), 
	.B2(n266), 
	.B1(\ram[107][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n138));
   AO22CHD U3731 (.O(n2306), 
	.B2(n266), 
	.B1(\ram[107][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n138));
   AO22CHD U3732 (.O(n2307), 
	.B2(n266), 
	.B1(\ram[107][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n138));
   AO22CHD U3733 (.O(n2308), 
	.B2(n266), 
	.B1(\ram[107][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n138));
   AO22CHD U3734 (.O(n2309), 
	.B2(n266), 
	.B1(\ram[107][15] ), 
	.A2(n23), 
	.A1(n138));
   AO22CHD U3735 (.O(n2310), 
	.B2(n268), 
	.B1(\ram[108][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n141));
   AO22CHD U3736 (.O(n2311), 
	.B2(n268), 
	.B1(\ram[108][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n141));
   AO22CHD U3737 (.O(n2312), 
	.B2(n268), 
	.B1(\ram[108][2] ), 
	.A2(n10), 
	.A1(n141));
   AO22CHD U3738 (.O(n2313), 
	.B2(n268), 
	.B1(\ram[108][3] ), 
	.A2(n11), 
	.A1(n141));
   AO22CHD U3739 (.O(n2314), 
	.B2(n268), 
	.B1(\ram[108][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n141));
   AO22CHD U3740 (.O(n2315), 
	.B2(n268), 
	.B1(\ram[108][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n141));
   AO22CHD U3741 (.O(n2316), 
	.B2(n268), 
	.B1(\ram[108][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n141));
   AO22CHD U3742 (.O(n2317), 
	.B2(n268), 
	.B1(\ram[108][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n141));
   AO22CHD U3743 (.O(n2318), 
	.B2(n268), 
	.B1(\ram[108][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n141));
   AO22CHD U3744 (.O(n2319), 
	.B2(n268), 
	.B1(\ram[108][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n141));
   AO22CHD U3745 (.O(n2320), 
	.B2(n268), 
	.B1(\ram[108][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n141));
   AO22CHD U3746 (.O(n2321), 
	.B2(n268), 
	.B1(\ram[108][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n141));
   AO22CHD U3747 (.O(n2322), 
	.B2(n268), 
	.B1(\ram[108][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n141));
   AO22CHD U3748 (.O(n2323), 
	.B2(n268), 
	.B1(\ram[108][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n141));
   AO22CHD U3749 (.O(n2324), 
	.B2(n268), 
	.B1(\ram[108][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n141));
   AO22CHD U3750 (.O(n2325), 
	.B2(n268), 
	.B1(\ram[108][15] ), 
	.A2(n23), 
	.A1(n141));
   AO22CHD U3751 (.O(n2326), 
	.B2(n270), 
	.B1(\ram[109][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n143));
   AO22CHD U3752 (.O(n2327), 
	.B2(n270), 
	.B1(\ram[109][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n143));
   AO22CHD U3753 (.O(n2328), 
	.B2(n270), 
	.B1(\ram[109][2] ), 
	.A2(n10), 
	.A1(n143));
   AO22CHD U3754 (.O(n2329), 
	.B2(n270), 
	.B1(\ram[109][3] ), 
	.A2(n11), 
	.A1(n143));
   AO22CHD U3755 (.O(n2330), 
	.B2(n270), 
	.B1(\ram[109][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n143));
   AO22CHD U3756 (.O(n2331), 
	.B2(n270), 
	.B1(\ram[109][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n143));
   AO22CHD U3757 (.O(n2332), 
	.B2(n270), 
	.B1(\ram[109][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n143));
   AO22CHD U3758 (.O(n2333), 
	.B2(n270), 
	.B1(\ram[109][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n143));
   AO22CHD U3759 (.O(n2334), 
	.B2(n270), 
	.B1(\ram[109][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n143));
   AO22CHD U3760 (.O(n2335), 
	.B2(n270), 
	.B1(\ram[109][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n143));
   AO22CHD U3761 (.O(n2336), 
	.B2(n270), 
	.B1(\ram[109][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n143));
   AO22CHD U3762 (.O(n2337), 
	.B2(n270), 
	.B1(\ram[109][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n143));
   AO22CHD U3763 (.O(n2338), 
	.B2(n270), 
	.B1(\ram[109][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n143));
   AO22CHD U3764 (.O(n2339), 
	.B2(n270), 
	.B1(\ram[109][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n143));
   AO22CHD U3765 (.O(n2340), 
	.B2(n270), 
	.B1(\ram[109][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n143));
   AO22CHD U3766 (.O(n2341), 
	.B2(n270), 
	.B1(\ram[109][15] ), 
	.A2(n23), 
	.A1(n143));
   AO22CHD U3767 (.O(n2342), 
	.B2(n272), 
	.B1(\ram[110][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n144));
   AO22CHD U3768 (.O(n2343), 
	.B2(n272), 
	.B1(\ram[110][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n144));
   AO22CHD U3769 (.O(n2344), 
	.B2(n272), 
	.B1(\ram[110][2] ), 
	.A2(n10), 
	.A1(n144));
   AO22CHD U3770 (.O(n2345), 
	.B2(n272), 
	.B1(\ram[110][3] ), 
	.A2(n11), 
	.A1(n144));
   AO22CHD U3771 (.O(n2346), 
	.B2(n272), 
	.B1(\ram[110][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n144));
   AO22CHD U3772 (.O(n2347), 
	.B2(n272), 
	.B1(\ram[110][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n144));
   AO22CHD U3773 (.O(n2348), 
	.B2(n272), 
	.B1(\ram[110][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n144));
   AO22CHD U3774 (.O(n2349), 
	.B2(n272), 
	.B1(\ram[110][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n144));
   AO22CHD U3775 (.O(n2350), 
	.B2(n272), 
	.B1(\ram[110][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n144));
   AO22CHD U3776 (.O(n2351), 
	.B2(n272), 
	.B1(\ram[110][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n144));
   AO22CHD U3777 (.O(n2352), 
	.B2(n272), 
	.B1(\ram[110][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n144));
   AO22CHD U3778 (.O(n2353), 
	.B2(n272), 
	.B1(\ram[110][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n144));
   AO22CHD U3779 (.O(n2354), 
	.B2(n272), 
	.B1(\ram[110][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n144));
   AO22CHD U3780 (.O(n2355), 
	.B2(n272), 
	.B1(\ram[110][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n144));
   AO22CHD U3781 (.O(n2356), 
	.B2(n272), 
	.B1(\ram[110][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n144));
   AO22CHD U3782 (.O(n2357), 
	.B2(n272), 
	.B1(\ram[110][15] ), 
	.A2(n23), 
	.A1(n144));
   AO22CHD U3783 (.O(n2358), 
	.B2(n274), 
	.B1(\ram[111][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n146));
   AO22CHD U3784 (.O(n2359), 
	.B2(n274), 
	.B1(\ram[111][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n146));
   AO22CHD U3785 (.O(n2360), 
	.B2(n274), 
	.B1(\ram[111][2] ), 
	.A2(n10), 
	.A1(n146));
   AO22CHD U3786 (.O(n2361), 
	.B2(n274), 
	.B1(\ram[111][3] ), 
	.A2(n11), 
	.A1(n146));
   AO22CHD U3787 (.O(n2362), 
	.B2(n274), 
	.B1(\ram[111][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n146));
   AO22CHD U3788 (.O(n2363), 
	.B2(n274), 
	.B1(\ram[111][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n146));
   AO22CHD U3789 (.O(n2364), 
	.B2(n274), 
	.B1(\ram[111][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n146));
   AO22CHD U3790 (.O(n2365), 
	.B2(n274), 
	.B1(\ram[111][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n146));
   AO22CHD U3791 (.O(n2366), 
	.B2(n274), 
	.B1(\ram[111][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n146));
   AO22CHD U3792 (.O(n2367), 
	.B2(n274), 
	.B1(\ram[111][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n146));
   AO22CHD U3793 (.O(n2368), 
	.B2(n274), 
	.B1(\ram[111][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n146));
   AO22CHD U3794 (.O(n2369), 
	.B2(n274), 
	.B1(\ram[111][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n146));
   AO22CHD U3795 (.O(n2370), 
	.B2(n274), 
	.B1(\ram[111][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n146));
   AO22CHD U3796 (.O(n2371), 
	.B2(n274), 
	.B1(\ram[111][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n146));
   AO22CHD U3797 (.O(n2372), 
	.B2(n274), 
	.B1(\ram[111][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n146));
   AO22CHD U3798 (.O(n2373), 
	.B2(n274), 
	.B1(\ram[111][15] ), 
	.A2(n23), 
	.A1(n146));
   AO22CHD U3799 (.O(n2374), 
	.B2(n276), 
	.B1(\ram[112][0] ), 
	.A2(n6), 
	.A1(n148));
   AO22CHD U3800 (.O(n2375), 
	.B2(n276), 
	.B1(\ram[112][1] ), 
	.A2(n9), 
	.A1(n148));
   AO22CHD U3801 (.O(n2376), 
	.B2(n276), 
	.B1(\ram[112][2] ), 
	.A2(n10), 
	.A1(n148));
   AO22CHD U3802 (.O(n2377), 
	.B2(n276), 
	.B1(\ram[112][3] ), 
	.A2(n11), 
	.A1(n148));
   AO22CHD U3803 (.O(n2378), 
	.B2(n276), 
	.B1(\ram[112][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n148));
   AO22CHD U3804 (.O(n2379), 
	.B2(n276), 
	.B1(\ram[112][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n148));
   AO22CHD U3805 (.O(n2380), 
	.B2(n276), 
	.B1(\ram[112][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n148));
   AO22CHD U3806 (.O(n2381), 
	.B2(n276), 
	.B1(\ram[112][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n148));
   AO22CHD U3807 (.O(n2382), 
	.B2(n276), 
	.B1(\ram[112][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n148));
   AO22CHD U3808 (.O(n2383), 
	.B2(n276), 
	.B1(\ram[112][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n148));
   AO22CHD U3809 (.O(n2384), 
	.B2(n276), 
	.B1(\ram[112][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n148));
   AO22CHD U3810 (.O(n2385), 
	.B2(n276), 
	.B1(\ram[112][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n148));
   AO22CHD U3811 (.O(n2386), 
	.B2(n276), 
	.B1(\ram[112][12] ), 
	.A2(n20), 
	.A1(n148));
   AO22CHD U3812 (.O(n2387), 
	.B2(n276), 
	.B1(\ram[112][13] ), 
	.A2(n21), 
	.A1(n148));
   AO22CHD U3813 (.O(n2388), 
	.B2(n276), 
	.B1(\ram[112][14] ), 
	.A2(n22), 
	.A1(n148));
   AO22CHD U3814 (.O(n2389), 
	.B2(n276), 
	.B1(\ram[112][15] ), 
	.A2(n23), 
	.A1(n148));
   AO22CHD U3815 (.O(n2390), 
	.B2(n279), 
	.B1(\ram[113][0] ), 
	.A2(n6), 
	.A1(n150));
   AO22CHD U3816 (.O(n2391), 
	.B2(n279), 
	.B1(\ram[113][1] ), 
	.A2(n9), 
	.A1(n150));
   AO22CHD U3817 (.O(n2392), 
	.B2(n279), 
	.B1(\ram[113][2] ), 
	.A2(n10), 
	.A1(n150));
   AO22CHD U3818 (.O(n2393), 
	.B2(n279), 
	.B1(\ram[113][3] ), 
	.A2(n11), 
	.A1(n150));
   AO22CHD U3819 (.O(n2394), 
	.B2(n279), 
	.B1(\ram[113][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n150));
   AO22CHD U3820 (.O(n2395), 
	.B2(n279), 
	.B1(\ram[113][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n150));
   AO22CHD U3821 (.O(n2396), 
	.B2(n279), 
	.B1(\ram[113][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n150));
   AO22CHD U3822 (.O(n2397), 
	.B2(n279), 
	.B1(\ram[113][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n150));
   AO22CHD U3823 (.O(n2398), 
	.B2(n279), 
	.B1(\ram[113][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n150));
   AO22CHD U3824 (.O(n2399), 
	.B2(n279), 
	.B1(\ram[113][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n150));
   AO22CHD U3825 (.O(n2400), 
	.B2(n279), 
	.B1(\ram[113][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n150));
   AO22CHD U3826 (.O(n2401), 
	.B2(n279), 
	.B1(\ram[113][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n150));
   AO22CHD U3827 (.O(n2402), 
	.B2(n279), 
	.B1(\ram[113][12] ), 
	.A2(n20), 
	.A1(n150));
   AO22CHD U3828 (.O(n2403), 
	.B2(n279), 
	.B1(\ram[113][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n150));
   AO22CHD U3829 (.O(n2404), 
	.B2(n279), 
	.B1(\ram[113][14] ), 
	.A2(n22), 
	.A1(n150));
   AO22CHD U3830 (.O(n2405), 
	.B2(n279), 
	.B1(\ram[113][15] ), 
	.A2(n23), 
	.A1(n150));
   AO22CHD U3831 (.O(n2406), 
	.B2(n281), 
	.B1(\ram[114][0] ), 
	.A2(n6), 
	.A1(n152));
   AO22CHD U3832 (.O(n2407), 
	.B2(n281), 
	.B1(\ram[114][1] ), 
	.A2(n9), 
	.A1(n152));
   AO22CHD U3833 (.O(n2408), 
	.B2(n281), 
	.B1(\ram[114][2] ), 
	.A2(n10), 
	.A1(n152));
   AO22CHD U3834 (.O(n2409), 
	.B2(n281), 
	.B1(\ram[114][3] ), 
	.A2(n11), 
	.A1(n152));
   AO22CHD U3835 (.O(n2410), 
	.B2(n281), 
	.B1(\ram[114][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n152));
   AO22CHD U3836 (.O(n2411), 
	.B2(n281), 
	.B1(\ram[114][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n152));
   AO22CHD U3837 (.O(n2412), 
	.B2(n281), 
	.B1(\ram[114][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n152));
   AO22CHD U3838 (.O(n2413), 
	.B2(n281), 
	.B1(\ram[114][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n152));
   AO22CHD U3839 (.O(n2414), 
	.B2(n281), 
	.B1(\ram[114][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n152));
   AO22CHD U3840 (.O(n2415), 
	.B2(n281), 
	.B1(\ram[114][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n152));
   AO22CHD U3841 (.O(n2416), 
	.B2(n281), 
	.B1(\ram[114][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n152));
   AO22CHD U3842 (.O(n2417), 
	.B2(n281), 
	.B1(\ram[114][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n152));
   AO22CHD U3843 (.O(n2418), 
	.B2(n281), 
	.B1(\ram[114][12] ), 
	.A2(n20), 
	.A1(n152));
   AO22CHD U3844 (.O(n2419), 
	.B2(n281), 
	.B1(\ram[114][13] ), 
	.A2(n21), 
	.A1(n152));
   AO22CHD U3845 (.O(n2420), 
	.B2(n281), 
	.B1(\ram[114][14] ), 
	.A2(n22), 
	.A1(n152));
   AO22CHD U3846 (.O(n2421), 
	.B2(n281), 
	.B1(\ram[114][15] ), 
	.A2(n23), 
	.A1(n152));
   AO22CHD U3847 (.O(n2422), 
	.B2(n283), 
	.B1(\ram[115][0] ), 
	.A2(n6), 
	.A1(n154));
   AO22CHD U3848 (.O(n2423), 
	.B2(n283), 
	.B1(\ram[115][1] ), 
	.A2(n9), 
	.A1(n154));
   AO22CHD U3849 (.O(n2424), 
	.B2(n283), 
	.B1(\ram[115][2] ), 
	.A2(n10), 
	.A1(n154));
   AO22CHD U3850 (.O(n2425), 
	.B2(n283), 
	.B1(\ram[115][3] ), 
	.A2(n11), 
	.A1(n154));
   AO22CHD U3851 (.O(n2426), 
	.B2(n283), 
	.B1(\ram[115][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n154));
   AO22CHD U3852 (.O(n2427), 
	.B2(n283), 
	.B1(\ram[115][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n154));
   AO22CHD U3853 (.O(n2428), 
	.B2(n283), 
	.B1(\ram[115][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n154));
   AO22CHD U3854 (.O(n2429), 
	.B2(n283), 
	.B1(\ram[115][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n154));
   AO22CHD U3855 (.O(n2430), 
	.B2(n283), 
	.B1(\ram[115][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n154));
   AO22CHD U3856 (.O(n2431), 
	.B2(n283), 
	.B1(\ram[115][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n154));
   AO22CHD U3857 (.O(n2432), 
	.B2(n283), 
	.B1(\ram[115][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n154));
   AO22CHD U3858 (.O(n2433), 
	.B2(n283), 
	.B1(\ram[115][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n154));
   AO22CHD U3859 (.O(n2434), 
	.B2(n283), 
	.B1(\ram[115][12] ), 
	.A2(n20), 
	.A1(n154));
   AO22CHD U3860 (.O(n2435), 
	.B2(n283), 
	.B1(\ram[115][13] ), 
	.A2(n21), 
	.A1(n154));
   AO22CHD U3861 (.O(n2436), 
	.B2(n283), 
	.B1(\ram[115][14] ), 
	.A2(n22), 
	.A1(n154));
   AO22CHD U3862 (.O(n2437), 
	.B2(n283), 
	.B1(\ram[115][15] ), 
	.A2(n23), 
	.A1(n154));
   AO22CHD U3863 (.O(n2438), 
	.B2(n285), 
	.B1(\ram[116][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n156));
   AO22CHD U3864 (.O(n2439), 
	.B2(n285), 
	.B1(\ram[116][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n156));
   AO22CHD U3865 (.O(n2440), 
	.B2(n285), 
	.B1(\ram[116][2] ), 
	.A2(n10), 
	.A1(n156));
   AO22CHD U3866 (.O(n2441), 
	.B2(n285), 
	.B1(\ram[116][3] ), 
	.A2(n11), 
	.A1(n156));
   AO22CHD U3867 (.O(n2442), 
	.B2(n285), 
	.B1(\ram[116][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n156));
   AO22CHD U3868 (.O(n2443), 
	.B2(n285), 
	.B1(\ram[116][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n156));
   AO22CHD U3869 (.O(n2444), 
	.B2(n285), 
	.B1(\ram[116][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n156));
   AO22CHD U3870 (.O(n2445), 
	.B2(n285), 
	.B1(\ram[116][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n156));
   AO22CHD U3871 (.O(n2446), 
	.B2(n285), 
	.B1(\ram[116][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n156));
   AO22CHD U3872 (.O(n2447), 
	.B2(n285), 
	.B1(\ram[116][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n156));
   AO22CHD U3873 (.O(n2448), 
	.B2(n285), 
	.B1(\ram[116][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n156));
   AO22CHD U3874 (.O(n2449), 
	.B2(n285), 
	.B1(\ram[116][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n156));
   AO22CHD U3875 (.O(n2450), 
	.B2(n285), 
	.B1(\ram[116][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n156));
   AO22CHD U3876 (.O(n2451), 
	.B2(n285), 
	.B1(\ram[116][13] ), 
	.A2(n21), 
	.A1(n156));
   AO22CHD U3877 (.O(n2452), 
	.B2(n285), 
	.B1(\ram[116][14] ), 
	.A2(n22), 
	.A1(n156));
   AO22CHD U3878 (.O(n2453), 
	.B2(n285), 
	.B1(\ram[116][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n156));
   AO22CHD U3879 (.O(n2454), 
	.B2(n287), 
	.B1(\ram[117][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n158));
   AO22CHD U3880 (.O(n2455), 
	.B2(n287), 
	.B1(\ram[117][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n158));
   AO22CHD U3881 (.O(n2456), 
	.B2(n287), 
	.B1(\ram[117][2] ), 
	.A2(n10), 
	.A1(n158));
   AO22CHD U3882 (.O(n2457), 
	.B2(n287), 
	.B1(\ram[117][3] ), 
	.A2(n11), 
	.A1(n158));
   AO22CHD U3883 (.O(n2458), 
	.B2(n287), 
	.B1(\ram[117][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n158));
   AO22CHD U3884 (.O(n2459), 
	.B2(n287), 
	.B1(\ram[117][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n158));
   AO22CHD U3885 (.O(n2460), 
	.B2(n287), 
	.B1(\ram[117][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n158));
   AO22CHD U3886 (.O(n2461), 
	.B2(n287), 
	.B1(\ram[117][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n158));
   AO22CHD U3887 (.O(n2462), 
	.B2(n287), 
	.B1(\ram[117][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n158));
   AO22CHD U3888 (.O(n2463), 
	.B2(n287), 
	.B1(\ram[117][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n158));
   AO22CHD U3889 (.O(n2464), 
	.B2(n287), 
	.B1(\ram[117][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n158));
   AO22CHD U3890 (.O(n2465), 
	.B2(n287), 
	.B1(\ram[117][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n158));
   AO22CHD U3891 (.O(n2466), 
	.B2(n287), 
	.B1(\ram[117][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n158));
   AO22CHD U3892 (.O(n2467), 
	.B2(n287), 
	.B1(\ram[117][13] ), 
	.A2(n21), 
	.A1(n158));
   AO22CHD U3893 (.O(n2468), 
	.B2(n287), 
	.B1(\ram[117][14] ), 
	.A2(n22), 
	.A1(n158));
   AO22CHD U3894 (.O(n2469), 
	.B2(n287), 
	.B1(\ram[117][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n158));
   AO22CHD U3895 (.O(n2470), 
	.B2(n289), 
	.B1(\ram[118][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n160));
   AO22CHD U3896 (.O(n2471), 
	.B2(n289), 
	.B1(\ram[118][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n160));
   AO22CHD U3897 (.O(n2472), 
	.B2(n289), 
	.B1(\ram[118][2] ), 
	.A2(n10), 
	.A1(n160));
   AO22CHD U3898 (.O(n2473), 
	.B2(n289), 
	.B1(\ram[118][3] ), 
	.A2(n11), 
	.A1(n160));
   AO22CHD U3899 (.O(n2474), 
	.B2(n289), 
	.B1(\ram[118][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n160));
   AO22CHD U3900 (.O(n2475), 
	.B2(n289), 
	.B1(\ram[118][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n160));
   AO22CHD U3901 (.O(n2476), 
	.B2(n289), 
	.B1(\ram[118][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n160));
   AO22CHD U3902 (.O(n2477), 
	.B2(n289), 
	.B1(\ram[118][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n160));
   AO22CHD U3903 (.O(n2478), 
	.B2(n289), 
	.B1(\ram[118][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n160));
   AO22CHD U3904 (.O(n2479), 
	.B2(n289), 
	.B1(\ram[118][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n160));
   AO22CHD U3905 (.O(n2480), 
	.B2(n289), 
	.B1(\ram[118][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n160));
   AO22CHD U3906 (.O(n2481), 
	.B2(n289), 
	.B1(\ram[118][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n160));
   AO22CHD U3907 (.O(n2482), 
	.B2(n289), 
	.B1(\ram[118][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n160));
   AO22CHD U3908 (.O(n2483), 
	.B2(n289), 
	.B1(\ram[118][13] ), 
	.A2(n21), 
	.A1(n160));
   AO22CHD U3909 (.O(n2484), 
	.B2(n289), 
	.B1(\ram[118][14] ), 
	.A2(n22), 
	.A1(n160));
   AO22CHD U3910 (.O(n2485), 
	.B2(n289), 
	.B1(\ram[118][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n160));
   AO22CHD U3911 (.O(n2486), 
	.B2(n291), 
	.B1(\ram[119][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n162));
   AO22CHD U3912 (.O(n2487), 
	.B2(n291), 
	.B1(\ram[119][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n162));
   AO22CHD U3913 (.O(n2488), 
	.B2(n291), 
	.B1(\ram[119][2] ), 
	.A2(n10), 
	.A1(n162));
   AO22CHD U3914 (.O(n2489), 
	.B2(n291), 
	.B1(\ram[119][3] ), 
	.A2(n11), 
	.A1(n162));
   AO22CHD U3915 (.O(n2490), 
	.B2(n291), 
	.B1(\ram[119][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n162));
   AO22CHD U3916 (.O(n2491), 
	.B2(n291), 
	.B1(\ram[119][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n162));
   AO22CHD U3917 (.O(n2492), 
	.B2(n291), 
	.B1(\ram[119][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n162));
   AO22CHD U3918 (.O(n2493), 
	.B2(n291), 
	.B1(\ram[119][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n162));
   AO22CHD U3919 (.O(n2494), 
	.B2(n291), 
	.B1(\ram[119][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n162));
   AO22CHD U3920 (.O(n2495), 
	.B2(n291), 
	.B1(\ram[119][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n162));
   AO22CHD U3921 (.O(n2496), 
	.B2(n291), 
	.B1(\ram[119][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n162));
   AO22CHD U3922 (.O(n2497), 
	.B2(n291), 
	.B1(\ram[119][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n162));
   AO22CHD U3923 (.O(n2498), 
	.B2(n291), 
	.B1(\ram[119][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n162));
   AO22CHD U3924 (.O(n2499), 
	.B2(n291), 
	.B1(\ram[119][13] ), 
	.A2(n21), 
	.A1(n162));
   AO22CHD U3925 (.O(n2500), 
	.B2(n291), 
	.B1(\ram[119][14] ), 
	.A2(n22), 
	.A1(n162));
   AO22CHD U3926 (.O(n2501), 
	.B2(n291), 
	.B1(\ram[119][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n162));
   AO22CHD U3927 (.O(n2502), 
	.B2(n293), 
	.B1(\ram[120][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n164));
   AO22CHD U3928 (.O(n2503), 
	.B2(n293), 
	.B1(\ram[120][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n164));
   AO22CHD U3929 (.O(n2504), 
	.B2(n293), 
	.B1(\ram[120][2] ), 
	.A2(n10), 
	.A1(n164));
   AO22CHD U3930 (.O(n2505), 
	.B2(n293), 
	.B1(\ram[120][3] ), 
	.A2(n11), 
	.A1(n164));
   AO22CHD U3931 (.O(n2506), 
	.B2(n293), 
	.B1(\ram[120][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n164));
   AO22CHD U3932 (.O(n2507), 
	.B2(n293), 
	.B1(\ram[120][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n164));
   AO22CHD U3933 (.O(n2508), 
	.B2(n293), 
	.B1(\ram[120][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n164));
   AO22CHD U3934 (.O(n2509), 
	.B2(n293), 
	.B1(\ram[120][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n164));
   AO22CHD U3935 (.O(n2510), 
	.B2(n293), 
	.B1(\ram[120][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n164));
   AO22CHD U3936 (.O(n2511), 
	.B2(n293), 
	.B1(\ram[120][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n164));
   AO22CHD U3937 (.O(n2512), 
	.B2(n293), 
	.B1(\ram[120][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n164));
   AO22CHD U3938 (.O(n2513), 
	.B2(n293), 
	.B1(\ram[120][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n164));
   AO22CHD U3939 (.O(n2514), 
	.B2(n293), 
	.B1(\ram[120][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n164));
   AO22CHD U3940 (.O(n2515), 
	.B2(n293), 
	.B1(\ram[120][13] ), 
	.A2(n21), 
	.A1(n164));
   AO22CHD U3941 (.O(n2516), 
	.B2(n293), 
	.B1(\ram[120][14] ), 
	.A2(n22), 
	.A1(n164));
   AO22CHD U3942 (.O(n2517), 
	.B2(n293), 
	.B1(\ram[120][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n164));
   AO22CHD U3943 (.O(n2518), 
	.B2(n295), 
	.B1(\ram[121][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n166));
   AO22CHD U3944 (.O(n2519), 
	.B2(n295), 
	.B1(\ram[121][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n166));
   AO22CHD U3945 (.O(n2520), 
	.B2(n295), 
	.B1(\ram[121][2] ), 
	.A2(n10), 
	.A1(n166));
   AO22CHD U3946 (.O(n2521), 
	.B2(n295), 
	.B1(\ram[121][3] ), 
	.A2(n11), 
	.A1(n166));
   AO22CHD U3947 (.O(n2522), 
	.B2(n295), 
	.B1(\ram[121][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n166));
   AO22CHD U3948 (.O(n2523), 
	.B2(n295), 
	.B1(\ram[121][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n166));
   AO22CHD U3949 (.O(n2524), 
	.B2(n295), 
	.B1(\ram[121][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n166));
   AO22CHD U3950 (.O(n2525), 
	.B2(n295), 
	.B1(\ram[121][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n166));
   AO22CHD U3951 (.O(n2526), 
	.B2(n295), 
	.B1(\ram[121][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n166));
   AO22CHD U3952 (.O(n2527), 
	.B2(n295), 
	.B1(\ram[121][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n166));
   AO22CHD U3953 (.O(n2528), 
	.B2(n295), 
	.B1(\ram[121][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n166));
   AO22CHD U3954 (.O(n2529), 
	.B2(n295), 
	.B1(\ram[121][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n166));
   AO22CHD U3955 (.O(n2530), 
	.B2(n295), 
	.B1(\ram[121][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n166));
   AO22CHD U3956 (.O(n2531), 
	.B2(n295), 
	.B1(\ram[121][13] ), 
	.A2(n21), 
	.A1(n166));
   AO22CHD U3957 (.O(n2532), 
	.B2(n295), 
	.B1(\ram[121][14] ), 
	.A2(n22), 
	.A1(n166));
   AO22CHD U3958 (.O(n2533), 
	.B2(n295), 
	.B1(\ram[121][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n166));
   AO22CHD U3959 (.O(n2534), 
	.B2(n297), 
	.B1(\ram[122][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n168));
   AO22CHD U3960 (.O(n2535), 
	.B2(n297), 
	.B1(\ram[122][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n168));
   AO22CHD U3961 (.O(n2536), 
	.B2(n297), 
	.B1(\ram[122][2] ), 
	.A2(n10), 
	.A1(n168));
   AO22CHD U3962 (.O(n2537), 
	.B2(n297), 
	.B1(\ram[122][3] ), 
	.A2(n11), 
	.A1(n168));
   AO22CHD U3963 (.O(n2538), 
	.B2(n297), 
	.B1(\ram[122][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n168));
   AO22CHD U3964 (.O(n2539), 
	.B2(n297), 
	.B1(\ram[122][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n168));
   AO22CHD U3965 (.O(n2540), 
	.B2(n297), 
	.B1(\ram[122][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n168));
   AO22CHD U3966 (.O(n2541), 
	.B2(n297), 
	.B1(\ram[122][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n168));
   AO22CHD U3967 (.O(n2542), 
	.B2(n297), 
	.B1(\ram[122][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n168));
   AO22CHD U3968 (.O(n2543), 
	.B2(n297), 
	.B1(\ram[122][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n168));
   AO22CHD U3969 (.O(n2544), 
	.B2(n297), 
	.B1(\ram[122][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n168));
   AO22CHD U3970 (.O(n2545), 
	.B2(n297), 
	.B1(\ram[122][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n168));
   AO22CHD U3971 (.O(n2546), 
	.B2(n297), 
	.B1(\ram[122][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n168));
   AO22CHD U3972 (.O(n2547), 
	.B2(n297), 
	.B1(\ram[122][13] ), 
	.A2(n21), 
	.A1(n168));
   AO22CHD U3973 (.O(n2548), 
	.B2(n297), 
	.B1(\ram[122][14] ), 
	.A2(n22), 
	.A1(n168));
   AO22CHD U3974 (.O(n2549), 
	.B2(n297), 
	.B1(\ram[122][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n168));
   AO22CHD U3975 (.O(n2550), 
	.B2(n299), 
	.B1(\ram[123][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n170));
   AO22CHD U3976 (.O(n2551), 
	.B2(n299), 
	.B1(\ram[123][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n170));
   AO22CHD U3977 (.O(n2552), 
	.B2(n299), 
	.B1(\ram[123][2] ), 
	.A2(n10), 
	.A1(n170));
   AO22CHD U3978 (.O(n2553), 
	.B2(n299), 
	.B1(\ram[123][3] ), 
	.A2(n11), 
	.A1(n170));
   AO22CHD U3979 (.O(n2554), 
	.B2(n299), 
	.B1(\ram[123][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n170));
   AO22CHD U3980 (.O(n2555), 
	.B2(n299), 
	.B1(\ram[123][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n170));
   AO22CHD U3981 (.O(n2556), 
	.B2(n299), 
	.B1(\ram[123][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n170));
   AO22CHD U3982 (.O(n2557), 
	.B2(n299), 
	.B1(\ram[123][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n170));
   AO22CHD U3983 (.O(n2558), 
	.B2(n299), 
	.B1(\ram[123][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n170));
   AO22CHD U3984 (.O(n2559), 
	.B2(n299), 
	.B1(\ram[123][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n170));
   AO22CHD U3985 (.O(n2560), 
	.B2(n299), 
	.B1(\ram[123][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n170));
   AO22CHD U3986 (.O(n2561), 
	.B2(n299), 
	.B1(\ram[123][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n170));
   AO22CHD U3987 (.O(n2562), 
	.B2(n299), 
	.B1(\ram[123][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n170));
   AO22CHD U3988 (.O(n2563), 
	.B2(n299), 
	.B1(\ram[123][13] ), 
	.A2(n21), 
	.A1(n170));
   AO22CHD U3989 (.O(n2564), 
	.B2(n299), 
	.B1(\ram[123][14] ), 
	.A2(n22), 
	.A1(n170));
   AO22CHD U3990 (.O(n2565), 
	.B2(n299), 
	.B1(\ram[123][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n170));
   AO22CHD U3991 (.O(n2566), 
	.B2(n301), 
	.B1(\ram[124][0] ), 
	.A2(n6), 
	.A1(n172));
   AO22CHD U3992 (.O(n2567), 
	.B2(n301), 
	.B1(\ram[124][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n172));
   AO22CHD U3993 (.O(n2568), 
	.B2(n301), 
	.B1(\ram[124][2] ), 
	.A2(n10), 
	.A1(n172));
   AO22CHD U3994 (.O(n2569), 
	.B2(n301), 
	.B1(\ram[124][3] ), 
	.A2(n11), 
	.A1(n172));
   AO22CHD U3995 (.O(n2570), 
	.B2(n301), 
	.B1(\ram[124][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n172));
   AO22CHD U3996 (.O(n2571), 
	.B2(n301), 
	.B1(\ram[124][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n172));
   AO22CHD U3997 (.O(n2572), 
	.B2(n301), 
	.B1(\ram[124][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n172));
   AO22CHD U3998 (.O(n2573), 
	.B2(n301), 
	.B1(\ram[124][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n172));
   AO22CHD U3999 (.O(n2574), 
	.B2(n301), 
	.B1(\ram[124][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n172));
   AO22CHD U4000 (.O(n2575), 
	.B2(n301), 
	.B1(\ram[124][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n172));
   AO22CHD U4001 (.O(n2576), 
	.B2(n301), 
	.B1(\ram[124][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n172));
   AO22CHD U4002 (.O(n2577), 
	.B2(n301), 
	.B1(\ram[124][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n172));
   AO22CHD U4003 (.O(n2578), 
	.B2(n301), 
	.B1(\ram[124][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n172));
   AO22CHD U4004 (.O(n2579), 
	.B2(n301), 
	.B1(\ram[124][13] ), 
	.A2(n21), 
	.A1(n172));
   AO22CHD U4005 (.O(n2580), 
	.B2(n301), 
	.B1(\ram[124][14] ), 
	.A2(n22), 
	.A1(n172));
   AO22CHD U4006 (.O(n2581), 
	.B2(n301), 
	.B1(\ram[124][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n172));
   AO22CHD U4007 (.O(n2582), 
	.B2(n303), 
	.B1(\ram[125][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n175));
   AO22CHD U4008 (.O(n2583), 
	.B2(n303), 
	.B1(\ram[125][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n175));
   AO22CHD U4009 (.O(n2584), 
	.B2(n303), 
	.B1(\ram[125][2] ), 
	.A2(n10), 
	.A1(n175));
   AO22CHD U4010 (.O(n2585), 
	.B2(n303), 
	.B1(\ram[125][3] ), 
	.A2(n11), 
	.A1(n175));
   AO22CHD U4011 (.O(n2586), 
	.B2(n303), 
	.B1(\ram[125][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n175));
   AO22CHD U4012 (.O(n2587), 
	.B2(n303), 
	.B1(\ram[125][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n175));
   AO22CHD U4013 (.O(n2588), 
	.B2(n303), 
	.B1(\ram[125][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n175));
   AO22CHD U4014 (.O(n2589), 
	.B2(n303), 
	.B1(\ram[125][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n175));
   AO22CHD U4015 (.O(n2590), 
	.B2(n303), 
	.B1(\ram[125][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n175));
   AO22CHD U4016 (.O(n2591), 
	.B2(n303), 
	.B1(\ram[125][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n175));
   AO22CHD U4017 (.O(n2592), 
	.B2(n303), 
	.B1(\ram[125][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n175));
   AO22CHD U4018 (.O(n2593), 
	.B2(n303), 
	.B1(\ram[125][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n175));
   AO22CHD U4019 (.O(n2594), 
	.B2(n303), 
	.B1(\ram[125][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n175));
   AO22CHD U4020 (.O(n2595), 
	.B2(n303), 
	.B1(\ram[125][13] ), 
	.A2(n21), 
	.A1(n175));
   AO22CHD U4021 (.O(n2596), 
	.B2(n303), 
	.B1(\ram[125][14] ), 
	.A2(n22), 
	.A1(n175));
   AO22CHD U4022 (.O(n2597), 
	.B2(n303), 
	.B1(\ram[125][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n175));
   AO22CHD U4023 (.O(n2598), 
	.B2(n305), 
	.B1(\ram[126][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n177));
   AO22CHD U4024 (.O(n2599), 
	.B2(n305), 
	.B1(\ram[126][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n177));
   AO22CHD U4025 (.O(n2600), 
	.B2(n305), 
	.B1(\ram[126][2] ), 
	.A2(n10), 
	.A1(n177));
   AO22CHD U4026 (.O(n2601), 
	.B2(n305), 
	.B1(\ram[126][3] ), 
	.A2(n11), 
	.A1(n177));
   AO22CHD U4027 (.O(n2602), 
	.B2(n305), 
	.B1(\ram[126][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n177));
   AO22CHD U4028 (.O(n2603), 
	.B2(n305), 
	.B1(\ram[126][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n177));
   AO22CHD U4029 (.O(n2604), 
	.B2(n305), 
	.B1(\ram[126][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n177));
   AO22CHD U4030 (.O(n2605), 
	.B2(n305), 
	.B1(\ram[126][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n177));
   AO22CHD U4031 (.O(n2606), 
	.B2(n305), 
	.B1(\ram[126][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n177));
   AO22CHD U4032 (.O(n2607), 
	.B2(n305), 
	.B1(\ram[126][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n177));
   AO22CHD U4033 (.O(n2608), 
	.B2(n305), 
	.B1(\ram[126][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n177));
   AO22CHD U4034 (.O(n2609), 
	.B2(n305), 
	.B1(\ram[126][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n177));
   AO22CHD U4035 (.O(n2610), 
	.B2(n305), 
	.B1(\ram[126][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n177));
   AO22CHD U4036 (.O(n2611), 
	.B2(n305), 
	.B1(\ram[126][13] ), 
	.A2(n21), 
	.A1(n177));
   AO22CHD U4037 (.O(n2612), 
	.B2(n305), 
	.B1(\ram[126][14] ), 
	.A2(n22), 
	.A1(n177));
   AO22CHD U4038 (.O(n2613), 
	.B2(n305), 
	.B1(\ram[126][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n177));
   AO22CHD U4039 (.O(n2614), 
	.B2(n307), 
	.B1(\ram[127][0] ), 
	.A2(n6), 
	.A1(n178));
   AO22CHD U4040 (.O(n2615), 
	.B2(n307), 
	.B1(\ram[127][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n178));
   AO22CHD U4041 (.O(n2616), 
	.B2(n307), 
	.B1(\ram[127][2] ), 
	.A2(n10), 
	.A1(n178));
   AO22CHD U4042 (.O(n2617), 
	.B2(n307), 
	.B1(\ram[127][3] ), 
	.A2(n11), 
	.A1(n178));
   AO22CHD U4043 (.O(n2618), 
	.B2(n307), 
	.B1(\ram[127][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n178));
   AO22CHD U4044 (.O(n2619), 
	.B2(n307), 
	.B1(\ram[127][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n178));
   AO22CHD U4045 (.O(n2620), 
	.B2(n307), 
	.B1(\ram[127][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n178));
   AO22CHD U4046 (.O(n2621), 
	.B2(n307), 
	.B1(\ram[127][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n178));
   AO22CHD U4047 (.O(n2622), 
	.B2(n307), 
	.B1(\ram[127][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n178));
   AO22CHD U4048 (.O(n2623), 
	.B2(n307), 
	.B1(\ram[127][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n178));
   AO22CHD U4049 (.O(n2624), 
	.B2(n307), 
	.B1(\ram[127][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n178));
   AO22CHD U4050 (.O(n2625), 
	.B2(n307), 
	.B1(\ram[127][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n178));
   AO22CHD U4051 (.O(n2626), 
	.B2(n307), 
	.B1(\ram[127][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n178));
   AO22CHD U4052 (.O(n2627), 
	.B2(n307), 
	.B1(\ram[127][13] ), 
	.A2(n21), 
	.A1(n178));
   AO22CHD U4053 (.O(n2628), 
	.B2(n307), 
	.B1(\ram[127][14] ), 
	.A2(n22), 
	.A1(n178));
   AO22CHD U4054 (.O(n2629), 
	.B2(n307), 
	.B1(\ram[127][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n178));
   AO22CHD U4055 (.O(n2630), 
	.B2(n309), 
	.B1(\ram[128][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n180));
   AO22CHD U4056 (.O(n2631), 
	.B2(n309), 
	.B1(\ram[128][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n180));
   AO22CHD U4057 (.O(n2632), 
	.B2(n309), 
	.B1(\ram[128][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n180));
   AO22CHD U4058 (.O(n2633), 
	.B2(n309), 
	.B1(\ram[128][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n180));
   AO22CHD U4059 (.O(n2634), 
	.B2(n309), 
	.B1(\ram[128][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n180));
   AO22CHD U4060 (.O(n2635), 
	.B2(n309), 
	.B1(\ram[128][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n180));
   AO22CHD U4061 (.O(n2636), 
	.B2(n309), 
	.B1(\ram[128][6] ), 
	.A2(n14), 
	.A1(n180));
   AO22CHD U4062 (.O(n2637), 
	.B2(n309), 
	.B1(\ram[128][7] ), 
	.A2(n15), 
	.A1(n180));
   AO22CHD U4063 (.O(n2638), 
	.B2(n309), 
	.B1(\ram[128][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n180));
   AO22CHD U4064 (.O(n2639), 
	.B2(n309), 
	.B1(\ram[128][9] ), 
	.A2(n17), 
	.A1(n180));
   AO22CHD U4065 (.O(n2640), 
	.B2(n309), 
	.B1(\ram[128][10] ), 
	.A2(n18), 
	.A1(n180));
   AO22CHD U4066 (.O(n2641), 
	.B2(n309), 
	.B1(\ram[128][11] ), 
	.A2(n19), 
	.A1(n180));
   AO22CHD U4067 (.O(n2642), 
	.B2(n309), 
	.B1(\ram[128][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n180));
   AO22CHD U4068 (.O(n2643), 
	.B2(n309), 
	.B1(\ram[128][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n180));
   AO22CHD U4069 (.O(n2644), 
	.B2(n309), 
	.B1(\ram[128][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n180));
   AO22CHD U4070 (.O(n2645), 
	.B2(n309), 
	.B1(\ram[128][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n180));
   AO22CHD U4071 (.O(n2646), 
	.B2(n312), 
	.B1(\ram[129][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n182));
   AO22CHD U4072 (.O(n2647), 
	.B2(n312), 
	.B1(\ram[129][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n182));
   AO22CHD U4073 (.O(n2648), 
	.B2(n312), 
	.B1(\ram[129][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n182));
   AO22CHD U4074 (.O(n2649), 
	.B2(n312), 
	.B1(\ram[129][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n182));
   AO22CHD U4075 (.O(n2650), 
	.B2(n312), 
	.B1(\ram[129][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n182));
   AO22CHD U4076 (.O(n2651), 
	.B2(n312), 
	.B1(\ram[129][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n182));
   AO22CHD U4077 (.O(n2652), 
	.B2(n312), 
	.B1(\ram[129][6] ), 
	.A2(n14), 
	.A1(n182));
   AO22CHD U4078 (.O(n2653), 
	.B2(n312), 
	.B1(\ram[129][7] ), 
	.A2(n15), 
	.A1(n182));
   AO22CHD U4079 (.O(n2654), 
	.B2(n312), 
	.B1(\ram[129][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n182));
   AO22CHD U4080 (.O(n2655), 
	.B2(n312), 
	.B1(\ram[129][9] ), 
	.A2(n17), 
	.A1(n182));
   AO22CHD U4081 (.O(n2656), 
	.B2(n312), 
	.B1(\ram[129][10] ), 
	.A2(n18), 
	.A1(n182));
   AO22CHD U4082 (.O(n2657), 
	.B2(n312), 
	.B1(\ram[129][11] ), 
	.A2(n19), 
	.A1(n182));
   AO22CHD U4083 (.O(n2658), 
	.B2(n312), 
	.B1(\ram[129][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n182));
   AO22CHD U4084 (.O(n2659), 
	.B2(n312), 
	.B1(\ram[129][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n182));
   AO22CHD U4085 (.O(n2660), 
	.B2(n312), 
	.B1(\ram[129][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n182));
   AO22CHD U4086 (.O(n2661), 
	.B2(n312), 
	.B1(\ram[129][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n182));
   AO22CHD U4087 (.O(n2662), 
	.B2(n314), 
	.B1(\ram[130][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n184));
   AO22CHD U4088 (.O(n2663), 
	.B2(n314), 
	.B1(\ram[130][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n184));
   AO22CHD U4089 (.O(n2664), 
	.B2(n314), 
	.B1(\ram[130][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n184));
   AO22CHD U4090 (.O(n2665), 
	.B2(n314), 
	.B1(\ram[130][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n184));
   AO22CHD U4091 (.O(n2666), 
	.B2(n314), 
	.B1(\ram[130][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n184));
   AO22CHD U4092 (.O(n2667), 
	.B2(n314), 
	.B1(\ram[130][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n184));
   AO22CHD U4093 (.O(n2668), 
	.B2(n314), 
	.B1(\ram[130][6] ), 
	.A2(n14), 
	.A1(n184));
   AO22CHD U4094 (.O(n2669), 
	.B2(n314), 
	.B1(\ram[130][7] ), 
	.A2(n15), 
	.A1(n184));
   AO22CHD U4095 (.O(n2670), 
	.B2(n314), 
	.B1(\ram[130][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n184));
   AO22CHD U4096 (.O(n2671), 
	.B2(n314), 
	.B1(\ram[130][9] ), 
	.A2(n17), 
	.A1(n184));
   AO22CHD U4097 (.O(n2672), 
	.B2(n314), 
	.B1(\ram[130][10] ), 
	.A2(n18), 
	.A1(n184));
   AO22CHD U4098 (.O(n2673), 
	.B2(n314), 
	.B1(\ram[130][11] ), 
	.A2(n19), 
	.A1(n184));
   AO22CHD U4099 (.O(n2674), 
	.B2(n314), 
	.B1(\ram[130][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n184));
   AO22CHD U4100 (.O(n2675), 
	.B2(n314), 
	.B1(\ram[130][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n184));
   AO22CHD U4101 (.O(n2676), 
	.B2(n314), 
	.B1(\ram[130][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n184));
   AO22CHD U4102 (.O(n2677), 
	.B2(n314), 
	.B1(\ram[130][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n184));
   AO22CHD U4103 (.O(n2678), 
	.B2(n316), 
	.B1(\ram[131][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n186));
   AO22CHD U4104 (.O(n2679), 
	.B2(n316), 
	.B1(\ram[131][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n186));
   AO22CHD U4105 (.O(n2680), 
	.B2(n316), 
	.B1(\ram[131][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n186));
   AO22CHD U4106 (.O(n2681), 
	.B2(n316), 
	.B1(\ram[131][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n186));
   AO22CHD U4107 (.O(n2682), 
	.B2(n316), 
	.B1(\ram[131][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n186));
   AO22CHD U4108 (.O(n2683), 
	.B2(n316), 
	.B1(\ram[131][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n186));
   AO22CHD U4109 (.O(n2684), 
	.B2(n316), 
	.B1(\ram[131][6] ), 
	.A2(n14), 
	.A1(n186));
   AO22CHD U4110 (.O(n2685), 
	.B2(n316), 
	.B1(\ram[131][7] ), 
	.A2(n15), 
	.A1(n186));
   AO22CHD U4111 (.O(n2686), 
	.B2(n316), 
	.B1(\ram[131][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n186));
   AO22CHD U4112 (.O(n2687), 
	.B2(n316), 
	.B1(\ram[131][9] ), 
	.A2(n17), 
	.A1(n186));
   AO22CHD U4113 (.O(n2688), 
	.B2(n316), 
	.B1(\ram[131][10] ), 
	.A2(n18), 
	.A1(n186));
   AO22CHD U4114 (.O(n2689), 
	.B2(n316), 
	.B1(\ram[131][11] ), 
	.A2(n19), 
	.A1(n186));
   AO22CHD U4115 (.O(n2690), 
	.B2(n316), 
	.B1(\ram[131][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n186));
   AO22CHD U4116 (.O(n2691), 
	.B2(n316), 
	.B1(\ram[131][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n186));
   AO22CHD U4117 (.O(n2692), 
	.B2(n316), 
	.B1(\ram[131][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n186));
   AO22CHD U4118 (.O(n2693), 
	.B2(n316), 
	.B1(\ram[131][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n186));
   AO22CHD U4119 (.O(n2694), 
	.B2(n318), 
	.B1(\ram[132][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n188));
   AO22CHD U4120 (.O(n2695), 
	.B2(n318), 
	.B1(\ram[132][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n188));
   AO22CHD U4121 (.O(n2696), 
	.B2(n318), 
	.B1(\ram[132][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n188));
   AO22CHD U4122 (.O(n2697), 
	.B2(n318), 
	.B1(\ram[132][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n188));
   AO22CHD U4123 (.O(n2698), 
	.B2(n318), 
	.B1(\ram[132][4] ), 
	.A2(n12), 
	.A1(n188));
   AO22CHD U4124 (.O(n2699), 
	.B2(n318), 
	.B1(\ram[132][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n188));
   AO22CHD U4125 (.O(n2700), 
	.B2(n318), 
	.B1(\ram[132][6] ), 
	.A2(n14), 
	.A1(n188));
   AO22CHD U4126 (.O(n2701), 
	.B2(n318), 
	.B1(\ram[132][7] ), 
	.A2(n15), 
	.A1(n188));
   AO22CHD U4127 (.O(n2702), 
	.B2(n318), 
	.B1(\ram[132][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n188));
   AO22CHD U4128 (.O(n2703), 
	.B2(n318), 
	.B1(\ram[132][9] ), 
	.A2(n17), 
	.A1(n188));
   AO22CHD U4129 (.O(n2704), 
	.B2(n318), 
	.B1(\ram[132][10] ), 
	.A2(n18), 
	.A1(n188));
   AO22CHD U4130 (.O(n2705), 
	.B2(n318), 
	.B1(\ram[132][11] ), 
	.A2(n19), 
	.A1(n188));
   AO22CHD U4131 (.O(n2706), 
	.B2(n318), 
	.B1(\ram[132][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n188));
   AO22CHD U4132 (.O(n2707), 
	.B2(n318), 
	.B1(\ram[132][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n188));
   AO22CHD U4133 (.O(n2708), 
	.B2(n318), 
	.B1(\ram[132][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n188));
   AO22CHD U4134 (.O(n2709), 
	.B2(n318), 
	.B1(\ram[132][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n188));
   AO22CHD U4135 (.O(n2710), 
	.B2(n320), 
	.B1(\ram[133][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n190));
   AO22CHD U4136 (.O(n2711), 
	.B2(n320), 
	.B1(\ram[133][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n190));
   AO22CHD U4137 (.O(n2712), 
	.B2(n320), 
	.B1(\ram[133][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n190));
   AO22CHD U4138 (.O(n2713), 
	.B2(n320), 
	.B1(\ram[133][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n190));
   AO22CHD U4139 (.O(n2714), 
	.B2(n320), 
	.B1(\ram[133][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n190));
   AO22CHD U4140 (.O(n2715), 
	.B2(n320), 
	.B1(\ram[133][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n190));
   AO22CHD U4141 (.O(n2716), 
	.B2(n320), 
	.B1(\ram[133][6] ), 
	.A2(n14), 
	.A1(n190));
   AO22CHD U4142 (.O(n2717), 
	.B2(n320), 
	.B1(\ram[133][7] ), 
	.A2(n15), 
	.A1(n190));
   AO22CHD U4143 (.O(n2718), 
	.B2(n320), 
	.B1(\ram[133][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n190));
   AO22CHD U4144 (.O(n2719), 
	.B2(n320), 
	.B1(\ram[133][9] ), 
	.A2(n17), 
	.A1(n190));
   AO22CHD U4145 (.O(n2720), 
	.B2(n320), 
	.B1(\ram[133][10] ), 
	.A2(n18), 
	.A1(n190));
   AO22CHD U4146 (.O(n2721), 
	.B2(n320), 
	.B1(\ram[133][11] ), 
	.A2(n19), 
	.A1(n190));
   AO22CHD U4147 (.O(n2722), 
	.B2(n320), 
	.B1(\ram[133][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n190));
   AO22CHD U4148 (.O(n2723), 
	.B2(n320), 
	.B1(\ram[133][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n190));
   AO22CHD U4149 (.O(n2724), 
	.B2(n320), 
	.B1(\ram[133][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n190));
   AO22CHD U4150 (.O(n2725), 
	.B2(n320), 
	.B1(\ram[133][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n190));
   AO22CHD U4151 (.O(n2726), 
	.B2(n322), 
	.B1(\ram[134][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n192));
   AO22CHD U4152 (.O(n2727), 
	.B2(n322), 
	.B1(\ram[134][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n192));
   AO22CHD U4153 (.O(n2728), 
	.B2(n322), 
	.B1(\ram[134][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n192));
   AO22CHD U4154 (.O(n2729), 
	.B2(n322), 
	.B1(\ram[134][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n192));
   AO22CHD U4155 (.O(n2730), 
	.B2(n322), 
	.B1(\ram[134][4] ), 
	.A2(n12), 
	.A1(n192));
   AO22CHD U4156 (.O(n2731), 
	.B2(n322), 
	.B1(\ram[134][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n192));
   AO22CHD U4157 (.O(n2732), 
	.B2(n322), 
	.B1(\ram[134][6] ), 
	.A2(n14), 
	.A1(n192));
   AO22CHD U4158 (.O(n2733), 
	.B2(n322), 
	.B1(\ram[134][7] ), 
	.A2(n15), 
	.A1(n192));
   AO22CHD U4159 (.O(n2734), 
	.B2(n322), 
	.B1(\ram[134][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n192));
   AO22CHD U4160 (.O(n2735), 
	.B2(n322), 
	.B1(\ram[134][9] ), 
	.A2(n17), 
	.A1(n192));
   AO22CHD U4161 (.O(n2736), 
	.B2(n322), 
	.B1(\ram[134][10] ), 
	.A2(n18), 
	.A1(n192));
   AO22CHD U4162 (.O(n2737), 
	.B2(n322), 
	.B1(\ram[134][11] ), 
	.A2(n19), 
	.A1(n192));
   AO22CHD U4163 (.O(n2738), 
	.B2(n322), 
	.B1(\ram[134][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n192));
   AO22CHD U4164 (.O(n2739), 
	.B2(n322), 
	.B1(\ram[134][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n192));
   AO22CHD U4165 (.O(n2740), 
	.B2(n322), 
	.B1(\ram[134][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n192));
   AO22CHD U4166 (.O(n2741), 
	.B2(n322), 
	.B1(\ram[134][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n192));
   AO22CHD U4167 (.O(n2742), 
	.B2(n324), 
	.B1(\ram[135][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n194));
   AO22CHD U4168 (.O(n2743), 
	.B2(n324), 
	.B1(\ram[135][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n194));
   AO22CHD U4169 (.O(n2744), 
	.B2(n324), 
	.B1(\ram[135][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n194));
   AO22CHD U4170 (.O(n2745), 
	.B2(n324), 
	.B1(\ram[135][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n194));
   AO22CHD U4171 (.O(n2746), 
	.B2(n324), 
	.B1(\ram[135][4] ), 
	.A2(n12), 
	.A1(n194));
   AO22CHD U4172 (.O(n2747), 
	.B2(n324), 
	.B1(\ram[135][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n194));
   AO22CHD U4173 (.O(n2748), 
	.B2(n324), 
	.B1(\ram[135][6] ), 
	.A2(n14), 
	.A1(n194));
   AO22CHD U4174 (.O(n2749), 
	.B2(n324), 
	.B1(\ram[135][7] ), 
	.A2(n15), 
	.A1(n194));
   AO22CHD U4175 (.O(n2750), 
	.B2(n324), 
	.B1(\ram[135][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n194));
   AO22CHD U4176 (.O(n2751), 
	.B2(n324), 
	.B1(\ram[135][9] ), 
	.A2(n17), 
	.A1(n194));
   AO22CHD U4177 (.O(n2752), 
	.B2(n324), 
	.B1(\ram[135][10] ), 
	.A2(n18), 
	.A1(n194));
   AO22CHD U4178 (.O(n2753), 
	.B2(n324), 
	.B1(\ram[135][11] ), 
	.A2(n19), 
	.A1(n194));
   AO22CHD U4179 (.O(n2754), 
	.B2(n324), 
	.B1(\ram[135][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n194));
   AO22CHD U4180 (.O(n2755), 
	.B2(n324), 
	.B1(\ram[135][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n194));
   AO22CHD U4181 (.O(n2756), 
	.B2(n324), 
	.B1(\ram[135][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n194));
   AO22CHD U4182 (.O(n2757), 
	.B2(n324), 
	.B1(\ram[135][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n194));
   AO22CHD U4183 (.O(n2758), 
	.B2(n326), 
	.B1(\ram[136][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n196));
   AO22CHD U4184 (.O(n2759), 
	.B2(n326), 
	.B1(\ram[136][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n196));
   AO22CHD U4185 (.O(n2760), 
	.B2(n326), 
	.B1(\ram[136][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n196));
   AO22CHD U4186 (.O(n2761), 
	.B2(n326), 
	.B1(\ram[136][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n196));
   AO22CHD U4187 (.O(n2762), 
	.B2(n326), 
	.B1(\ram[136][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n196));
   AO22CHD U4188 (.O(n2763), 
	.B2(n326), 
	.B1(\ram[136][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n196));
   AO22CHD U4189 (.O(n2764), 
	.B2(n326), 
	.B1(\ram[136][6] ), 
	.A2(n14), 
	.A1(n196));
   AO22CHD U4190 (.O(n2765), 
	.B2(n326), 
	.B1(\ram[136][7] ), 
	.A2(n15), 
	.A1(n196));
   AO22CHD U4191 (.O(n2766), 
	.B2(n326), 
	.B1(\ram[136][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n196));
   AO22CHD U4192 (.O(n2767), 
	.B2(n326), 
	.B1(\ram[136][9] ), 
	.A2(n17), 
	.A1(n196));
   AO22CHD U4193 (.O(n2768), 
	.B2(n326), 
	.B1(\ram[136][10] ), 
	.A2(n18), 
	.A1(n196));
   AO22CHD U4194 (.O(n2769), 
	.B2(n326), 
	.B1(\ram[136][11] ), 
	.A2(n19), 
	.A1(n196));
   AO22CHD U4195 (.O(n2770), 
	.B2(n326), 
	.B1(\ram[136][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n196));
   AO22CHD U4196 (.O(n2771), 
	.B2(n326), 
	.B1(\ram[136][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n196));
   AO22CHD U4197 (.O(n2772), 
	.B2(n326), 
	.B1(\ram[136][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n196));
   AO22CHD U4198 (.O(n2773), 
	.B2(n326), 
	.B1(\ram[136][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n196));
   AO22CHD U4199 (.O(n2774), 
	.B2(n328), 
	.B1(\ram[137][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n198));
   AO22CHD U4200 (.O(n2775), 
	.B2(n328), 
	.B1(\ram[137][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n198));
   AO22CHD U4201 (.O(n2776), 
	.B2(n328), 
	.B1(\ram[137][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n198));
   AO22CHD U4202 (.O(n2777), 
	.B2(n328), 
	.B1(\ram[137][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n198));
   AO22CHD U4203 (.O(n2778), 
	.B2(n328), 
	.B1(\ram[137][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n198));
   AO22CHD U4204 (.O(n2779), 
	.B2(n328), 
	.B1(\ram[137][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n198));
   AO22CHD U4205 (.O(n2780), 
	.B2(n328), 
	.B1(\ram[137][6] ), 
	.A2(n14), 
	.A1(n198));
   AO22CHD U4206 (.O(n2781), 
	.B2(n328), 
	.B1(\ram[137][7] ), 
	.A2(n15), 
	.A1(n198));
   AO22CHD U4207 (.O(n2782), 
	.B2(n328), 
	.B1(\ram[137][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n198));
   AO22CHD U4208 (.O(n2783), 
	.B2(n328), 
	.B1(\ram[137][9] ), 
	.A2(n17), 
	.A1(n198));
   AO22CHD U4209 (.O(n2784), 
	.B2(n328), 
	.B1(\ram[137][10] ), 
	.A2(n18), 
	.A1(n198));
   AO22CHD U4210 (.O(n2785), 
	.B2(n328), 
	.B1(\ram[137][11] ), 
	.A2(n19), 
	.A1(n198));
   AO22CHD U4211 (.O(n2786), 
	.B2(n328), 
	.B1(\ram[137][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n198));
   AO22CHD U4212 (.O(n2787), 
	.B2(n328), 
	.B1(\ram[137][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n198));
   AO22CHD U4213 (.O(n2788), 
	.B2(n328), 
	.B1(\ram[137][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n198));
   AO22CHD U4214 (.O(n2789), 
	.B2(n328), 
	.B1(\ram[137][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n198));
   AO22CHD U4215 (.O(n2790), 
	.B2(n330), 
	.B1(\ram[138][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n200));
   AO22CHD U4216 (.O(n2791), 
	.B2(n330), 
	.B1(\ram[138][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n200));
   AO22CHD U4217 (.O(n2792), 
	.B2(n330), 
	.B1(\ram[138][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n200));
   AO22CHD U4218 (.O(n2793), 
	.B2(n330), 
	.B1(\ram[138][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n200));
   AO22CHD U4219 (.O(n2794), 
	.B2(n330), 
	.B1(\ram[138][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n200));
   AO22CHD U4220 (.O(n2795), 
	.B2(n330), 
	.B1(\ram[138][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n200));
   AO22CHD U4221 (.O(n2796), 
	.B2(n330), 
	.B1(\ram[138][6] ), 
	.A2(n14), 
	.A1(n200));
   AO22CHD U4222 (.O(n2797), 
	.B2(n330), 
	.B1(\ram[138][7] ), 
	.A2(n15), 
	.A1(n200));
   AO22CHD U4223 (.O(n2798), 
	.B2(n330), 
	.B1(\ram[138][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n200));
   AO22CHD U4224 (.O(n2799), 
	.B2(n330), 
	.B1(\ram[138][9] ), 
	.A2(n17), 
	.A1(n200));
   AO22CHD U4225 (.O(n2800), 
	.B2(n330), 
	.B1(\ram[138][10] ), 
	.A2(n18), 
	.A1(n200));
   AO22CHD U4226 (.O(n2801), 
	.B2(n330), 
	.B1(\ram[138][11] ), 
	.A2(n19), 
	.A1(n200));
   AO22CHD U4227 (.O(n2802), 
	.B2(n330), 
	.B1(\ram[138][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n200));
   AO22CHD U4228 (.O(n2803), 
	.B2(n330), 
	.B1(\ram[138][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n200));
   AO22CHD U4229 (.O(n2804), 
	.B2(n330), 
	.B1(\ram[138][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n200));
   AO22CHD U4230 (.O(n2805), 
	.B2(n330), 
	.B1(\ram[138][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n200));
   AO22CHD U4231 (.O(n2806), 
	.B2(n332), 
	.B1(\ram[139][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n202));
   AO22CHD U4232 (.O(n2807), 
	.B2(n332), 
	.B1(\ram[139][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n202));
   AO22CHD U4233 (.O(n2808), 
	.B2(n332), 
	.B1(\ram[139][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n202));
   AO22CHD U4234 (.O(n2809), 
	.B2(n332), 
	.B1(\ram[139][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n202));
   AO22CHD U4235 (.O(n2810), 
	.B2(n332), 
	.B1(\ram[139][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n202));
   AO22CHD U4236 (.O(n2811), 
	.B2(n332), 
	.B1(\ram[139][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n202));
   AO22CHD U4237 (.O(n2812), 
	.B2(n332), 
	.B1(\ram[139][6] ), 
	.A2(n14), 
	.A1(n202));
   AO22CHD U4238 (.O(n2813), 
	.B2(n332), 
	.B1(\ram[139][7] ), 
	.A2(n15), 
	.A1(n202));
   AO22CHD U4239 (.O(n2814), 
	.B2(n332), 
	.B1(\ram[139][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n202));
   AO22CHD U4240 (.O(n2815), 
	.B2(n332), 
	.B1(\ram[139][9] ), 
	.A2(n17), 
	.A1(n202));
   AO22CHD U4241 (.O(n2816), 
	.B2(n332), 
	.B1(\ram[139][10] ), 
	.A2(n18), 
	.A1(n202));
   AO22CHD U4242 (.O(n2817), 
	.B2(n332), 
	.B1(\ram[139][11] ), 
	.A2(n19), 
	.A1(n202));
   AO22CHD U4243 (.O(n2818), 
	.B2(n332), 
	.B1(\ram[139][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n202));
   AO22CHD U4244 (.O(n2819), 
	.B2(n332), 
	.B1(\ram[139][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n202));
   AO22CHD U4245 (.O(n2820), 
	.B2(n332), 
	.B1(\ram[139][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n202));
   AO22CHD U4246 (.O(n2821), 
	.B2(n332), 
	.B1(\ram[139][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n202));
   AO22CHD U4247 (.O(n2822), 
	.B2(n334), 
	.B1(\ram[140][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n204));
   AO22CHD U4248 (.O(n2823), 
	.B2(n334), 
	.B1(\ram[140][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n204));
   AO22CHD U4249 (.O(n2824), 
	.B2(n334), 
	.B1(\ram[140][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n204));
   AO22CHD U4250 (.O(n2825), 
	.B2(n334), 
	.B1(\ram[140][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n204));
   AO22CHD U4251 (.O(n2826), 
	.B2(n334), 
	.B1(\ram[140][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n204));
   AO22CHD U4252 (.O(n2827), 
	.B2(n334), 
	.B1(\ram[140][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n204));
   AO22CHD U4253 (.O(n2828), 
	.B2(n334), 
	.B1(\ram[140][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n204));
   AO22CHD U4254 (.O(n2829), 
	.B2(n334), 
	.B1(\ram[140][7] ), 
	.A2(n15), 
	.A1(n204));
   AO22CHD U4255 (.O(n2830), 
	.B2(n334), 
	.B1(\ram[140][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n204));
   AO22CHD U4256 (.O(n2831), 
	.B2(n334), 
	.B1(\ram[140][9] ), 
	.A2(n17), 
	.A1(n204));
   AO22CHD U4257 (.O(n2832), 
	.B2(n334), 
	.B1(\ram[140][10] ), 
	.A2(n18), 
	.A1(n204));
   AO22CHD U4258 (.O(n2833), 
	.B2(n334), 
	.B1(\ram[140][11] ), 
	.A2(n19), 
	.A1(n204));
   AO22CHD U4259 (.O(n2834), 
	.B2(n334), 
	.B1(\ram[140][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n204));
   AO22CHD U4260 (.O(n2835), 
	.B2(n334), 
	.B1(\ram[140][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n204));
   AO22CHD U4261 (.O(n2836), 
	.B2(n334), 
	.B1(\ram[140][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n204));
   AO22CHD U4262 (.O(n2837), 
	.B2(n334), 
	.B1(\ram[140][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n204));
   AO22CHD U4263 (.O(n2838), 
	.B2(n336), 
	.B1(\ram[141][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n206));
   AO22CHD U4264 (.O(n2839), 
	.B2(n336), 
	.B1(\ram[141][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n206));
   AO22CHD U4265 (.O(n2840), 
	.B2(n336), 
	.B1(\ram[141][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n206));
   AO22CHD U4266 (.O(n2841), 
	.B2(n336), 
	.B1(\ram[141][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n206));
   AO22CHD U4267 (.O(n2842), 
	.B2(n336), 
	.B1(\ram[141][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n206));
   AO22CHD U4268 (.O(n2843), 
	.B2(n336), 
	.B1(\ram[141][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n206));
   AO22CHD U4269 (.O(n2844), 
	.B2(n336), 
	.B1(\ram[141][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n206));
   AO22CHD U4270 (.O(n2845), 
	.B2(n336), 
	.B1(\ram[141][7] ), 
	.A2(n15), 
	.A1(n206));
   AO22CHD U4271 (.O(n2846), 
	.B2(n336), 
	.B1(\ram[141][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n206));
   AO22CHD U4272 (.O(n2847), 
	.B2(n336), 
	.B1(\ram[141][9] ), 
	.A2(n17), 
	.A1(n206));
   AO22CHD U4273 (.O(n2848), 
	.B2(n336), 
	.B1(\ram[141][10] ), 
	.A2(n18), 
	.A1(n206));
   AO22CHD U4274 (.O(n2849), 
	.B2(n336), 
	.B1(\ram[141][11] ), 
	.A2(n19), 
	.A1(n206));
   AO22CHD U4275 (.O(n2850), 
	.B2(n336), 
	.B1(\ram[141][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n206));
   AO22CHD U4276 (.O(n2851), 
	.B2(n336), 
	.B1(\ram[141][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n206));
   AO22CHD U4277 (.O(n2852), 
	.B2(n336), 
	.B1(\ram[141][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n206));
   AO22CHD U4278 (.O(n2853), 
	.B2(n336), 
	.B1(\ram[141][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n206));
   AO22CHD U4279 (.O(n2854), 
	.B2(n338), 
	.B1(\ram[142][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n209));
   AO22CHD U4280 (.O(n2855), 
	.B2(n338), 
	.B1(\ram[142][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n209));
   AO22CHD U4281 (.O(n2856), 
	.B2(n338), 
	.B1(\ram[142][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n209));
   AO22CHD U4282 (.O(n2857), 
	.B2(n338), 
	.B1(\ram[142][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n209));
   AO22CHD U4283 (.O(n2858), 
	.B2(n338), 
	.B1(\ram[142][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n209));
   AO22CHD U4284 (.O(n2859), 
	.B2(n338), 
	.B1(\ram[142][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n209));
   AO22CHD U4285 (.O(n2860), 
	.B2(n338), 
	.B1(\ram[142][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n209));
   AO22CHD U4286 (.O(n2861), 
	.B2(n338), 
	.B1(\ram[142][7] ), 
	.A2(n15), 
	.A1(n209));
   AO22CHD U4287 (.O(n2862), 
	.B2(n338), 
	.B1(\ram[142][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n209));
   AO22CHD U4288 (.O(n2863), 
	.B2(n338), 
	.B1(\ram[142][9] ), 
	.A2(n17), 
	.A1(n209));
   AO22CHD U4289 (.O(n2864), 
	.B2(n338), 
	.B1(\ram[142][10] ), 
	.A2(n18), 
	.A1(n209));
   AO22CHD U4290 (.O(n2865), 
	.B2(n338), 
	.B1(\ram[142][11] ), 
	.A2(n19), 
	.A1(n209));
   AO22CHD U4291 (.O(n2866), 
	.B2(n338), 
	.B1(\ram[142][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n209));
   AO22CHD U4292 (.O(n2867), 
	.B2(n338), 
	.B1(\ram[142][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n209));
   AO22CHD U4293 (.O(n2868), 
	.B2(n338), 
	.B1(\ram[142][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n209));
   AO22CHD U4294 (.O(n2869), 
	.B2(n338), 
	.B1(\ram[142][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n209));
   AO22CHD U4295 (.O(n2870), 
	.B2(n340), 
	.B1(\ram[143][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n211));
   AO22CHD U4296 (.O(n2871), 
	.B2(n340), 
	.B1(\ram[143][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n211));
   AO22CHD U4297 (.O(n2872), 
	.B2(n340), 
	.B1(\ram[143][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n211));
   AO22CHD U4298 (.O(n2873), 
	.B2(n340), 
	.B1(\ram[143][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n211));
   AO22CHD U4299 (.O(n2874), 
	.B2(n340), 
	.B1(\ram[143][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n211));
   AO22CHD U4300 (.O(n2875), 
	.B2(n340), 
	.B1(\ram[143][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n211));
   AO22CHD U4301 (.O(n2876), 
	.B2(n340), 
	.B1(\ram[143][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n211));
   AO22CHD U4302 (.O(n2877), 
	.B2(n340), 
	.B1(\ram[143][7] ), 
	.A2(n15), 
	.A1(n211));
   AO22CHD U4303 (.O(n2878), 
	.B2(n340), 
	.B1(\ram[143][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n211));
   AO22CHD U4304 (.O(n2879), 
	.B2(n340), 
	.B1(\ram[143][9] ), 
	.A2(n17), 
	.A1(n211));
   AO22CHD U4305 (.O(n2880), 
	.B2(n340), 
	.B1(\ram[143][10] ), 
	.A2(n18), 
	.A1(n211));
   AO22CHD U4306 (.O(n2881), 
	.B2(n340), 
	.B1(\ram[143][11] ), 
	.A2(n19), 
	.A1(n211));
   AO22CHD U4307 (.O(n2882), 
	.B2(n340), 
	.B1(\ram[143][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n211));
   AO22CHD U4308 (.O(n2883), 
	.B2(n340), 
	.B1(\ram[143][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n211));
   AO22CHD U4309 (.O(n2884), 
	.B2(n340), 
	.B1(\ram[143][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n211));
   AO22CHD U4310 (.O(n2885), 
	.B2(n340), 
	.B1(\ram[143][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n211));
   AO22CHD U4311 (.O(n2886), 
	.B2(n343), 
	.B1(\ram[144][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n212));
   AO22CHD U4312 (.O(n2887), 
	.B2(n343), 
	.B1(\ram[144][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n212));
   AO22CHD U4313 (.O(n2888), 
	.B2(n343), 
	.B1(\ram[144][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n212));
   AO22CHD U4314 (.O(n2889), 
	.B2(n343), 
	.B1(\ram[144][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n212));
   AO22CHD U4315 (.O(n2890), 
	.B2(n343), 
	.B1(\ram[144][4] ), 
	.A2(n12), 
	.A1(n212));
   AO22CHD U4316 (.O(n2891), 
	.B2(n343), 
	.B1(\ram[144][5] ), 
	.A2(n13), 
	.A1(n212));
   AO22CHD U4317 (.O(n2892), 
	.B2(n343), 
	.B1(\ram[144][6] ), 
	.A2(n14), 
	.A1(n212));
   AO22CHD U4318 (.O(n2893), 
	.B2(n343), 
	.B1(\ram[144][7] ), 
	.A2(n15), 
	.A1(n212));
   AO22CHD U4319 (.O(n2894), 
	.B2(n343), 
	.B1(\ram[144][8] ), 
	.A2(n16), 
	.A1(n212));
   AO22CHD U4320 (.O(n2895), 
	.B2(n343), 
	.B1(\ram[144][9] ), 
	.A2(n17), 
	.A1(n212));
   AO22CHD U4321 (.O(n2896), 
	.B2(n343), 
	.B1(\ram[144][10] ), 
	.A2(n18), 
	.A1(n212));
   AO22CHD U4322 (.O(n2897), 
	.B2(n343), 
	.B1(\ram[144][11] ), 
	.A2(n19), 
	.A1(n212));
   AO22CHD U4323 (.O(n2898), 
	.B2(n343), 
	.B1(\ram[144][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n212));
   AO22CHD U4324 (.O(n2899), 
	.B2(n343), 
	.B1(\ram[144][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n212));
   AO22CHD U4325 (.O(n2900), 
	.B2(n343), 
	.B1(\ram[144][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n212));
   AO22CHD U4326 (.O(n2901), 
	.B2(n343), 
	.B1(\ram[144][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n212));
   AO22CHD U4327 (.O(n2902), 
	.B2(n346), 
	.B1(\ram[145][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n214));
   AO22CHD U4328 (.O(n2903), 
	.B2(n346), 
	.B1(\ram[145][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n214));
   AO22CHD U4329 (.O(n2904), 
	.B2(n346), 
	.B1(\ram[145][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n214));
   AO22CHD U4330 (.O(n2905), 
	.B2(n346), 
	.B1(\ram[145][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n214));
   AO22CHD U4331 (.O(n2906), 
	.B2(n346), 
	.B1(\ram[145][4] ), 
	.A2(n12), 
	.A1(n214));
   AO22CHD U4332 (.O(n2907), 
	.B2(n346), 
	.B1(\ram[145][5] ), 
	.A2(n13), 
	.A1(n214));
   AO22CHD U4333 (.O(n2908), 
	.B2(n346), 
	.B1(\ram[145][6] ), 
	.A2(n14), 
	.A1(n214));
   AO22CHD U4334 (.O(n2909), 
	.B2(n346), 
	.B1(\ram[145][7] ), 
	.A2(n15), 
	.A1(n214));
   AO22CHD U4335 (.O(n2910), 
	.B2(n346), 
	.B1(\ram[145][8] ), 
	.A2(n16), 
	.A1(n214));
   AO22CHD U4336 (.O(n2911), 
	.B2(n346), 
	.B1(\ram[145][9] ), 
	.A2(n17), 
	.A1(n214));
   AO22CHD U4337 (.O(n2912), 
	.B2(n346), 
	.B1(\ram[145][10] ), 
	.A2(n18), 
	.A1(n214));
   AO22CHD U4338 (.O(n2913), 
	.B2(n346), 
	.B1(\ram[145][11] ), 
	.A2(n19), 
	.A1(n214));
   AO22CHD U4339 (.O(n2914), 
	.B2(n346), 
	.B1(\ram[145][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n214));
   AO22CHD U4340 (.O(n2915), 
	.B2(n346), 
	.B1(\ram[145][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n214));
   AO22CHD U4341 (.O(n2916), 
	.B2(n346), 
	.B1(\ram[145][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n214));
   AO22CHD U4342 (.O(n2917), 
	.B2(n346), 
	.B1(\ram[145][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n214));
   AO22CHD U4343 (.O(n2918), 
	.B2(n348), 
	.B1(\ram[146][0] ), 
	.A2(n6), 
	.A1(n216));
   AO22CHD U4344 (.O(n2919), 
	.B2(n348), 
	.B1(\ram[146][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n216));
   AO22CHD U4345 (.O(n2920), 
	.B2(n348), 
	.B1(\ram[146][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n216));
   AO22CHD U4346 (.O(n2921), 
	.B2(n348), 
	.B1(\ram[146][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n216));
   AO22CHD U4347 (.O(n2922), 
	.B2(n348), 
	.B1(\ram[146][4] ), 
	.A2(n12), 
	.A1(n216));
   AO22CHD U4348 (.O(n2923), 
	.B2(n348), 
	.B1(\ram[146][5] ), 
	.A2(n13), 
	.A1(n216));
   AO22CHD U4349 (.O(n2924), 
	.B2(n348), 
	.B1(\ram[146][6] ), 
	.A2(n14), 
	.A1(n216));
   AO22CHD U4350 (.O(n2925), 
	.B2(n348), 
	.B1(\ram[146][7] ), 
	.A2(n15), 
	.A1(n216));
   AO22CHD U4351 (.O(n2926), 
	.B2(n348), 
	.B1(\ram[146][8] ), 
	.A2(n16), 
	.A1(n216));
   AO22CHD U4352 (.O(n2927), 
	.B2(n348), 
	.B1(\ram[146][9] ), 
	.A2(n17), 
	.A1(n216));
   AO22CHD U4353 (.O(n2928), 
	.B2(n348), 
	.B1(\ram[146][10] ), 
	.A2(n18), 
	.A1(n216));
   AO22CHD U4354 (.O(n2929), 
	.B2(n348), 
	.B1(\ram[146][11] ), 
	.A2(n19), 
	.A1(n216));
   AO22CHD U4355 (.O(n2930), 
	.B2(n348), 
	.B1(\ram[146][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n216));
   AO22CHD U4356 (.O(n2931), 
	.B2(n348), 
	.B1(\ram[146][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n216));
   AO22CHD U4357 (.O(n2932), 
	.B2(n348), 
	.B1(\ram[146][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n216));
   AO22CHD U4358 (.O(n2933), 
	.B2(n348), 
	.B1(\ram[146][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n216));
   AO22CHD U4359 (.O(n2934), 
	.B2(n350), 
	.B1(\ram[147][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n218));
   AO22CHD U4360 (.O(n2935), 
	.B2(n350), 
	.B1(\ram[147][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n218));
   AO22CHD U4361 (.O(n2936), 
	.B2(n350), 
	.B1(\ram[147][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n218));
   AO22CHD U4362 (.O(n2937), 
	.B2(n350), 
	.B1(\ram[147][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n218));
   AO22CHD U4363 (.O(n2938), 
	.B2(n350), 
	.B1(\ram[147][4] ), 
	.A2(n12), 
	.A1(n218));
   AO22CHD U4364 (.O(n2939), 
	.B2(n350), 
	.B1(\ram[147][5] ), 
	.A2(n13), 
	.A1(n218));
   AO22CHD U4365 (.O(n2940), 
	.B2(n350), 
	.B1(\ram[147][6] ), 
	.A2(n14), 
	.A1(n218));
   AO22CHD U4366 (.O(n2941), 
	.B2(n350), 
	.B1(\ram[147][7] ), 
	.A2(n15), 
	.A1(n218));
   AO22CHD U4367 (.O(n2942), 
	.B2(n350), 
	.B1(\ram[147][8] ), 
	.A2(n16), 
	.A1(n218));
   AO22CHD U4368 (.O(n2943), 
	.B2(n350), 
	.B1(\ram[147][9] ), 
	.A2(n17), 
	.A1(n218));
   AO22CHD U4369 (.O(n2944), 
	.B2(n350), 
	.B1(\ram[147][10] ), 
	.A2(n18), 
	.A1(n218));
   AO22CHD U4370 (.O(n2945), 
	.B2(n350), 
	.B1(\ram[147][11] ), 
	.A2(n19), 
	.A1(n218));
   AO22CHD U4371 (.O(n2946), 
	.B2(n350), 
	.B1(\ram[147][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n218));
   AO22CHD U4372 (.O(n2947), 
	.B2(n350), 
	.B1(\ram[147][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n218));
   AO22CHD U4373 (.O(n2948), 
	.B2(n350), 
	.B1(\ram[147][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n218));
   AO22CHD U4374 (.O(n2949), 
	.B2(n350), 
	.B1(\ram[147][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n218));
   AO22CHD U4375 (.O(n2950), 
	.B2(n352), 
	.B1(\ram[148][0] ), 
	.A2(n6), 
	.A1(n220));
   AO22CHD U4376 (.O(n2951), 
	.B2(n352), 
	.B1(\ram[148][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n220));
   AO22CHD U4377 (.O(n2952), 
	.B2(n352), 
	.B1(\ram[148][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n220));
   AO22CHD U4378 (.O(n2953), 
	.B2(n352), 
	.B1(\ram[148][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n220));
   AO22CHD U4379 (.O(n2954), 
	.B2(n352), 
	.B1(\ram[148][4] ), 
	.A2(n12), 
	.A1(n220));
   AO22CHD U4380 (.O(n2955), 
	.B2(n352), 
	.B1(\ram[148][5] ), 
	.A2(n13), 
	.A1(n220));
   AO22CHD U4381 (.O(n2956), 
	.B2(n352), 
	.B1(\ram[148][6] ), 
	.A2(n14), 
	.A1(n220));
   AO22CHD U4382 (.O(n2957), 
	.B2(n352), 
	.B1(\ram[148][7] ), 
	.A2(n15), 
	.A1(n220));
   AO22CHD U4383 (.O(n2958), 
	.B2(n352), 
	.B1(\ram[148][8] ), 
	.A2(n16), 
	.A1(n220));
   AO22CHD U4384 (.O(n2959), 
	.B2(n352), 
	.B1(\ram[148][9] ), 
	.A2(n17), 
	.A1(n220));
   AO22CHD U4385 (.O(n2960), 
	.B2(n352), 
	.B1(\ram[148][10] ), 
	.A2(n18), 
	.A1(n220));
   AO22CHD U4386 (.O(n2961), 
	.B2(n352), 
	.B1(\ram[148][11] ), 
	.A2(n19), 
	.A1(n220));
   AO22CHD U4387 (.O(n2962), 
	.B2(n352), 
	.B1(\ram[148][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n220));
   AO22CHD U4388 (.O(n2963), 
	.B2(n352), 
	.B1(\ram[148][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n220));
   AO22CHD U4389 (.O(n2964), 
	.B2(n352), 
	.B1(\ram[148][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n220));
   AO22CHD U4390 (.O(n2965), 
	.B2(n352), 
	.B1(\ram[148][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n220));
   AO22CHD U4391 (.O(n2966), 
	.B2(n354), 
	.B1(\ram[149][0] ), 
	.A2(n6), 
	.A1(n222));
   AO22CHD U4392 (.O(n2967), 
	.B2(n354), 
	.B1(\ram[149][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n222));
   AO22CHD U4393 (.O(n2968), 
	.B2(n354), 
	.B1(\ram[149][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n222));
   AO22CHD U4394 (.O(n2969), 
	.B2(n354), 
	.B1(\ram[149][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n222));
   AO22CHD U4395 (.O(n2970), 
	.B2(n354), 
	.B1(\ram[149][4] ), 
	.A2(n12), 
	.A1(n222));
   AO22CHD U4396 (.O(n2971), 
	.B2(n354), 
	.B1(\ram[149][5] ), 
	.A2(n13), 
	.A1(n222));
   AO22CHD U4397 (.O(n2972), 
	.B2(n354), 
	.B1(\ram[149][6] ), 
	.A2(n14), 
	.A1(n222));
   AO22CHD U4398 (.O(n2973), 
	.B2(n354), 
	.B1(\ram[149][7] ), 
	.A2(n15), 
	.A1(n222));
   AO22CHD U4399 (.O(n2974), 
	.B2(n354), 
	.B1(\ram[149][8] ), 
	.A2(n16), 
	.A1(n222));
   AO22CHD U4400 (.O(n2975), 
	.B2(n354), 
	.B1(\ram[149][9] ), 
	.A2(n17), 
	.A1(n222));
   AO22CHD U4401 (.O(n2976), 
	.B2(n354), 
	.B1(\ram[149][10] ), 
	.A2(n18), 
	.A1(n222));
   AO22CHD U4402 (.O(n2977), 
	.B2(n354), 
	.B1(\ram[149][11] ), 
	.A2(n19), 
	.A1(n222));
   AO22CHD U4403 (.O(n2978), 
	.B2(n354), 
	.B1(\ram[149][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n222));
   AO22CHD U4404 (.O(n2979), 
	.B2(n354), 
	.B1(\ram[149][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n222));
   AO22CHD U4405 (.O(n2980), 
	.B2(n354), 
	.B1(\ram[149][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n222));
   AO22CHD U4406 (.O(n2981), 
	.B2(n354), 
	.B1(\ram[149][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n222));
   AO22CHD U4407 (.O(n2982), 
	.B2(n356), 
	.B1(\ram[150][0] ), 
	.A2(n6), 
	.A1(n224));
   AO22CHD U4408 (.O(n2983), 
	.B2(n356), 
	.B1(\ram[150][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n224));
   AO22CHD U4409 (.O(n2984), 
	.B2(n356), 
	.B1(\ram[150][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n224));
   AO22CHD U4410 (.O(n2985), 
	.B2(n356), 
	.B1(\ram[150][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n224));
   AO22CHD U4411 (.O(n2986), 
	.B2(n356), 
	.B1(\ram[150][4] ), 
	.A2(n12), 
	.A1(n224));
   AO22CHD U4412 (.O(n2987), 
	.B2(n356), 
	.B1(\ram[150][5] ), 
	.A2(n13), 
	.A1(n224));
   AO22CHD U4413 (.O(n2988), 
	.B2(n356), 
	.B1(\ram[150][6] ), 
	.A2(n14), 
	.A1(n224));
   AO22CHD U4414 (.O(n2989), 
	.B2(n356), 
	.B1(\ram[150][7] ), 
	.A2(n15), 
	.A1(n224));
   AO22CHD U4415 (.O(n2990), 
	.B2(n356), 
	.B1(\ram[150][8] ), 
	.A2(n16), 
	.A1(n224));
   AO22CHD U4416 (.O(n2991), 
	.B2(n356), 
	.B1(\ram[150][9] ), 
	.A2(n17), 
	.A1(n224));
   AO22CHD U4417 (.O(n2992), 
	.B2(n356), 
	.B1(\ram[150][10] ), 
	.A2(n18), 
	.A1(n224));
   AO22CHD U4418 (.O(n2993), 
	.B2(n356), 
	.B1(\ram[150][11] ), 
	.A2(n19), 
	.A1(n224));
   AO22CHD U4419 (.O(n2994), 
	.B2(n356), 
	.B1(\ram[150][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n224));
   AO22CHD U4420 (.O(n2995), 
	.B2(n356), 
	.B1(\ram[150][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n224));
   AO22CHD U4421 (.O(n2996), 
	.B2(n356), 
	.B1(\ram[150][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n224));
   AO22CHD U4422 (.O(n2997), 
	.B2(n356), 
	.B1(\ram[150][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n224));
   AO22CHD U4423 (.O(n2998), 
	.B2(n358), 
	.B1(\ram[151][0] ), 
	.A2(n6), 
	.A1(n226));
   AO22CHD U4424 (.O(n2999), 
	.B2(n358), 
	.B1(\ram[151][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n226));
   AO22CHD U4425 (.O(n3000), 
	.B2(n358), 
	.B1(\ram[151][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n226));
   AO22CHD U4426 (.O(n3001), 
	.B2(n358), 
	.B1(\ram[151][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n226));
   AO22CHD U4427 (.O(n3002), 
	.B2(n358), 
	.B1(\ram[151][4] ), 
	.A2(n12), 
	.A1(n226));
   AO22CHD U4428 (.O(n3003), 
	.B2(n358), 
	.B1(\ram[151][5] ), 
	.A2(n13), 
	.A1(n226));
   AO22CHD U4429 (.O(n3004), 
	.B2(n358), 
	.B1(\ram[151][6] ), 
	.A2(n14), 
	.A1(n226));
   AO22CHD U4430 (.O(n3005), 
	.B2(n358), 
	.B1(\ram[151][7] ), 
	.A2(n15), 
	.A1(n226));
   AO22CHD U4431 (.O(n3006), 
	.B2(n358), 
	.B1(\ram[151][8] ), 
	.A2(n16), 
	.A1(n226));
   AO22CHD U4432 (.O(n3007), 
	.B2(n358), 
	.B1(\ram[151][9] ), 
	.A2(n17), 
	.A1(n226));
   AO22CHD U4433 (.O(n3008), 
	.B2(n358), 
	.B1(\ram[151][10] ), 
	.A2(n18), 
	.A1(n226));
   AO22CHD U4434 (.O(n3009), 
	.B2(n358), 
	.B1(\ram[151][11] ), 
	.A2(n19), 
	.A1(n226));
   AO22CHD U4435 (.O(n3010), 
	.B2(n358), 
	.B1(\ram[151][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n226));
   AO22CHD U4436 (.O(n3011), 
	.B2(n358), 
	.B1(\ram[151][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n226));
   AO22CHD U4437 (.O(n3012), 
	.B2(n358), 
	.B1(\ram[151][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n226));
   AO22CHD U4438 (.O(n3013), 
	.B2(n358), 
	.B1(\ram[151][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n226));
   AO22CHD U4439 (.O(n3014), 
	.B2(n360), 
	.B1(\ram[152][0] ), 
	.A2(n6), 
	.A1(n228));
   AO22CHD U4440 (.O(n3015), 
	.B2(n360), 
	.B1(\ram[152][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n228));
   AO22CHD U4441 (.O(n3016), 
	.B2(n360), 
	.B1(\ram[152][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n228));
   AO22CHD U4442 (.O(n3017), 
	.B2(n360), 
	.B1(\ram[152][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n228));
   AO22CHD U4443 (.O(n3018), 
	.B2(n360), 
	.B1(\ram[152][4] ), 
	.A2(n12), 
	.A1(n228));
   AO22CHD U4444 (.O(n3019), 
	.B2(n360), 
	.B1(\ram[152][5] ), 
	.A2(n13), 
	.A1(n228));
   AO22CHD U4445 (.O(n3020), 
	.B2(n360), 
	.B1(\ram[152][6] ), 
	.A2(n14), 
	.A1(n228));
   AO22CHD U4446 (.O(n3021), 
	.B2(n360), 
	.B1(\ram[152][7] ), 
	.A2(n15), 
	.A1(n228));
   AO22CHD U4447 (.O(n3022), 
	.B2(n360), 
	.B1(\ram[152][8] ), 
	.A2(n16), 
	.A1(n228));
   AO22CHD U4448 (.O(n3023), 
	.B2(n360), 
	.B1(\ram[152][9] ), 
	.A2(n17), 
	.A1(n228));
   AO22CHD U4449 (.O(n3024), 
	.B2(n360), 
	.B1(\ram[152][10] ), 
	.A2(n18), 
	.A1(n228));
   AO22CHD U4450 (.O(n3025), 
	.B2(n360), 
	.B1(\ram[152][11] ), 
	.A2(n19), 
	.A1(n228));
   AO22CHD U4451 (.O(n3026), 
	.B2(n360), 
	.B1(\ram[152][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n228));
   AO22CHD U4452 (.O(n3027), 
	.B2(n360), 
	.B1(\ram[152][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n228));
   AO22CHD U4453 (.O(n3028), 
	.B2(n360), 
	.B1(\ram[152][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n228));
   AO22CHD U4454 (.O(n3029), 
	.B2(n360), 
	.B1(\ram[152][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n228));
   AO22CHD U4455 (.O(n3030), 
	.B2(n362), 
	.B1(\ram[153][0] ), 
	.A2(n6), 
	.A1(n230));
   AO22CHD U4456 (.O(n3031), 
	.B2(n362), 
	.B1(\ram[153][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n230));
   AO22CHD U4457 (.O(n3032), 
	.B2(n362), 
	.B1(\ram[153][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n230));
   AO22CHD U4458 (.O(n3033), 
	.B2(n362), 
	.B1(\ram[153][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n230));
   AO22CHD U4459 (.O(n3034), 
	.B2(n362), 
	.B1(\ram[153][4] ), 
	.A2(n12), 
	.A1(n230));
   AO22CHD U4460 (.O(n3035), 
	.B2(n362), 
	.B1(\ram[153][5] ), 
	.A2(n13), 
	.A1(n230));
   AO22CHD U4461 (.O(n3036), 
	.B2(n362), 
	.B1(\ram[153][6] ), 
	.A2(n14), 
	.A1(n230));
   AO22CHD U4462 (.O(n3037), 
	.B2(n362), 
	.B1(\ram[153][7] ), 
	.A2(n15), 
	.A1(n230));
   AO22CHD U4463 (.O(n3038), 
	.B2(n362), 
	.B1(\ram[153][8] ), 
	.A2(n16), 
	.A1(n230));
   AO22CHD U4464 (.O(n3039), 
	.B2(n362), 
	.B1(\ram[153][9] ), 
	.A2(n17), 
	.A1(n230));
   AO22CHD U4465 (.O(n3040), 
	.B2(n362), 
	.B1(\ram[153][10] ), 
	.A2(n18), 
	.A1(n230));
   AO22CHD U4466 (.O(n3041), 
	.B2(n362), 
	.B1(\ram[153][11] ), 
	.A2(n19), 
	.A1(n230));
   AO22CHD U4467 (.O(n3042), 
	.B2(n362), 
	.B1(\ram[153][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n230));
   AO22CHD U4468 (.O(n3043), 
	.B2(n362), 
	.B1(\ram[153][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n230));
   AO22CHD U4469 (.O(n3044), 
	.B2(n362), 
	.B1(\ram[153][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n230));
   AO22CHD U4470 (.O(n3045), 
	.B2(n362), 
	.B1(\ram[153][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n230));
   AO22CHD U4471 (.O(n3046), 
	.B2(n364), 
	.B1(\ram[154][0] ), 
	.A2(n6), 
	.A1(n232));
   AO22CHD U4472 (.O(n3047), 
	.B2(n364), 
	.B1(\ram[154][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n232));
   AO22CHD U4473 (.O(n3048), 
	.B2(n364), 
	.B1(\ram[154][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n232));
   AO22CHD U4474 (.O(n3049), 
	.B2(n364), 
	.B1(\ram[154][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n232));
   AO22CHD U4475 (.O(n3050), 
	.B2(n364), 
	.B1(\ram[154][4] ), 
	.A2(n12), 
	.A1(n232));
   AO22CHD U4476 (.O(n3051), 
	.B2(n364), 
	.B1(\ram[154][5] ), 
	.A2(n13), 
	.A1(n232));
   AO22CHD U4477 (.O(n3052), 
	.B2(n364), 
	.B1(\ram[154][6] ), 
	.A2(n14), 
	.A1(n232));
   AO22CHD U4478 (.O(n3053), 
	.B2(n364), 
	.B1(\ram[154][7] ), 
	.A2(n15), 
	.A1(n232));
   AO22CHD U4479 (.O(n3054), 
	.B2(n364), 
	.B1(\ram[154][8] ), 
	.A2(n16), 
	.A1(n232));
   AO22CHD U4480 (.O(n3055), 
	.B2(n364), 
	.B1(\ram[154][9] ), 
	.A2(n17), 
	.A1(n232));
   AO22CHD U4481 (.O(n3056), 
	.B2(n364), 
	.B1(\ram[154][10] ), 
	.A2(n18), 
	.A1(n232));
   AO22CHD U4482 (.O(n3057), 
	.B2(n364), 
	.B1(\ram[154][11] ), 
	.A2(n19), 
	.A1(n232));
   AO22CHD U4483 (.O(n3058), 
	.B2(n364), 
	.B1(\ram[154][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n232));
   AO22CHD U4484 (.O(n3059), 
	.B2(n364), 
	.B1(\ram[154][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n232));
   AO22CHD U4485 (.O(n3060), 
	.B2(n364), 
	.B1(\ram[154][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n232));
   AO22CHD U4486 (.O(n3061), 
	.B2(n364), 
	.B1(\ram[154][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n232));
   AO22CHD U4487 (.O(n3062), 
	.B2(n366), 
	.B1(\ram[155][0] ), 
	.A2(n6), 
	.A1(n234));
   AO22CHD U4488 (.O(n3063), 
	.B2(n366), 
	.B1(\ram[155][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n234));
   AO22CHD U4489 (.O(n3064), 
	.B2(n366), 
	.B1(\ram[155][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n234));
   AO22CHD U4490 (.O(n3065), 
	.B2(n366), 
	.B1(\ram[155][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n234));
   AO22CHD U4491 (.O(n3066), 
	.B2(n366), 
	.B1(\ram[155][4] ), 
	.A2(n12), 
	.A1(n234));
   AO22CHD U4492 (.O(n3067), 
	.B2(n366), 
	.B1(\ram[155][5] ), 
	.A2(n13), 
	.A1(n234));
   AO22CHD U4493 (.O(n3068), 
	.B2(n366), 
	.B1(\ram[155][6] ), 
	.A2(n14), 
	.A1(n234));
   AO22CHD U4494 (.O(n3069), 
	.B2(n366), 
	.B1(\ram[155][7] ), 
	.A2(n15), 
	.A1(n234));
   AO22CHD U4495 (.O(n3070), 
	.B2(n366), 
	.B1(\ram[155][8] ), 
	.A2(n16), 
	.A1(n234));
   AO22CHD U4496 (.O(n3071), 
	.B2(n366), 
	.B1(\ram[155][9] ), 
	.A2(n17), 
	.A1(n234));
   AO22CHD U4497 (.O(n3072), 
	.B2(n366), 
	.B1(\ram[155][10] ), 
	.A2(n18), 
	.A1(n234));
   AO22CHD U4498 (.O(n3073), 
	.B2(n366), 
	.B1(\ram[155][11] ), 
	.A2(n19), 
	.A1(n234));
   AO22CHD U4499 (.O(n3074), 
	.B2(n366), 
	.B1(\ram[155][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n234));
   AO22CHD U4500 (.O(n3075), 
	.B2(n366), 
	.B1(\ram[155][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n234));
   AO22CHD U4501 (.O(n3076), 
	.B2(n366), 
	.B1(\ram[155][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n234));
   AO22CHD U4502 (.O(n3077), 
	.B2(n366), 
	.B1(\ram[155][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n234));
   AO22CHD U4503 (.O(n3078), 
	.B2(n368), 
	.B1(\ram[156][0] ), 
	.A2(n6), 
	.A1(n236));
   AO22CHD U4504 (.O(n3079), 
	.B2(n368), 
	.B1(\ram[156][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n236));
   AO22CHD U4505 (.O(n3080), 
	.B2(n368), 
	.B1(\ram[156][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n236));
   AO22CHD U4506 (.O(n3081), 
	.B2(n368), 
	.B1(\ram[156][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n236));
   AO22CHD U4507 (.O(n3082), 
	.B2(n368), 
	.B1(\ram[156][4] ), 
	.A2(n12), 
	.A1(n236));
   AO22CHD U4508 (.O(n3083), 
	.B2(n368), 
	.B1(\ram[156][5] ), 
	.A2(n13), 
	.A1(n236));
   AO22CHD U4509 (.O(n3084), 
	.B2(n368), 
	.B1(\ram[156][6] ), 
	.A2(n14), 
	.A1(n236));
   AO22CHD U4510 (.O(n3085), 
	.B2(n368), 
	.B1(\ram[156][7] ), 
	.A2(n15), 
	.A1(n236));
   AO22CHD U4511 (.O(n3086), 
	.B2(n368), 
	.B1(\ram[156][8] ), 
	.A2(n16), 
	.A1(n236));
   AO22CHD U4512 (.O(n3087), 
	.B2(n368), 
	.B1(\ram[156][9] ), 
	.A2(n17), 
	.A1(n236));
   AO22CHD U4513 (.O(n3088), 
	.B2(n368), 
	.B1(\ram[156][10] ), 
	.A2(n18), 
	.A1(n236));
   AO22CHD U4514 (.O(n3089), 
	.B2(n368), 
	.B1(\ram[156][11] ), 
	.A2(n19), 
	.A1(n236));
   AO22CHD U4515 (.O(n3090), 
	.B2(n368), 
	.B1(\ram[156][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n236));
   AO22CHD U4516 (.O(n3091), 
	.B2(n368), 
	.B1(\ram[156][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n236));
   AO22CHD U4517 (.O(n3092), 
	.B2(n368), 
	.B1(\ram[156][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n236));
   AO22CHD U4518 (.O(n3093), 
	.B2(n368), 
	.B1(\ram[156][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n236));
   AO22CHD U4519 (.O(n3094), 
	.B2(n370), 
	.B1(\ram[157][0] ), 
	.A2(n6), 
	.A1(n238));
   AO22CHD U4520 (.O(n3095), 
	.B2(n370), 
	.B1(\ram[157][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n238));
   AO22CHD U4521 (.O(n3096), 
	.B2(n370), 
	.B1(\ram[157][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n238));
   AO22CHD U4522 (.O(n3097), 
	.B2(n370), 
	.B1(\ram[157][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n238));
   AO22CHD U4523 (.O(n3098), 
	.B2(n370), 
	.B1(\ram[157][4] ), 
	.A2(n12), 
	.A1(n238));
   AO22CHD U4524 (.O(n3099), 
	.B2(n370), 
	.B1(\ram[157][5] ), 
	.A2(n13), 
	.A1(n238));
   AO22CHD U4525 (.O(n3100), 
	.B2(n370), 
	.B1(\ram[157][6] ), 
	.A2(n14), 
	.A1(n238));
   AO22CHD U4526 (.O(n3101), 
	.B2(n370), 
	.B1(\ram[157][7] ), 
	.A2(n15), 
	.A1(n238));
   AO22CHD U4527 (.O(n3102), 
	.B2(n370), 
	.B1(\ram[157][8] ), 
	.A2(n16), 
	.A1(n238));
   AO22CHD U4528 (.O(n3103), 
	.B2(n370), 
	.B1(\ram[157][9] ), 
	.A2(n17), 
	.A1(n238));
   AO22CHD U4529 (.O(n3104), 
	.B2(n370), 
	.B1(\ram[157][10] ), 
	.A2(n18), 
	.A1(n238));
   AO22CHD U4530 (.O(n3105), 
	.B2(n370), 
	.B1(\ram[157][11] ), 
	.A2(n19), 
	.A1(n238));
   AO22CHD U4531 (.O(n3106), 
	.B2(n370), 
	.B1(\ram[157][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n238));
   AO22CHD U4532 (.O(n3107), 
	.B2(n370), 
	.B1(\ram[157][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n238));
   AO22CHD U4533 (.O(n3108), 
	.B2(n370), 
	.B1(\ram[157][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n238));
   AO22CHD U4534 (.O(n3109), 
	.B2(n370), 
	.B1(\ram[157][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n238));
   AO22CHD U4535 (.O(n3110), 
	.B2(n372), 
	.B1(\ram[158][0] ), 
	.A2(n6), 
	.A1(n240));
   AO22CHD U4536 (.O(n3111), 
	.B2(n372), 
	.B1(\ram[158][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n240));
   AO22CHD U4537 (.O(n3112), 
	.B2(n372), 
	.B1(\ram[158][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n240));
   AO22CHD U4538 (.O(n3113), 
	.B2(n372), 
	.B1(\ram[158][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n240));
   AO22CHD U4539 (.O(n3114), 
	.B2(n372), 
	.B1(\ram[158][4] ), 
	.A2(n12), 
	.A1(n240));
   AO22CHD U4540 (.O(n3115), 
	.B2(n372), 
	.B1(\ram[158][5] ), 
	.A2(n13), 
	.A1(n240));
   AO22CHD U4541 (.O(n3116), 
	.B2(n372), 
	.B1(\ram[158][6] ), 
	.A2(n14), 
	.A1(n240));
   AO22CHD U4542 (.O(n3117), 
	.B2(n372), 
	.B1(\ram[158][7] ), 
	.A2(n15), 
	.A1(n240));
   AO22CHD U4543 (.O(n3118), 
	.B2(n372), 
	.B1(\ram[158][8] ), 
	.A2(n16), 
	.A1(n240));
   AO22CHD U4544 (.O(n3119), 
	.B2(n372), 
	.B1(\ram[158][9] ), 
	.A2(n17), 
	.A1(n240));
   AO22CHD U4545 (.O(n3120), 
	.B2(n372), 
	.B1(\ram[158][10] ), 
	.A2(n18), 
	.A1(n240));
   AO22CHD U4546 (.O(n3121), 
	.B2(n372), 
	.B1(\ram[158][11] ), 
	.A2(n19), 
	.A1(n240));
   AO22CHD U4547 (.O(n3122), 
	.B2(n372), 
	.B1(\ram[158][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n240));
   AO22CHD U4548 (.O(n3123), 
	.B2(n372), 
	.B1(\ram[158][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n240));
   AO22CHD U4549 (.O(n3124), 
	.B2(n372), 
	.B1(\ram[158][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n240));
   AO22CHD U4550 (.O(n3125), 
	.B2(n372), 
	.B1(\ram[158][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n240));
   AO22CHD U4551 (.O(n3126), 
	.B2(n374), 
	.B1(\ram[159][0] ), 
	.A2(n6), 
	.A1(n242));
   AO22CHD U4552 (.O(n3127), 
	.B2(n374), 
	.B1(\ram[159][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n242));
   AO22CHD U4553 (.O(n3128), 
	.B2(n374), 
	.B1(\ram[159][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n242));
   AO22CHD U4554 (.O(n3129), 
	.B2(n374), 
	.B1(\ram[159][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n242));
   AO22CHD U4555 (.O(n3130), 
	.B2(n374), 
	.B1(\ram[159][4] ), 
	.A2(n12), 
	.A1(n242));
   AO22CHD U4556 (.O(n3131), 
	.B2(n374), 
	.B1(\ram[159][5] ), 
	.A2(n13), 
	.A1(n242));
   AO22CHD U4557 (.O(n3132), 
	.B2(n374), 
	.B1(\ram[159][6] ), 
	.A2(n14), 
	.A1(n242));
   AO22CHD U4558 (.O(n3133), 
	.B2(n374), 
	.B1(\ram[159][7] ), 
	.A2(n15), 
	.A1(n242));
   AO22CHD U4559 (.O(n3134), 
	.B2(n374), 
	.B1(\ram[159][8] ), 
	.A2(n16), 
	.A1(n242));
   AO22CHD U4560 (.O(n3135), 
	.B2(n374), 
	.B1(\ram[159][9] ), 
	.A2(n17), 
	.A1(n242));
   AO22CHD U4561 (.O(n3136), 
	.B2(n374), 
	.B1(\ram[159][10] ), 
	.A2(n18), 
	.A1(n242));
   AO22CHD U4562 (.O(n3137), 
	.B2(n374), 
	.B1(\ram[159][11] ), 
	.A2(n19), 
	.A1(n242));
   AO22CHD U4563 (.O(n3138), 
	.B2(n374), 
	.B1(\ram[159][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n242));
   AO22CHD U4564 (.O(n3139), 
	.B2(n374), 
	.B1(\ram[159][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n242));
   AO22CHD U4565 (.O(n3140), 
	.B2(n374), 
	.B1(\ram[159][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n242));
   AO22CHD U4566 (.O(n3141), 
	.B2(n374), 
	.B1(\ram[159][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n242));
   AO22CHD U4567 (.O(n3142), 
	.B2(n376), 
	.B1(\ram[160][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n244));
   AO22CHD U4568 (.O(n3143), 
	.B2(n376), 
	.B1(\ram[160][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n244));
   AO22CHD U4569 (.O(n3144), 
	.B2(n376), 
	.B1(\ram[160][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n244));
   AO22CHD U4570 (.O(n3145), 
	.B2(n376), 
	.B1(\ram[160][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n244));
   AO22CHD U4571 (.O(n3146), 
	.B2(n376), 
	.B1(\ram[160][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n244));
   AO22CHD U4572 (.O(n3147), 
	.B2(n376), 
	.B1(\ram[160][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n244));
   AO22CHD U4573 (.O(n3148), 
	.B2(n376), 
	.B1(\ram[160][6] ), 
	.A2(n14), 
	.A1(n244));
   AO22CHD U4574 (.O(n3149), 
	.B2(n376), 
	.B1(\ram[160][7] ), 
	.A2(n15), 
	.A1(n244));
   AO22CHD U4575 (.O(n3150), 
	.B2(n376), 
	.B1(\ram[160][8] ), 
	.A2(n16), 
	.A1(n244));
   AO22CHD U4576 (.O(n3151), 
	.B2(n376), 
	.B1(\ram[160][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n244));
   AO22CHD U4577 (.O(n3152), 
	.B2(n376), 
	.B1(\ram[160][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n244));
   AO22CHD U4578 (.O(n3153), 
	.B2(n376), 
	.B1(\ram[160][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n244));
   AO22CHD U4579 (.O(n3154), 
	.B2(n376), 
	.B1(\ram[160][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n244));
   AO22CHD U4580 (.O(n3155), 
	.B2(n376), 
	.B1(\ram[160][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n244));
   AO22CHD U4581 (.O(n3156), 
	.B2(n376), 
	.B1(\ram[160][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n244));
   AO22CHD U4582 (.O(n3157), 
	.B2(n376), 
	.B1(\ram[160][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n244));
   AO22CHD U4583 (.O(n3158), 
	.B2(n379), 
	.B1(\ram[161][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n245));
   AO22CHD U4584 (.O(n3159), 
	.B2(n379), 
	.B1(\ram[161][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n245));
   AO22CHD U4585 (.O(n3160), 
	.B2(n379), 
	.B1(\ram[161][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n245));
   AO22CHD U4586 (.O(n3161), 
	.B2(n379), 
	.B1(\ram[161][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n245));
   AO22CHD U4587 (.O(n3162), 
	.B2(n379), 
	.B1(\ram[161][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n245));
   AO22CHD U4588 (.O(n3163), 
	.B2(n379), 
	.B1(\ram[161][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n245));
   AO22CHD U4589 (.O(n3164), 
	.B2(n379), 
	.B1(\ram[161][6] ), 
	.A2(n14), 
	.A1(n245));
   AO22CHD U4590 (.O(n3165), 
	.B2(n379), 
	.B1(\ram[161][7] ), 
	.A2(n15), 
	.A1(n245));
   AO22CHD U4591 (.O(n3166), 
	.B2(n379), 
	.B1(\ram[161][8] ), 
	.A2(n16), 
	.A1(n245));
   AO22CHD U4592 (.O(n3167), 
	.B2(n379), 
	.B1(\ram[161][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n245));
   AO22CHD U4593 (.O(n3168), 
	.B2(n379), 
	.B1(\ram[161][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n245));
   AO22CHD U4594 (.O(n3169), 
	.B2(n379), 
	.B1(\ram[161][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n245));
   AO22CHD U4595 (.O(n3170), 
	.B2(n379), 
	.B1(\ram[161][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n245));
   AO22CHD U4596 (.O(n3171), 
	.B2(n379), 
	.B1(\ram[161][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n245));
   AO22CHD U4597 (.O(n3172), 
	.B2(n379), 
	.B1(\ram[161][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n245));
   AO22CHD U4598 (.O(n3173), 
	.B2(n379), 
	.B1(\ram[161][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n245));
   AO22CHD U4599 (.O(n3174), 
	.B2(n381), 
	.B1(\ram[162][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n247));
   AO22CHD U4600 (.O(n3175), 
	.B2(n381), 
	.B1(\ram[162][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n247));
   AO22CHD U4601 (.O(n3176), 
	.B2(n381), 
	.B1(\ram[162][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n247));
   AO22CHD U4602 (.O(n3177), 
	.B2(n381), 
	.B1(\ram[162][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n247));
   AO22CHD U4603 (.O(n3178), 
	.B2(n381), 
	.B1(\ram[162][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n247));
   AO22CHD U4604 (.O(n3179), 
	.B2(n381), 
	.B1(\ram[162][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n247));
   AO22CHD U4605 (.O(n3180), 
	.B2(n381), 
	.B1(\ram[162][6] ), 
	.A2(n14), 
	.A1(n247));
   AO22CHD U4606 (.O(n3181), 
	.B2(n381), 
	.B1(\ram[162][7] ), 
	.A2(n15), 
	.A1(n247));
   AO22CHD U4607 (.O(n3182), 
	.B2(n381), 
	.B1(\ram[162][8] ), 
	.A2(n16), 
	.A1(n247));
   AO22CHD U4608 (.O(n3183), 
	.B2(n381), 
	.B1(\ram[162][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n247));
   AO22CHD U4609 (.O(n3184), 
	.B2(n381), 
	.B1(\ram[162][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n247));
   AO22CHD U4610 (.O(n3185), 
	.B2(n381), 
	.B1(\ram[162][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n247));
   AO22CHD U4611 (.O(n3186), 
	.B2(n381), 
	.B1(\ram[162][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n247));
   AO22CHD U4612 (.O(n3187), 
	.B2(n381), 
	.B1(\ram[162][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n247));
   AO22CHD U4613 (.O(n3188), 
	.B2(n381), 
	.B1(\ram[162][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n247));
   AO22CHD U4614 (.O(n3189), 
	.B2(n381), 
	.B1(\ram[162][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n247));
   AO22CHD U4615 (.O(n3190), 
	.B2(n383), 
	.B1(\ram[163][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n249));
   AO22CHD U4616 (.O(n3191), 
	.B2(n383), 
	.B1(\ram[163][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n249));
   AO22CHD U4617 (.O(n3192), 
	.B2(n383), 
	.B1(\ram[163][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n249));
   AO22CHD U4618 (.O(n3193), 
	.B2(n383), 
	.B1(\ram[163][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n249));
   AO22CHD U4619 (.O(n3194), 
	.B2(n383), 
	.B1(\ram[163][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n249));
   AO22CHD U4620 (.O(n3195), 
	.B2(n383), 
	.B1(\ram[163][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n249));
   AO22CHD U4621 (.O(n3196), 
	.B2(n383), 
	.B1(\ram[163][6] ), 
	.A2(n14), 
	.A1(n249));
   AO22CHD U4622 (.O(n3197), 
	.B2(n383), 
	.B1(\ram[163][7] ), 
	.A2(n15), 
	.A1(n249));
   AO22CHD U4623 (.O(n3198), 
	.B2(n383), 
	.B1(\ram[163][8] ), 
	.A2(n16), 
	.A1(n249));
   AO22CHD U4624 (.O(n3199), 
	.B2(n383), 
	.B1(\ram[163][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n249));
   AO22CHD U4625 (.O(n3200), 
	.B2(n383), 
	.B1(\ram[163][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n249));
   AO22CHD U4626 (.O(n3201), 
	.B2(n383), 
	.B1(\ram[163][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n249));
   AO22CHD U4627 (.O(n3202), 
	.B2(n383), 
	.B1(\ram[163][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n249));
   AO22CHD U4628 (.O(n3203), 
	.B2(n383), 
	.B1(\ram[163][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n249));
   AO22CHD U4629 (.O(n3204), 
	.B2(n383), 
	.B1(\ram[163][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n249));
   AO22CHD U4630 (.O(n3205), 
	.B2(n383), 
	.B1(\ram[163][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n249));
   AO22CHD U4631 (.O(n3206), 
	.B2(n385), 
	.B1(\ram[164][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n251));
   AO22CHD U4632 (.O(n3207), 
	.B2(n385), 
	.B1(\ram[164][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n251));
   AO22CHD U4633 (.O(n3208), 
	.B2(n385), 
	.B1(\ram[164][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n251));
   AO22CHD U4634 (.O(n3209), 
	.B2(n385), 
	.B1(\ram[164][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n251));
   AO22CHD U4635 (.O(n3210), 
	.B2(n385), 
	.B1(\ram[164][4] ), 
	.A2(n12), 
	.A1(n251));
   AO22CHD U4636 (.O(n3211), 
	.B2(n385), 
	.B1(\ram[164][5] ), 
	.A2(n13), 
	.A1(n251));
   AO22CHD U4637 (.O(n3212), 
	.B2(n385), 
	.B1(\ram[164][6] ), 
	.A2(n14), 
	.A1(n251));
   AO22CHD U4638 (.O(n3213), 
	.B2(n385), 
	.B1(\ram[164][7] ), 
	.A2(n15), 
	.A1(n251));
   AO22CHD U4639 (.O(n3214), 
	.B2(n385), 
	.B1(\ram[164][8] ), 
	.A2(n16), 
	.A1(n251));
   AO22CHD U4640 (.O(n3215), 
	.B2(n385), 
	.B1(\ram[164][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n251));
   AO22CHD U4641 (.O(n3216), 
	.B2(n385), 
	.B1(\ram[164][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n251));
   AO22CHD U4642 (.O(n3217), 
	.B2(n385), 
	.B1(\ram[164][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n251));
   AO22CHD U4643 (.O(n3218), 
	.B2(n385), 
	.B1(\ram[164][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n251));
   AO22CHD U4644 (.O(n3219), 
	.B2(n385), 
	.B1(\ram[164][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n251));
   AO22CHD U4645 (.O(n3220), 
	.B2(n385), 
	.B1(\ram[164][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n251));
   AO22CHD U4646 (.O(n3221), 
	.B2(n385), 
	.B1(\ram[164][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n251));
   AO22CHD U4647 (.O(n3222), 
	.B2(n387), 
	.B1(\ram[165][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n253));
   AO22CHD U4648 (.O(n3223), 
	.B2(n387), 
	.B1(\ram[165][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n253));
   AO22CHD U4649 (.O(n3224), 
	.B2(n387), 
	.B1(\ram[165][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n253));
   AO22CHD U4650 (.O(n3225), 
	.B2(n387), 
	.B1(\ram[165][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n253));
   AO22CHD U4651 (.O(n3226), 
	.B2(n387), 
	.B1(\ram[165][4] ), 
	.A2(n12), 
	.A1(n253));
   AO22CHD U4652 (.O(n3227), 
	.B2(n387), 
	.B1(\ram[165][5] ), 
	.A2(n13), 
	.A1(n253));
   AO22CHD U4653 (.O(n3228), 
	.B2(n387), 
	.B1(\ram[165][6] ), 
	.A2(n14), 
	.A1(n253));
   AO22CHD U4654 (.O(n3229), 
	.B2(n387), 
	.B1(\ram[165][7] ), 
	.A2(n15), 
	.A1(n253));
   AO22CHD U4655 (.O(n3230), 
	.B2(n387), 
	.B1(\ram[165][8] ), 
	.A2(n16), 
	.A1(n253));
   AO22CHD U4656 (.O(n3231), 
	.B2(n387), 
	.B1(\ram[165][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n253));
   AO22CHD U4657 (.O(n3232), 
	.B2(n387), 
	.B1(\ram[165][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n253));
   AO22CHD U4658 (.O(n3233), 
	.B2(n387), 
	.B1(\ram[165][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n253));
   AO22CHD U4659 (.O(n3234), 
	.B2(n387), 
	.B1(\ram[165][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n253));
   AO22CHD U4660 (.O(n3235), 
	.B2(n387), 
	.B1(\ram[165][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n253));
   AO22CHD U4661 (.O(n3236), 
	.B2(n387), 
	.B1(\ram[165][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n253));
   AO22CHD U4662 (.O(n3237), 
	.B2(n387), 
	.B1(\ram[165][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n253));
   AO22CHD U4663 (.O(n3238), 
	.B2(n389), 
	.B1(\ram[166][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n255));
   AO22CHD U4664 (.O(n3239), 
	.B2(n389), 
	.B1(\ram[166][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n255));
   AO22CHD U4665 (.O(n3240), 
	.B2(n389), 
	.B1(\ram[166][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n255));
   AO22CHD U4666 (.O(n3241), 
	.B2(n389), 
	.B1(\ram[166][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n255));
   AO22CHD U4667 (.O(n3242), 
	.B2(n389), 
	.B1(\ram[166][4] ), 
	.A2(n12), 
	.A1(n255));
   AO22CHD U4668 (.O(n3243), 
	.B2(n389), 
	.B1(\ram[166][5] ), 
	.A2(n13), 
	.A1(n255));
   AO22CHD U4669 (.O(n3244), 
	.B2(n389), 
	.B1(\ram[166][6] ), 
	.A2(n14), 
	.A1(n255));
   AO22CHD U4670 (.O(n3245), 
	.B2(n389), 
	.B1(\ram[166][7] ), 
	.A2(n15), 
	.A1(n255));
   AO22CHD U4671 (.O(n3246), 
	.B2(n389), 
	.B1(\ram[166][8] ), 
	.A2(n16), 
	.A1(n255));
   AO22CHD U4672 (.O(n3247), 
	.B2(n389), 
	.B1(\ram[166][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n255));
   AO22CHD U4673 (.O(n3248), 
	.B2(n389), 
	.B1(\ram[166][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n255));
   AO22CHD U4674 (.O(n3249), 
	.B2(n389), 
	.B1(\ram[166][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n255));
   AO22CHD U4675 (.O(n3250), 
	.B2(n389), 
	.B1(\ram[166][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n255));
   AO22CHD U4676 (.O(n3251), 
	.B2(n389), 
	.B1(\ram[166][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n255));
   AO22CHD U4677 (.O(n3252), 
	.B2(n389), 
	.B1(\ram[166][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n255));
   AO22CHD U4678 (.O(n3253), 
	.B2(n389), 
	.B1(\ram[166][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n255));
   AO22CHD U4679 (.O(n3254), 
	.B2(n391), 
	.B1(\ram[167][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n257));
   AO22CHD U4680 (.O(n3255), 
	.B2(n391), 
	.B1(\ram[167][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n257));
   AO22CHD U4681 (.O(n3256), 
	.B2(n391), 
	.B1(\ram[167][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n257));
   AO22CHD U4682 (.O(n3257), 
	.B2(n391), 
	.B1(\ram[167][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n257));
   AO22CHD U4683 (.O(n3258), 
	.B2(n391), 
	.B1(\ram[167][4] ), 
	.A2(n12), 
	.A1(n257));
   AO22CHD U4684 (.O(n3259), 
	.B2(n391), 
	.B1(\ram[167][5] ), 
	.A2(n13), 
	.A1(n257));
   AO22CHD U4685 (.O(n3260), 
	.B2(n391), 
	.B1(\ram[167][6] ), 
	.A2(n14), 
	.A1(n257));
   AO22CHD U4686 (.O(n3261), 
	.B2(n391), 
	.B1(\ram[167][7] ), 
	.A2(n15), 
	.A1(n257));
   AO22CHD U4687 (.O(n3262), 
	.B2(n391), 
	.B1(\ram[167][8] ), 
	.A2(n16), 
	.A1(n257));
   AO22CHD U4688 (.O(n3263), 
	.B2(n391), 
	.B1(\ram[167][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n257));
   AO22CHD U4689 (.O(n3264), 
	.B2(n391), 
	.B1(\ram[167][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n257));
   AO22CHD U4690 (.O(n3265), 
	.B2(n391), 
	.B1(\ram[167][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n257));
   AO22CHD U4691 (.O(n3266), 
	.B2(n391), 
	.B1(\ram[167][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n257));
   AO22CHD U4692 (.O(n3267), 
	.B2(n391), 
	.B1(\ram[167][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n257));
   AO22CHD U4693 (.O(n3268), 
	.B2(n391), 
	.B1(\ram[167][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n257));
   AO22CHD U4694 (.O(n3269), 
	.B2(n391), 
	.B1(\ram[167][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n257));
   AO22CHD U4695 (.O(n3270), 
	.B2(n393), 
	.B1(\ram[168][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n259));
   AO22CHD U4696 (.O(n3271), 
	.B2(n393), 
	.B1(\ram[168][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n259));
   AO22CHD U4697 (.O(n3272), 
	.B2(n393), 
	.B1(\ram[168][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n259));
   AO22CHD U4698 (.O(n3273), 
	.B2(n393), 
	.B1(\ram[168][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n259));
   AO22CHD U4699 (.O(n3274), 
	.B2(n393), 
	.B1(\ram[168][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n259));
   AO22CHD U4700 (.O(n3275), 
	.B2(n393), 
	.B1(\ram[168][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n259));
   AO22CHD U4701 (.O(n3276), 
	.B2(n393), 
	.B1(\ram[168][6] ), 
	.A2(n14), 
	.A1(n259));
   AO22CHD U4702 (.O(n3277), 
	.B2(n393), 
	.B1(\ram[168][7] ), 
	.A2(n15), 
	.A1(n259));
   AO22CHD U4703 (.O(n3278), 
	.B2(n393), 
	.B1(\ram[168][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n259));
   AO22CHD U4704 (.O(n3279), 
	.B2(n393), 
	.B1(\ram[168][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n259));
   AO22CHD U4705 (.O(n3280), 
	.B2(n393), 
	.B1(\ram[168][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n259));
   AO22CHD U4706 (.O(n3281), 
	.B2(n393), 
	.B1(\ram[168][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n259));
   AO22CHD U4707 (.O(n3282), 
	.B2(n393), 
	.B1(\ram[168][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n259));
   AO22CHD U4708 (.O(n3283), 
	.B2(n393), 
	.B1(\ram[168][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n259));
   AO22CHD U4709 (.O(n3284), 
	.B2(n393), 
	.B1(\ram[168][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n259));
   AO22CHD U4710 (.O(n3285), 
	.B2(n393), 
	.B1(\ram[168][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n259));
   AO22CHD U4711 (.O(n3286), 
	.B2(n395), 
	.B1(\ram[169][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n261));
   AO22CHD U4712 (.O(n3287), 
	.B2(n395), 
	.B1(\ram[169][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n261));
   AO22CHD U4713 (.O(n3288), 
	.B2(n395), 
	.B1(\ram[169][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n261));
   AO22CHD U4714 (.O(n3289), 
	.B2(n395), 
	.B1(\ram[169][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n261));
   AO22CHD U4715 (.O(n3290), 
	.B2(n395), 
	.B1(\ram[169][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n261));
   AO22CHD U4716 (.O(n3291), 
	.B2(n395), 
	.B1(\ram[169][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n261));
   AO22CHD U4717 (.O(n3292), 
	.B2(n395), 
	.B1(\ram[169][6] ), 
	.A2(n14), 
	.A1(n261));
   AO22CHD U4718 (.O(n3293), 
	.B2(n395), 
	.B1(\ram[169][7] ), 
	.A2(n15), 
	.A1(n261));
   AO22CHD U4719 (.O(n3294), 
	.B2(n395), 
	.B1(\ram[169][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n261));
   AO22CHD U4720 (.O(n3295), 
	.B2(n395), 
	.B1(\ram[169][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n261));
   AO22CHD U4721 (.O(n3296), 
	.B2(n395), 
	.B1(\ram[169][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n261));
   AO22CHD U4722 (.O(n3297), 
	.B2(n395), 
	.B1(\ram[169][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n261));
   AO22CHD U4723 (.O(n3298), 
	.B2(n395), 
	.B1(\ram[169][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n261));
   AO22CHD U4724 (.O(n3299), 
	.B2(n395), 
	.B1(\ram[169][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n261));
   AO22CHD U4725 (.O(n3300), 
	.B2(n395), 
	.B1(\ram[169][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n261));
   AO22CHD U4726 (.O(n3301), 
	.B2(n395), 
	.B1(\ram[169][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n261));
   AO22CHD U4727 (.O(n3302), 
	.B2(n397), 
	.B1(\ram[170][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n263));
   AO22CHD U4728 (.O(n3303), 
	.B2(n397), 
	.B1(\ram[170][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n263));
   AO22CHD U4729 (.O(n3304), 
	.B2(n397), 
	.B1(\ram[170][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n263));
   AO22CHD U4730 (.O(n3305), 
	.B2(n397), 
	.B1(\ram[170][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n263));
   AO22CHD U4731 (.O(n3306), 
	.B2(n397), 
	.B1(\ram[170][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n263));
   AO22CHD U4732 (.O(n3307), 
	.B2(n397), 
	.B1(\ram[170][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n263));
   AO22CHD U4733 (.O(n3308), 
	.B2(n397), 
	.B1(\ram[170][6] ), 
	.A2(n14), 
	.A1(n263));
   AO22CHD U4734 (.O(n3309), 
	.B2(n397), 
	.B1(\ram[170][7] ), 
	.A2(n15), 
	.A1(n263));
   AO22CHD U4735 (.O(n3310), 
	.B2(n397), 
	.B1(\ram[170][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n263));
   AO22CHD U4736 (.O(n3311), 
	.B2(n397), 
	.B1(\ram[170][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n263));
   AO22CHD U4737 (.O(n3312), 
	.B2(n397), 
	.B1(\ram[170][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n263));
   AO22CHD U4738 (.O(n3313), 
	.B2(n397), 
	.B1(\ram[170][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n263));
   AO22CHD U4739 (.O(n3314), 
	.B2(n397), 
	.B1(\ram[170][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n263));
   AO22CHD U4740 (.O(n3315), 
	.B2(n397), 
	.B1(\ram[170][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n263));
   AO22CHD U4741 (.O(n3316), 
	.B2(n397), 
	.B1(\ram[170][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n263));
   AO22CHD U4742 (.O(n3317), 
	.B2(n397), 
	.B1(\ram[170][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n263));
   AO22CHD U4743 (.O(n3318), 
	.B2(n399), 
	.B1(\ram[171][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n265));
   AO22CHD U4744 (.O(n3319), 
	.B2(n399), 
	.B1(\ram[171][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n265));
   AO22CHD U4745 (.O(n3320), 
	.B2(n399), 
	.B1(\ram[171][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n265));
   AO22CHD U4746 (.O(n3321), 
	.B2(n399), 
	.B1(\ram[171][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n265));
   AO22CHD U4747 (.O(n3322), 
	.B2(n399), 
	.B1(\ram[171][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n265));
   AO22CHD U4748 (.O(n3323), 
	.B2(n399), 
	.B1(\ram[171][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n265));
   AO22CHD U4749 (.O(n3324), 
	.B2(n399), 
	.B1(\ram[171][6] ), 
	.A2(n14), 
	.A1(n265));
   AO22CHD U4750 (.O(n3325), 
	.B2(n399), 
	.B1(\ram[171][7] ), 
	.A2(n15), 
	.A1(n265));
   AO22CHD U4751 (.O(n3326), 
	.B2(n399), 
	.B1(\ram[171][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n265));
   AO22CHD U4752 (.O(n3327), 
	.B2(n399), 
	.B1(\ram[171][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n265));
   AO22CHD U4753 (.O(n3328), 
	.B2(n399), 
	.B1(\ram[171][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n265));
   AO22CHD U4754 (.O(n3329), 
	.B2(n399), 
	.B1(\ram[171][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n265));
   AO22CHD U4755 (.O(n3330), 
	.B2(n399), 
	.B1(\ram[171][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n265));
   AO22CHD U4756 (.O(n3331), 
	.B2(n399), 
	.B1(\ram[171][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n265));
   AO22CHD U4757 (.O(n3332), 
	.B2(n399), 
	.B1(\ram[171][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n265));
   AO22CHD U4758 (.O(n3333), 
	.B2(n399), 
	.B1(\ram[171][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n265));
   AO22CHD U4759 (.O(n3334), 
	.B2(n401), 
	.B1(\ram[172][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n267));
   AO22CHD U4760 (.O(n3335), 
	.B2(n401), 
	.B1(\ram[172][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n267));
   AO22CHD U4761 (.O(n3336), 
	.B2(n401), 
	.B1(\ram[172][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n267));
   AO22CHD U4762 (.O(n3337), 
	.B2(n401), 
	.B1(\ram[172][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n267));
   AO22CHD U4763 (.O(n3338), 
	.B2(n401), 
	.B1(\ram[172][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n267));
   AO22CHD U4764 (.O(n3339), 
	.B2(n401), 
	.B1(\ram[172][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n267));
   AO22CHD U4765 (.O(n3340), 
	.B2(n401), 
	.B1(\ram[172][6] ), 
	.A2(n14), 
	.A1(n267));
   AO22CHD U4766 (.O(n3341), 
	.B2(n401), 
	.B1(\ram[172][7] ), 
	.A2(n15), 
	.A1(n267));
   AO22CHD U4767 (.O(n3342), 
	.B2(n401), 
	.B1(\ram[172][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n267));
   AO22CHD U4768 (.O(n3343), 
	.B2(n401), 
	.B1(\ram[172][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n267));
   AO22CHD U4769 (.O(n3344), 
	.B2(n401), 
	.B1(\ram[172][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n267));
   AO22CHD U4770 (.O(n3345), 
	.B2(n401), 
	.B1(\ram[172][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n267));
   AO22CHD U4771 (.O(n3346), 
	.B2(n401), 
	.B1(\ram[172][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n267));
   AO22CHD U4772 (.O(n3347), 
	.B2(n401), 
	.B1(\ram[172][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n267));
   AO22CHD U4773 (.O(n3348), 
	.B2(n401), 
	.B1(\ram[172][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n267));
   AO22CHD U4774 (.O(n3349), 
	.B2(n401), 
	.B1(\ram[172][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n267));
   AO22CHD U4775 (.O(n3350), 
	.B2(n403), 
	.B1(\ram[173][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n269));
   AO22CHD U4776 (.O(n3351), 
	.B2(n403), 
	.B1(\ram[173][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n269));
   AO22CHD U4777 (.O(n3352), 
	.B2(n403), 
	.B1(\ram[173][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n269));
   AO22CHD U4778 (.O(n3353), 
	.B2(n403), 
	.B1(\ram[173][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n269));
   AO22CHD U4779 (.O(n3354), 
	.B2(n403), 
	.B1(\ram[173][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n269));
   AO22CHD U4780 (.O(n3355), 
	.B2(n403), 
	.B1(\ram[173][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n269));
   AO22CHD U4781 (.O(n3356), 
	.B2(n403), 
	.B1(\ram[173][6] ), 
	.A2(n14), 
	.A1(n269));
   AO22CHD U4782 (.O(n3357), 
	.B2(n403), 
	.B1(\ram[173][7] ), 
	.A2(n15), 
	.A1(n269));
   AO22CHD U4783 (.O(n3358), 
	.B2(n403), 
	.B1(\ram[173][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n269));
   AO22CHD U4784 (.O(n3359), 
	.B2(n403), 
	.B1(\ram[173][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n269));
   AO22CHD U4785 (.O(n3360), 
	.B2(n403), 
	.B1(\ram[173][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n269));
   AO22CHD U4786 (.O(n3361), 
	.B2(n403), 
	.B1(\ram[173][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n269));
   AO22CHD U4787 (.O(n3362), 
	.B2(n403), 
	.B1(\ram[173][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n269));
   AO22CHD U4788 (.O(n3363), 
	.B2(n403), 
	.B1(\ram[173][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n269));
   AO22CHD U4789 (.O(n3364), 
	.B2(n403), 
	.B1(\ram[173][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n269));
   AO22CHD U4790 (.O(n3365), 
	.B2(n403), 
	.B1(\ram[173][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n269));
   AO22CHD U4791 (.O(n3366), 
	.B2(n405), 
	.B1(\ram[174][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n271));
   AO22CHD U4792 (.O(n3367), 
	.B2(n405), 
	.B1(\ram[174][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n271));
   AO22CHD U4793 (.O(n3368), 
	.B2(n405), 
	.B1(\ram[174][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n271));
   AO22CHD U4794 (.O(n3369), 
	.B2(n405), 
	.B1(\ram[174][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n271));
   AO22CHD U4795 (.O(n3370), 
	.B2(n405), 
	.B1(\ram[174][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n271));
   AO22CHD U4796 (.O(n3371), 
	.B2(n405), 
	.B1(\ram[174][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n271));
   AO22CHD U4797 (.O(n3372), 
	.B2(n405), 
	.B1(\ram[174][6] ), 
	.A2(n14), 
	.A1(n271));
   AO22CHD U4798 (.O(n3373), 
	.B2(n405), 
	.B1(\ram[174][7] ), 
	.A2(n15), 
	.A1(n271));
   AO22CHD U4799 (.O(n3374), 
	.B2(n405), 
	.B1(\ram[174][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n271));
   AO22CHD U4800 (.O(n3375), 
	.B2(n405), 
	.B1(\ram[174][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n271));
   AO22CHD U4801 (.O(n3376), 
	.B2(n405), 
	.B1(\ram[174][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n271));
   AO22CHD U4802 (.O(n3377), 
	.B2(n405), 
	.B1(\ram[174][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n271));
   AO22CHD U4803 (.O(n3378), 
	.B2(n405), 
	.B1(\ram[174][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n271));
   AO22CHD U4804 (.O(n3379), 
	.B2(n405), 
	.B1(\ram[174][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n271));
   AO22CHD U4805 (.O(n3380), 
	.B2(n405), 
	.B1(\ram[174][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n271));
   AO22CHD U4806 (.O(n3381), 
	.B2(n405), 
	.B1(\ram[174][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n271));
   AO22CHD U4807 (.O(n3382), 
	.B2(n407), 
	.B1(\ram[175][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n273));
   AO22CHD U4808 (.O(n3383), 
	.B2(n407), 
	.B1(\ram[175][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n273));
   AO22CHD U4809 (.O(n3384), 
	.B2(n407), 
	.B1(\ram[175][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n273));
   AO22CHD U4810 (.O(n3385), 
	.B2(n407), 
	.B1(\ram[175][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n273));
   AO22CHD U4811 (.O(n3386), 
	.B2(n407), 
	.B1(\ram[175][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n273));
   AO22CHD U4812 (.O(n3387), 
	.B2(n407), 
	.B1(\ram[175][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n273));
   AO22CHD U4813 (.O(n3388), 
	.B2(n407), 
	.B1(\ram[175][6] ), 
	.A2(n14), 
	.A1(n273));
   AO22CHD U4814 (.O(n3389), 
	.B2(n407), 
	.B1(\ram[175][7] ), 
	.A2(n15), 
	.A1(n273));
   AO22CHD U4815 (.O(n3390), 
	.B2(n407), 
	.B1(\ram[175][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n273));
   AO22CHD U4816 (.O(n3391), 
	.B2(n407), 
	.B1(\ram[175][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n273));
   AO22CHD U4817 (.O(n3392), 
	.B2(n407), 
	.B1(\ram[175][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n273));
   AO22CHD U4818 (.O(n3393), 
	.B2(n407), 
	.B1(\ram[175][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n273));
   AO22CHD U4819 (.O(n3394), 
	.B2(n407), 
	.B1(\ram[175][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n273));
   AO22CHD U4820 (.O(n3395), 
	.B2(n407), 
	.B1(\ram[175][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n273));
   AO22CHD U4821 (.O(n3396), 
	.B2(n407), 
	.B1(\ram[175][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n273));
   AO22CHD U4822 (.O(n3397), 
	.B2(n407), 
	.B1(\ram[175][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n273));
   AO22CHD U4823 (.O(n3398), 
	.B2(n409), 
	.B1(\ram[176][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n275));
   AO22CHD U4824 (.O(n3399), 
	.B2(n409), 
	.B1(\ram[176][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n275));
   AO22CHD U4825 (.O(n3400), 
	.B2(n409), 
	.B1(\ram[176][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n275));
   AO22CHD U4826 (.O(n3401), 
	.B2(n409), 
	.B1(\ram[176][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n275));
   AO22CHD U4827 (.O(n3402), 
	.B2(n409), 
	.B1(\ram[176][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n275));
   AO22CHD U4828 (.O(n3403), 
	.B2(n409), 
	.B1(\ram[176][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n275));
   AO22CHD U4829 (.O(n3404), 
	.B2(n409), 
	.B1(\ram[176][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n275));
   AO22CHD U4830 (.O(n3405), 
	.B2(n409), 
	.B1(\ram[176][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n275));
   AO22CHD U4831 (.O(n3406), 
	.B2(n409), 
	.B1(\ram[176][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n275));
   AO22CHD U4832 (.O(n3407), 
	.B2(n409), 
	.B1(\ram[176][9] ), 
	.A2(n17), 
	.A1(n275));
   AO22CHD U4833 (.O(n3408), 
	.B2(n409), 
	.B1(\ram[176][10] ), 
	.A2(n18), 
	.A1(n275));
   AO22CHD U4834 (.O(n3409), 
	.B2(n409), 
	.B1(\ram[176][11] ), 
	.A2(n19), 
	.A1(n275));
   AO22CHD U4835 (.O(n3410), 
	.B2(n409), 
	.B1(\ram[176][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n275));
   AO22CHD U4836 (.O(n3411), 
	.B2(n409), 
	.B1(\ram[176][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n275));
   AO22CHD U4837 (.O(n3412), 
	.B2(n409), 
	.B1(\ram[176][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n275));
   AO22CHD U4838 (.O(n3413), 
	.B2(n409), 
	.B1(\ram[176][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n275));
   AO22CHD U4839 (.O(n3414), 
	.B2(n412), 
	.B1(\ram[177][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n277));
   AO22CHD U4840 (.O(n3415), 
	.B2(n412), 
	.B1(\ram[177][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n277));
   AO22CHD U4841 (.O(n3416), 
	.B2(n412), 
	.B1(\ram[177][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n277));
   AO22CHD U4842 (.O(n3417), 
	.B2(n412), 
	.B1(\ram[177][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n277));
   AO22CHD U4843 (.O(n3418), 
	.B2(n412), 
	.B1(\ram[177][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n277));
   AO22CHD U4844 (.O(n3419), 
	.B2(n412), 
	.B1(\ram[177][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n277));
   AO22CHD U4845 (.O(n3420), 
	.B2(n412), 
	.B1(\ram[177][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n277));
   AO22CHD U4846 (.O(n3421), 
	.B2(n412), 
	.B1(\ram[177][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n277));
   AO22CHD U4847 (.O(n3422), 
	.B2(n412), 
	.B1(\ram[177][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n277));
   AO22CHD U4848 (.O(n3423), 
	.B2(n412), 
	.B1(\ram[177][9] ), 
	.A2(n17), 
	.A1(n277));
   AO22CHD U4849 (.O(n3424), 
	.B2(n412), 
	.B1(\ram[177][10] ), 
	.A2(n18), 
	.A1(n277));
   AO22CHD U4850 (.O(n3425), 
	.B2(n412), 
	.B1(\ram[177][11] ), 
	.A2(n19), 
	.A1(n277));
   AO22CHD U4851 (.O(n3426), 
	.B2(n412), 
	.B1(\ram[177][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n277));
   AO22CHD U4852 (.O(n3427), 
	.B2(n412), 
	.B1(\ram[177][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n277));
   AO22CHD U4853 (.O(n3428), 
	.B2(n412), 
	.B1(\ram[177][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n277));
   AO22CHD U4854 (.O(n3429), 
	.B2(n412), 
	.B1(\ram[177][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n277));
   AO22CHD U4855 (.O(n3430), 
	.B2(n414), 
	.B1(\ram[178][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n278));
   AO22CHD U4856 (.O(n3431), 
	.B2(n414), 
	.B1(\ram[178][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n278));
   AO22CHD U4857 (.O(n3432), 
	.B2(n414), 
	.B1(\ram[178][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n278));
   AO22CHD U4858 (.O(n3433), 
	.B2(n414), 
	.B1(\ram[178][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n278));
   AO22CHD U4859 (.O(n3434), 
	.B2(n414), 
	.B1(\ram[178][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n278));
   AO22CHD U4860 (.O(n3435), 
	.B2(n414), 
	.B1(\ram[178][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n278));
   AO22CHD U4861 (.O(n3436), 
	.B2(n414), 
	.B1(\ram[178][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n278));
   AO22CHD U4862 (.O(n3437), 
	.B2(n414), 
	.B1(\ram[178][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n278));
   AO22CHD U4863 (.O(n3438), 
	.B2(n414), 
	.B1(\ram[178][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n278));
   AO22CHD U4864 (.O(n3439), 
	.B2(n414), 
	.B1(\ram[178][9] ), 
	.A2(n17), 
	.A1(n278));
   AO22CHD U4865 (.O(n3440), 
	.B2(n414), 
	.B1(\ram[178][10] ), 
	.A2(n18), 
	.A1(n278));
   AO22CHD U4866 (.O(n3441), 
	.B2(n414), 
	.B1(\ram[178][11] ), 
	.A2(n19), 
	.A1(n278));
   AO22CHD U4867 (.O(n3442), 
	.B2(n414), 
	.B1(\ram[178][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n278));
   AO22CHD U4868 (.O(n3443), 
	.B2(n414), 
	.B1(\ram[178][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n278));
   AO22CHD U4869 (.O(n3444), 
	.B2(n414), 
	.B1(\ram[178][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n278));
   AO22CHD U4870 (.O(n3445), 
	.B2(n414), 
	.B1(\ram[178][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n278));
   AO22CHD U4871 (.O(n3446), 
	.B2(n416), 
	.B1(\ram[179][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n280));
   AO22CHD U4872 (.O(n3447), 
	.B2(n416), 
	.B1(\ram[179][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n280));
   AO22CHD U4873 (.O(n3448), 
	.B2(n416), 
	.B1(\ram[179][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n280));
   AO22CHD U4874 (.O(n3449), 
	.B2(n416), 
	.B1(\ram[179][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n280));
   AO22CHD U4875 (.O(n3450), 
	.B2(n416), 
	.B1(\ram[179][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n280));
   AO22CHD U4876 (.O(n3451), 
	.B2(n416), 
	.B1(\ram[179][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n280));
   AO22CHD U4877 (.O(n3452), 
	.B2(n416), 
	.B1(\ram[179][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n280));
   AO22CHD U4878 (.O(n3453), 
	.B2(n416), 
	.B1(\ram[179][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n280));
   AO22CHD U4879 (.O(n3454), 
	.B2(n416), 
	.B1(\ram[179][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n280));
   AO22CHD U4880 (.O(n3455), 
	.B2(n416), 
	.B1(\ram[179][9] ), 
	.A2(n17), 
	.A1(n280));
   AO22CHD U4881 (.O(n3456), 
	.B2(n416), 
	.B1(\ram[179][10] ), 
	.A2(n18), 
	.A1(n280));
   AO22CHD U4882 (.O(n3457), 
	.B2(n416), 
	.B1(\ram[179][11] ), 
	.A2(n19), 
	.A1(n280));
   AO22CHD U4883 (.O(n3458), 
	.B2(n416), 
	.B1(\ram[179][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n280));
   AO22CHD U4884 (.O(n3459), 
	.B2(n416), 
	.B1(\ram[179][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n280));
   AO22CHD U4885 (.O(n3460), 
	.B2(n416), 
	.B1(\ram[179][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n280));
   AO22CHD U4886 (.O(n3461), 
	.B2(n416), 
	.B1(\ram[179][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n280));
   AO22CHD U4887 (.O(n3462), 
	.B2(n418), 
	.B1(\ram[180][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n282));
   AO22CHD U4888 (.O(n3463), 
	.B2(n418), 
	.B1(\ram[180][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n282));
   AO22CHD U4889 (.O(n3464), 
	.B2(n418), 
	.B1(\ram[180][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n282));
   AO22CHD U4890 (.O(n3465), 
	.B2(n418), 
	.B1(\ram[180][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n282));
   AO22CHD U4891 (.O(n3466), 
	.B2(n418), 
	.B1(\ram[180][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n282));
   AO22CHD U4892 (.O(n3467), 
	.B2(n418), 
	.B1(\ram[180][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n282));
   AO22CHD U4893 (.O(n3468), 
	.B2(n418), 
	.B1(\ram[180][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n282));
   AO22CHD U4894 (.O(n3469), 
	.B2(n418), 
	.B1(\ram[180][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n282));
   AO22CHD U4895 (.O(n3470), 
	.B2(n418), 
	.B1(\ram[180][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n282));
   AO22CHD U4896 (.O(n3471), 
	.B2(n418), 
	.B1(\ram[180][9] ), 
	.A2(n17), 
	.A1(n282));
   AO22CHD U4897 (.O(n3472), 
	.B2(n418), 
	.B1(\ram[180][10] ), 
	.A2(n18), 
	.A1(n282));
   AO22CHD U4898 (.O(n3473), 
	.B2(n418), 
	.B1(\ram[180][11] ), 
	.A2(n19), 
	.A1(n282));
   AO22CHD U4899 (.O(n3474), 
	.B2(n418), 
	.B1(\ram[180][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n282));
   AO22CHD U4900 (.O(n3475), 
	.B2(n418), 
	.B1(\ram[180][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n282));
   AO22CHD U4901 (.O(n3476), 
	.B2(n418), 
	.B1(\ram[180][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n282));
   AO22CHD U4902 (.O(n3477), 
	.B2(n418), 
	.B1(\ram[180][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n282));
   AO22CHD U4903 (.O(n3478), 
	.B2(n420), 
	.B1(\ram[181][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n284));
   AO22CHD U4904 (.O(n3479), 
	.B2(n420), 
	.B1(\ram[181][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n284));
   AO22CHD U4905 (.O(n3480), 
	.B2(n420), 
	.B1(\ram[181][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n284));
   AO22CHD U4906 (.O(n3481), 
	.B2(n420), 
	.B1(\ram[181][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n284));
   AO22CHD U4907 (.O(n3482), 
	.B2(n420), 
	.B1(\ram[181][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n284));
   AO22CHD U4908 (.O(n3483), 
	.B2(n420), 
	.B1(\ram[181][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n284));
   AO22CHD U4909 (.O(n3484), 
	.B2(n420), 
	.B1(\ram[181][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n284));
   AO22CHD U4910 (.O(n3485), 
	.B2(n420), 
	.B1(\ram[181][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n284));
   AO22CHD U4911 (.O(n3486), 
	.B2(n420), 
	.B1(\ram[181][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n284));
   AO22CHD U4912 (.O(n3487), 
	.B2(n420), 
	.B1(\ram[181][9] ), 
	.A2(n17), 
	.A1(n284));
   AO22CHD U4913 (.O(n3488), 
	.B2(n420), 
	.B1(\ram[181][10] ), 
	.A2(n18), 
	.A1(n284));
   AO22CHD U4914 (.O(n3489), 
	.B2(n420), 
	.B1(\ram[181][11] ), 
	.A2(n19), 
	.A1(n284));
   AO22CHD U4915 (.O(n3490), 
	.B2(n420), 
	.B1(\ram[181][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n284));
   AO22CHD U4916 (.O(n3491), 
	.B2(n420), 
	.B1(\ram[181][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n284));
   AO22CHD U4917 (.O(n3492), 
	.B2(n420), 
	.B1(\ram[181][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n284));
   AO22CHD U4918 (.O(n3493), 
	.B2(n420), 
	.B1(\ram[181][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n284));
   AO22CHD U4919 (.O(n3494), 
	.B2(n422), 
	.B1(\ram[182][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n286));
   AO22CHD U4920 (.O(n3495), 
	.B2(n422), 
	.B1(\ram[182][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n286));
   AO22CHD U4921 (.O(n3496), 
	.B2(n422), 
	.B1(\ram[182][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n286));
   AO22CHD U4922 (.O(n3497), 
	.B2(n422), 
	.B1(\ram[182][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n286));
   AO22CHD U4923 (.O(n3498), 
	.B2(n422), 
	.B1(\ram[182][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n286));
   AO22CHD U4924 (.O(n3499), 
	.B2(n422), 
	.B1(\ram[182][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n286));
   AO22CHD U4925 (.O(n3500), 
	.B2(n422), 
	.B1(\ram[182][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n286));
   AO22CHD U4926 (.O(n3501), 
	.B2(n422), 
	.B1(\ram[182][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n286));
   AO22CHD U4927 (.O(n3502), 
	.B2(n422), 
	.B1(\ram[182][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n286));
   AO22CHD U4928 (.O(n3503), 
	.B2(n422), 
	.B1(\ram[182][9] ), 
	.A2(n17), 
	.A1(n286));
   AO22CHD U4929 (.O(n3504), 
	.B2(n422), 
	.B1(\ram[182][10] ), 
	.A2(n18), 
	.A1(n286));
   AO22CHD U4930 (.O(n3505), 
	.B2(n422), 
	.B1(\ram[182][11] ), 
	.A2(n19), 
	.A1(n286));
   AO22CHD U4931 (.O(n3506), 
	.B2(n422), 
	.B1(\ram[182][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n286));
   AO22CHD U4932 (.O(n3507), 
	.B2(n422), 
	.B1(\ram[182][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n286));
   AO22CHD U4933 (.O(n3508), 
	.B2(n422), 
	.B1(\ram[182][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n286));
   AO22CHD U4934 (.O(n3509), 
	.B2(n422), 
	.B1(\ram[182][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n286));
   AO22CHD U4935 (.O(n3510), 
	.B2(n424), 
	.B1(\ram[183][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n288));
   AO22CHD U4936 (.O(n3511), 
	.B2(n424), 
	.B1(\ram[183][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n288));
   AO22CHD U4937 (.O(n3512), 
	.B2(n424), 
	.B1(\ram[183][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n288));
   AO22CHD U4938 (.O(n3513), 
	.B2(n424), 
	.B1(\ram[183][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n288));
   AO22CHD U4939 (.O(n3514), 
	.B2(n424), 
	.B1(\ram[183][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n288));
   AO22CHD U4940 (.O(n3515), 
	.B2(n424), 
	.B1(\ram[183][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n288));
   AO22CHD U4941 (.O(n3516), 
	.B2(n424), 
	.B1(\ram[183][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n288));
   AO22CHD U4942 (.O(n3517), 
	.B2(n424), 
	.B1(\ram[183][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n288));
   AO22CHD U4943 (.O(n3518), 
	.B2(n424), 
	.B1(\ram[183][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n288));
   AO22CHD U4944 (.O(n3519), 
	.B2(n424), 
	.B1(\ram[183][9] ), 
	.A2(n17), 
	.A1(n288));
   AO22CHD U4945 (.O(n3520), 
	.B2(n424), 
	.B1(\ram[183][10] ), 
	.A2(n18), 
	.A1(n288));
   AO22CHD U4946 (.O(n3521), 
	.B2(n424), 
	.B1(\ram[183][11] ), 
	.A2(n19), 
	.A1(n288));
   AO22CHD U4947 (.O(n3522), 
	.B2(n424), 
	.B1(\ram[183][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n288));
   AO22CHD U4948 (.O(n3523), 
	.B2(n424), 
	.B1(\ram[183][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n288));
   AO22CHD U4949 (.O(n3524), 
	.B2(n424), 
	.B1(\ram[183][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n288));
   AO22CHD U4950 (.O(n3525), 
	.B2(n424), 
	.B1(\ram[183][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n288));
   AO22CHD U4951 (.O(n3526), 
	.B2(n426), 
	.B1(\ram[184][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n290));
   AO22CHD U4952 (.O(n3527), 
	.B2(n426), 
	.B1(\ram[184][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n290));
   AO22CHD U4953 (.O(n3528), 
	.B2(n426), 
	.B1(\ram[184][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n290));
   AO22CHD U4954 (.O(n3529), 
	.B2(n426), 
	.B1(\ram[184][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n290));
   AO22CHD U4955 (.O(n3530), 
	.B2(n426), 
	.B1(\ram[184][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n290));
   AO22CHD U4956 (.O(n3531), 
	.B2(n426), 
	.B1(\ram[184][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n290));
   AO22CHD U4957 (.O(n3532), 
	.B2(n426), 
	.B1(\ram[184][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n290));
   AO22CHD U4958 (.O(n3533), 
	.B2(n426), 
	.B1(\ram[184][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n290));
   AO22CHD U4959 (.O(n3534), 
	.B2(n426), 
	.B1(\ram[184][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n290));
   AO22CHD U4960 (.O(n3535), 
	.B2(n426), 
	.B1(\ram[184][9] ), 
	.A2(n17), 
	.A1(n290));
   AO22CHD U4961 (.O(n3536), 
	.B2(n426), 
	.B1(\ram[184][10] ), 
	.A2(n18), 
	.A1(n290));
   AO22CHD U4962 (.O(n3537), 
	.B2(n426), 
	.B1(\ram[184][11] ), 
	.A2(n19), 
	.A1(n290));
   AO22CHD U4963 (.O(n3538), 
	.B2(n426), 
	.B1(\ram[184][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n290));
   AO22CHD U4964 (.O(n3539), 
	.B2(n426), 
	.B1(\ram[184][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n290));
   AO22CHD U4965 (.O(n3540), 
	.B2(n426), 
	.B1(\ram[184][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n290));
   AO22CHD U4966 (.O(n3541), 
	.B2(n426), 
	.B1(\ram[184][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n290));
   AO22CHD U4967 (.O(n3542), 
	.B2(n428), 
	.B1(\ram[185][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n292));
   AO22CHD U4968 (.O(n3543), 
	.B2(n428), 
	.B1(\ram[185][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n292));
   AO22CHD U4969 (.O(n3544), 
	.B2(n428), 
	.B1(\ram[185][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n292));
   AO22CHD U4970 (.O(n3545), 
	.B2(n428), 
	.B1(\ram[185][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n292));
   AO22CHD U4971 (.O(n3546), 
	.B2(n428), 
	.B1(\ram[185][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n292));
   AO22CHD U4972 (.O(n3547), 
	.B2(n428), 
	.B1(\ram[185][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n292));
   AO22CHD U4973 (.O(n3548), 
	.B2(n428), 
	.B1(\ram[185][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n292));
   AO22CHD U4974 (.O(n3549), 
	.B2(n428), 
	.B1(\ram[185][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n292));
   AO22CHD U4975 (.O(n3550), 
	.B2(n428), 
	.B1(\ram[185][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n292));
   AO22CHD U4976 (.O(n3551), 
	.B2(n428), 
	.B1(\ram[185][9] ), 
	.A2(n17), 
	.A1(n292));
   AO22CHD U4977 (.O(n3552), 
	.B2(n428), 
	.B1(\ram[185][10] ), 
	.A2(n18), 
	.A1(n292));
   AO22CHD U4978 (.O(n3553), 
	.B2(n428), 
	.B1(\ram[185][11] ), 
	.A2(n19), 
	.A1(n292));
   AO22CHD U4979 (.O(n3554), 
	.B2(n428), 
	.B1(\ram[185][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n292));
   AO22CHD U4980 (.O(n3555), 
	.B2(n428), 
	.B1(\ram[185][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n292));
   AO22CHD U4981 (.O(n3556), 
	.B2(n428), 
	.B1(\ram[185][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n292));
   AO22CHD U4982 (.O(n3557), 
	.B2(n428), 
	.B1(\ram[185][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n292));
   AO22CHD U4983 (.O(n3558), 
	.B2(n430), 
	.B1(\ram[186][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n294));
   AO22CHD U4984 (.O(n3559), 
	.B2(n430), 
	.B1(\ram[186][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n294));
   AO22CHD U4985 (.O(n3560), 
	.B2(n430), 
	.B1(\ram[186][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n294));
   AO22CHD U4986 (.O(n3561), 
	.B2(n430), 
	.B1(\ram[186][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n294));
   AO22CHD U4987 (.O(n3562), 
	.B2(n430), 
	.B1(\ram[186][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n294));
   AO22CHD U4988 (.O(n3563), 
	.B2(n430), 
	.B1(\ram[186][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n294));
   AO22CHD U4989 (.O(n3564), 
	.B2(n430), 
	.B1(\ram[186][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n294));
   AO22CHD U4990 (.O(n3565), 
	.B2(n430), 
	.B1(\ram[186][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n294));
   AO22CHD U4991 (.O(n3566), 
	.B2(n430), 
	.B1(\ram[186][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n294));
   AO22CHD U4992 (.O(n3567), 
	.B2(n430), 
	.B1(\ram[186][9] ), 
	.A2(n17), 
	.A1(n294));
   AO22CHD U4993 (.O(n3568), 
	.B2(n430), 
	.B1(\ram[186][10] ), 
	.A2(n18), 
	.A1(n294));
   AO22CHD U4994 (.O(n3569), 
	.B2(n430), 
	.B1(\ram[186][11] ), 
	.A2(n19), 
	.A1(n294));
   AO22CHD U4995 (.O(n3570), 
	.B2(n430), 
	.B1(\ram[186][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n294));
   AO22CHD U4996 (.O(n3571), 
	.B2(n430), 
	.B1(\ram[186][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n294));
   AO22CHD U4997 (.O(n3572), 
	.B2(n430), 
	.B1(\ram[186][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n294));
   AO22CHD U4998 (.O(n3573), 
	.B2(n430), 
	.B1(\ram[186][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n294));
   AO22CHD U4999 (.O(n3574), 
	.B2(n432), 
	.B1(\ram[187][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n296));
   AO22CHD U5000 (.O(n3575), 
	.B2(n432), 
	.B1(\ram[187][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n296));
   AO22CHD U5001 (.O(n3576), 
	.B2(n432), 
	.B1(\ram[187][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n296));
   AO22CHD U5002 (.O(n3577), 
	.B2(n432), 
	.B1(\ram[187][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n296));
   AO22CHD U5003 (.O(n3578), 
	.B2(n432), 
	.B1(\ram[187][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n296));
   AO22CHD U5004 (.O(n3579), 
	.B2(n432), 
	.B1(\ram[187][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n296));
   AO22CHD U5005 (.O(n3580), 
	.B2(n432), 
	.B1(\ram[187][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n296));
   AO22CHD U5006 (.O(n3581), 
	.B2(n432), 
	.B1(\ram[187][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n296));
   AO22CHD U5007 (.O(n3582), 
	.B2(n432), 
	.B1(\ram[187][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n296));
   AO22CHD U5008 (.O(n3583), 
	.B2(n432), 
	.B1(\ram[187][9] ), 
	.A2(n17), 
	.A1(n296));
   AO22CHD U5009 (.O(n3584), 
	.B2(n432), 
	.B1(\ram[187][10] ), 
	.A2(n18), 
	.A1(n296));
   AO22CHD U5010 (.O(n3585), 
	.B2(n432), 
	.B1(\ram[187][11] ), 
	.A2(n19), 
	.A1(n296));
   AO22CHD U5011 (.O(n3586), 
	.B2(n432), 
	.B1(\ram[187][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n296));
   AO22CHD U5012 (.O(n3587), 
	.B2(n432), 
	.B1(\ram[187][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n296));
   AO22CHD U5013 (.O(n3588), 
	.B2(n432), 
	.B1(\ram[187][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n296));
   AO22CHD U5014 (.O(n3589), 
	.B2(n432), 
	.B1(\ram[187][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n296));
   AO22CHD U5015 (.O(n3590), 
	.B2(n434), 
	.B1(\ram[188][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n298));
   AO22CHD U5016 (.O(n3591), 
	.B2(n434), 
	.B1(\ram[188][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n298));
   AO22CHD U5017 (.O(n3592), 
	.B2(n434), 
	.B1(\ram[188][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n298));
   AO22CHD U5018 (.O(n3593), 
	.B2(n434), 
	.B1(\ram[188][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n298));
   AO22CHD U5019 (.O(n3594), 
	.B2(n434), 
	.B1(\ram[188][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n298));
   AO22CHD U5020 (.O(n3595), 
	.B2(n434), 
	.B1(\ram[188][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n298));
   AO22CHD U5021 (.O(n3596), 
	.B2(n434), 
	.B1(\ram[188][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n298));
   AO22CHD U5022 (.O(n3597), 
	.B2(n434), 
	.B1(\ram[188][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n298));
   AO22CHD U5023 (.O(n3598), 
	.B2(n434), 
	.B1(\ram[188][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n298));
   AO22CHD U5024 (.O(n3599), 
	.B2(n434), 
	.B1(\ram[188][9] ), 
	.A2(n17), 
	.A1(n298));
   AO22CHD U5025 (.O(n3600), 
	.B2(n434), 
	.B1(\ram[188][10] ), 
	.A2(n18), 
	.A1(n298));
   AO22CHD U5026 (.O(n3601), 
	.B2(n434), 
	.B1(\ram[188][11] ), 
	.A2(n19), 
	.A1(n298));
   AO22CHD U5027 (.O(n3602), 
	.B2(n434), 
	.B1(\ram[188][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n298));
   AO22CHD U5028 (.O(n3603), 
	.B2(n434), 
	.B1(\ram[188][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n298));
   AO22CHD U5029 (.O(n3604), 
	.B2(n434), 
	.B1(\ram[188][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n298));
   AO22CHD U5030 (.O(n3605), 
	.B2(n434), 
	.B1(\ram[188][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n298));
   AO22CHD U5031 (.O(n3606), 
	.B2(n436), 
	.B1(\ram[189][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n300));
   AO22CHD U5032 (.O(n3607), 
	.B2(n436), 
	.B1(\ram[189][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n300));
   AO22CHD U5033 (.O(n3608), 
	.B2(n436), 
	.B1(\ram[189][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n300));
   AO22CHD U5034 (.O(n3609), 
	.B2(n436), 
	.B1(\ram[189][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n300));
   AO22CHD U5035 (.O(n3610), 
	.B2(n436), 
	.B1(\ram[189][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n300));
   AO22CHD U5036 (.O(n3611), 
	.B2(n436), 
	.B1(\ram[189][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n300));
   AO22CHD U5037 (.O(n3612), 
	.B2(n436), 
	.B1(\ram[189][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n300));
   AO22CHD U5038 (.O(n3613), 
	.B2(n436), 
	.B1(\ram[189][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n300));
   AO22CHD U5039 (.O(n3614), 
	.B2(n436), 
	.B1(\ram[189][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n300));
   AO22CHD U5040 (.O(n3615), 
	.B2(n436), 
	.B1(\ram[189][9] ), 
	.A2(n17), 
	.A1(n300));
   AO22CHD U5041 (.O(n3616), 
	.B2(n436), 
	.B1(\ram[189][10] ), 
	.A2(n18), 
	.A1(n300));
   AO22CHD U5042 (.O(n3617), 
	.B2(n436), 
	.B1(\ram[189][11] ), 
	.A2(n19), 
	.A1(n300));
   AO22CHD U5043 (.O(n3618), 
	.B2(n436), 
	.B1(\ram[189][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n300));
   AO22CHD U5044 (.O(n3619), 
	.B2(n436), 
	.B1(\ram[189][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n300));
   AO22CHD U5045 (.O(n3620), 
	.B2(n436), 
	.B1(\ram[189][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n300));
   AO22CHD U5046 (.O(n3621), 
	.B2(n436), 
	.B1(\ram[189][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n300));
   AO22CHD U5047 (.O(n3622), 
	.B2(n438), 
	.B1(\ram[190][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n302));
   AO22CHD U5048 (.O(n3623), 
	.B2(n438), 
	.B1(\ram[190][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n302));
   AO22CHD U5049 (.O(n3624), 
	.B2(n438), 
	.B1(\ram[190][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n302));
   AO22CHD U5050 (.O(n3625), 
	.B2(n438), 
	.B1(\ram[190][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n302));
   AO22CHD U5051 (.O(n3626), 
	.B2(n438), 
	.B1(\ram[190][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n302));
   AO22CHD U5052 (.O(n3627), 
	.B2(n438), 
	.B1(\ram[190][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n302));
   AO22CHD U5053 (.O(n3628), 
	.B2(n438), 
	.B1(\ram[190][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n302));
   AO22CHD U5054 (.O(n3629), 
	.B2(n438), 
	.B1(\ram[190][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n302));
   AO22CHD U5055 (.O(n3630), 
	.B2(n438), 
	.B1(\ram[190][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n302));
   AO22CHD U5056 (.O(n3631), 
	.B2(n438), 
	.B1(\ram[190][9] ), 
	.A2(n17), 
	.A1(n302));
   AO22CHD U5057 (.O(n3632), 
	.B2(n438), 
	.B1(\ram[190][10] ), 
	.A2(n18), 
	.A1(n302));
   AO22CHD U5058 (.O(n3633), 
	.B2(n438), 
	.B1(\ram[190][11] ), 
	.A2(n19), 
	.A1(n302));
   AO22CHD U5059 (.O(n3634), 
	.B2(n438), 
	.B1(\ram[190][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n302));
   AO22CHD U5060 (.O(n3635), 
	.B2(n438), 
	.B1(\ram[190][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n302));
   AO22CHD U5061 (.O(n3636), 
	.B2(n438), 
	.B1(\ram[190][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n302));
   AO22CHD U5062 (.O(n3637), 
	.B2(n438), 
	.B1(\ram[190][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n302));
   AO22CHD U5063 (.O(n3638), 
	.B2(n440), 
	.B1(\ram[191][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n304));
   AO22CHD U5064 (.O(n3639), 
	.B2(n440), 
	.B1(\ram[191][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n304));
   AO22CHD U5065 (.O(n3640), 
	.B2(n440), 
	.B1(\ram[191][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n304));
   AO22CHD U5066 (.O(n3641), 
	.B2(n440), 
	.B1(\ram[191][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n304));
   AO22CHD U5067 (.O(n3642), 
	.B2(n440), 
	.B1(\ram[191][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n304));
   AO22CHD U5068 (.O(n3643), 
	.B2(n440), 
	.B1(\ram[191][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n304));
   AO22CHD U5069 (.O(n3644), 
	.B2(n440), 
	.B1(\ram[191][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n304));
   AO22CHD U5070 (.O(n3645), 
	.B2(n440), 
	.B1(\ram[191][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n304));
   AO22CHD U5071 (.O(n3646), 
	.B2(n440), 
	.B1(\ram[191][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n304));
   AO22CHD U5072 (.O(n3647), 
	.B2(n440), 
	.B1(\ram[191][9] ), 
	.A2(n17), 
	.A1(n304));
   AO22CHD U5073 (.O(n3648), 
	.B2(n440), 
	.B1(\ram[191][10] ), 
	.A2(n18), 
	.A1(n304));
   AO22CHD U5074 (.O(n3649), 
	.B2(n440), 
	.B1(\ram[191][11] ), 
	.A2(n19), 
	.A1(n304));
   AO22CHD U5075 (.O(n3650), 
	.B2(n440), 
	.B1(\ram[191][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n304));
   AO22CHD U5076 (.O(n3651), 
	.B2(n440), 
	.B1(\ram[191][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n304));
   AO22CHD U5077 (.O(n3652), 
	.B2(n440), 
	.B1(\ram[191][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n304));
   AO22CHD U5078 (.O(n3653), 
	.B2(n440), 
	.B1(\ram[191][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n304));
   AO22CHD U5079 (.O(n3654), 
	.B2(n442), 
	.B1(\ram[192][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n306));
   AO22CHD U5080 (.O(n3655), 
	.B2(n442), 
	.B1(\ram[192][1] ), 
	.A2(n9), 
	.A1(n306));
   AO22CHD U5081 (.O(n3656), 
	.B2(n442), 
	.B1(\ram[192][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n306));
   AO22CHD U5082 (.O(n3657), 
	.B2(n442), 
	.B1(\ram[192][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n306));
   AO22CHD U5083 (.O(n3658), 
	.B2(n442), 
	.B1(\ram[192][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n306));
   AO22CHD U5084 (.O(n3659), 
	.B2(n442), 
	.B1(\ram[192][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n306));
   AO22CHD U5085 (.O(n3660), 
	.B2(n442), 
	.B1(\ram[192][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n306));
   AO22CHD U5086 (.O(n3661), 
	.B2(n442), 
	.B1(\ram[192][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n306));
   AO22CHD U5087 (.O(n3662), 
	.B2(n442), 
	.B1(\ram[192][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n306));
   AO22CHD U5088 (.O(n3663), 
	.B2(n442), 
	.B1(\ram[192][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n306));
   AO22CHD U5089 (.O(n3664), 
	.B2(n442), 
	.B1(\ram[192][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n306));
   AO22CHD U5090 (.O(n3665), 
	.B2(n442), 
	.B1(\ram[192][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n306));
   AO22CHD U5091 (.O(n3666), 
	.B2(n442), 
	.B1(\ram[192][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n306));
   AO22CHD U5092 (.O(n3667), 
	.B2(n442), 
	.B1(\ram[192][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n306));
   AO22CHD U5093 (.O(n3668), 
	.B2(n442), 
	.B1(\ram[192][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n306));
   AO22CHD U5094 (.O(n3669), 
	.B2(n442), 
	.B1(\ram[192][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n306));
   AO22CHD U5095 (.O(n3670), 
	.B2(n445), 
	.B1(\ram[193][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n308));
   AO22CHD U5096 (.O(n3671), 
	.B2(n445), 
	.B1(\ram[193][1] ), 
	.A2(n9), 
	.A1(n308));
   AO22CHD U5097 (.O(n3672), 
	.B2(n445), 
	.B1(\ram[193][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n308));
   AO22CHD U5098 (.O(n3673), 
	.B2(n445), 
	.B1(\ram[193][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n308));
   AO22CHD U5099 (.O(n3674), 
	.B2(n445), 
	.B1(\ram[193][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n308));
   AO22CHD U5100 (.O(n3675), 
	.B2(n445), 
	.B1(\ram[193][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n308));
   AO22CHD U5101 (.O(n3676), 
	.B2(n445), 
	.B1(\ram[193][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n308));
   AO22CHD U5102 (.O(n3677), 
	.B2(n445), 
	.B1(\ram[193][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n308));
   AO22CHD U5103 (.O(n3678), 
	.B2(n445), 
	.B1(\ram[193][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n308));
   AO22CHD U5104 (.O(n3679), 
	.B2(n445), 
	.B1(\ram[193][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n308));
   AO22CHD U5105 (.O(n3680), 
	.B2(n445), 
	.B1(\ram[193][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n308));
   AO22CHD U5106 (.O(n3681), 
	.B2(n445), 
	.B1(\ram[193][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n308));
   AO22CHD U5107 (.O(n3682), 
	.B2(n445), 
	.B1(\ram[193][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n308));
   AO22CHD U5108 (.O(n3683), 
	.B2(n445), 
	.B1(\ram[193][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n308));
   AO22CHD U5109 (.O(n3684), 
	.B2(n445), 
	.B1(\ram[193][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n308));
   AO22CHD U5110 (.O(n3685), 
	.B2(n445), 
	.B1(\ram[193][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n308));
   AO22CHD U5111 (.O(n3686), 
	.B2(n447), 
	.B1(\ram[194][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n310));
   AO22CHD U5112 (.O(n3687), 
	.B2(n447), 
	.B1(\ram[194][1] ), 
	.A2(n9), 
	.A1(n310));
   AO22CHD U5113 (.O(n3688), 
	.B2(n447), 
	.B1(\ram[194][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n310));
   AO22CHD U5114 (.O(n3689), 
	.B2(n447), 
	.B1(\ram[194][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n310));
   AO22CHD U5115 (.O(n3690), 
	.B2(n447), 
	.B1(\ram[194][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n310));
   AO22CHD U5116 (.O(n3691), 
	.B2(n447), 
	.B1(\ram[194][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n310));
   AO22CHD U5117 (.O(n3692), 
	.B2(n447), 
	.B1(\ram[194][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n310));
   AO22CHD U5118 (.O(n3693), 
	.B2(n447), 
	.B1(\ram[194][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n310));
   AO22CHD U5119 (.O(n3694), 
	.B2(n447), 
	.B1(\ram[194][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n310));
   AO22CHD U5120 (.O(n3695), 
	.B2(n447), 
	.B1(\ram[194][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n310));
   AO22CHD U5121 (.O(n3696), 
	.B2(n447), 
	.B1(\ram[194][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n310));
   AO22CHD U5122 (.O(n3697), 
	.B2(n447), 
	.B1(\ram[194][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n310));
   AO22CHD U5123 (.O(n3698), 
	.B2(n447), 
	.B1(\ram[194][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n310));
   AO22CHD U5124 (.O(n3699), 
	.B2(n447), 
	.B1(\ram[194][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n310));
   AO22CHD U5125 (.O(n3700), 
	.B2(n447), 
	.B1(\ram[194][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n310));
   AO22CHD U5126 (.O(n3701), 
	.B2(n447), 
	.B1(\ram[194][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n310));
   AO22CHD U5127 (.O(n3702), 
	.B2(n449), 
	.B1(\ram[195][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n311));
   AO22CHD U5128 (.O(n3703), 
	.B2(n449), 
	.B1(\ram[195][1] ), 
	.A2(n9), 
	.A1(n311));
   AO22CHD U5129 (.O(n3704), 
	.B2(n449), 
	.B1(\ram[195][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n311));
   AO22CHD U5130 (.O(n3705), 
	.B2(n449), 
	.B1(\ram[195][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n311));
   AO22CHD U5131 (.O(n3706), 
	.B2(n449), 
	.B1(\ram[195][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n311));
   AO22CHD U5132 (.O(n3707), 
	.B2(n449), 
	.B1(\ram[195][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n311));
   AO22CHD U5133 (.O(n3708), 
	.B2(n449), 
	.B1(\ram[195][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n311));
   AO22CHD U5134 (.O(n3709), 
	.B2(n449), 
	.B1(\ram[195][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n311));
   AO22CHD U5135 (.O(n3710), 
	.B2(n449), 
	.B1(\ram[195][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n311));
   AO22CHD U5136 (.O(n3711), 
	.B2(n449), 
	.B1(\ram[195][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n311));
   AO22CHD U5137 (.O(n3712), 
	.B2(n449), 
	.B1(\ram[195][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n311));
   AO22CHD U5138 (.O(n3713), 
	.B2(n449), 
	.B1(\ram[195][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n311));
   AO22CHD U5139 (.O(n3714), 
	.B2(n449), 
	.B1(\ram[195][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n311));
   AO22CHD U5140 (.O(n3715), 
	.B2(n449), 
	.B1(\ram[195][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n311));
   AO22CHD U5141 (.O(n3716), 
	.B2(n449), 
	.B1(\ram[195][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n311));
   AO22CHD U5142 (.O(n3717), 
	.B2(n449), 
	.B1(\ram[195][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n311));
   AO22CHD U5143 (.O(n3718), 
	.B2(n451), 
	.B1(\ram[196][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n313));
   AO22CHD U5144 (.O(n3719), 
	.B2(n451), 
	.B1(\ram[196][1] ), 
	.A2(n9), 
	.A1(n313));
   AO22CHD U5145 (.O(n3720), 
	.B2(n451), 
	.B1(\ram[196][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n313));
   AO22CHD U5146 (.O(n3721), 
	.B2(n451), 
	.B1(\ram[196][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n313));
   AO22CHD U5147 (.O(n3722), 
	.B2(n451), 
	.B1(\ram[196][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n313));
   AO22CHD U5148 (.O(n3723), 
	.B2(n451), 
	.B1(\ram[196][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n313));
   AO22CHD U5149 (.O(n3724), 
	.B2(n451), 
	.B1(\ram[196][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n313));
   AO22CHD U5150 (.O(n3725), 
	.B2(n451), 
	.B1(\ram[196][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n313));
   AO22CHD U5151 (.O(n3726), 
	.B2(n451), 
	.B1(\ram[196][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n313));
   AO22CHD U5152 (.O(n3727), 
	.B2(n451), 
	.B1(\ram[196][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n313));
   AO22CHD U5153 (.O(n3728), 
	.B2(n451), 
	.B1(\ram[196][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n313));
   AO22CHD U5154 (.O(n3729), 
	.B2(n451), 
	.B1(\ram[196][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n313));
   AO22CHD U5155 (.O(n3730), 
	.B2(n451), 
	.B1(\ram[196][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n313));
   AO22CHD U5156 (.O(n3731), 
	.B2(n451), 
	.B1(\ram[196][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n313));
   AO22CHD U5157 (.O(n3732), 
	.B2(n451), 
	.B1(\ram[196][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n313));
   AO22CHD U5158 (.O(n3733), 
	.B2(n451), 
	.B1(\ram[196][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n313));
   AO22CHD U5159 (.O(n3734), 
	.B2(n453), 
	.B1(\ram[197][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n315));
   AO22CHD U5160 (.O(n3735), 
	.B2(n453), 
	.B1(\ram[197][1] ), 
	.A2(n9), 
	.A1(n315));
   AO22CHD U5161 (.O(n3736), 
	.B2(n453), 
	.B1(\ram[197][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n315));
   AO22CHD U5162 (.O(n3737), 
	.B2(n453), 
	.B1(\ram[197][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n315));
   AO22CHD U5163 (.O(n3738), 
	.B2(n453), 
	.B1(\ram[197][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n315));
   AO22CHD U5164 (.O(n3739), 
	.B2(n453), 
	.B1(\ram[197][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n315));
   AO22CHD U5165 (.O(n3740), 
	.B2(n453), 
	.B1(\ram[197][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n315));
   AO22CHD U5166 (.O(n3741), 
	.B2(n453), 
	.B1(\ram[197][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n315));
   AO22CHD U5167 (.O(n3742), 
	.B2(n453), 
	.B1(\ram[197][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n315));
   AO22CHD U5168 (.O(n3743), 
	.B2(n453), 
	.B1(\ram[197][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n315));
   AO22CHD U5169 (.O(n3744), 
	.B2(n453), 
	.B1(\ram[197][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n315));
   AO22CHD U5170 (.O(n3745), 
	.B2(n453), 
	.B1(\ram[197][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n315));
   AO22CHD U5171 (.O(n3746), 
	.B2(n453), 
	.B1(\ram[197][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n315));
   AO22CHD U5172 (.O(n3747), 
	.B2(n453), 
	.B1(\ram[197][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n315));
   AO22CHD U5173 (.O(n3748), 
	.B2(n453), 
	.B1(\ram[197][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n315));
   AO22CHD U5174 (.O(n3749), 
	.B2(n453), 
	.B1(\ram[197][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n315));
   AO22CHD U5175 (.O(n3750), 
	.B2(n455), 
	.B1(\ram[198][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n317));
   AO22CHD U5176 (.O(n3751), 
	.B2(n455), 
	.B1(\ram[198][1] ), 
	.A2(n9), 
	.A1(n317));
   AO22CHD U5177 (.O(n3752), 
	.B2(n455), 
	.B1(\ram[198][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n317));
   AO22CHD U5178 (.O(n3753), 
	.B2(n455), 
	.B1(\ram[198][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n317));
   AO22CHD U5179 (.O(n3754), 
	.B2(n455), 
	.B1(\ram[198][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n317));
   AO22CHD U5180 (.O(n3755), 
	.B2(n455), 
	.B1(\ram[198][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n317));
   AO22CHD U5181 (.O(n3756), 
	.B2(n455), 
	.B1(\ram[198][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n317));
   AO22CHD U5182 (.O(n3757), 
	.B2(n455), 
	.B1(\ram[198][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n317));
   AO22CHD U5183 (.O(n3758), 
	.B2(n455), 
	.B1(\ram[198][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n317));
   AO22CHD U5184 (.O(n3759), 
	.B2(n455), 
	.B1(\ram[198][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n317));
   AO22CHD U5185 (.O(n3760), 
	.B2(n455), 
	.B1(\ram[198][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n317));
   AO22CHD U5186 (.O(n3761), 
	.B2(n455), 
	.B1(\ram[198][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n317));
   AO22CHD U5187 (.O(n3762), 
	.B2(n455), 
	.B1(\ram[198][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n317));
   AO22CHD U5188 (.O(n3763), 
	.B2(n455), 
	.B1(\ram[198][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n317));
   AO22CHD U5189 (.O(n3764), 
	.B2(n455), 
	.B1(\ram[198][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n317));
   AO22CHD U5190 (.O(n3765), 
	.B2(n455), 
	.B1(\ram[198][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n317));
   AO22CHD U5191 (.O(n3766), 
	.B2(n457), 
	.B1(\ram[199][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n319));
   AO22CHD U5192 (.O(n3767), 
	.B2(n457), 
	.B1(\ram[199][1] ), 
	.A2(n9), 
	.A1(n319));
   AO22CHD U5193 (.O(n3768), 
	.B2(n457), 
	.B1(\ram[199][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n319));
   AO22CHD U5194 (.O(n3769), 
	.B2(n457), 
	.B1(\ram[199][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n319));
   AO22CHD U5195 (.O(n3770), 
	.B2(n457), 
	.B1(\ram[199][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n319));
   AO22CHD U5196 (.O(n3771), 
	.B2(n457), 
	.B1(\ram[199][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n319));
   AO22CHD U5197 (.O(n3772), 
	.B2(n457), 
	.B1(\ram[199][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n319));
   AO22CHD U5198 (.O(n3773), 
	.B2(n457), 
	.B1(\ram[199][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n319));
   AO22CHD U5199 (.O(n3774), 
	.B2(n457), 
	.B1(\ram[199][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n319));
   AO22CHD U5200 (.O(n3775), 
	.B2(n457), 
	.B1(\ram[199][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n319));
   AO22CHD U5201 (.O(n3776), 
	.B2(n457), 
	.B1(\ram[199][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n319));
   AO22CHD U5202 (.O(n3777), 
	.B2(n457), 
	.B1(\ram[199][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n319));
   AO22CHD U5203 (.O(n3778), 
	.B2(n457), 
	.B1(\ram[199][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n319));
   AO22CHD U5204 (.O(n3779), 
	.B2(n457), 
	.B1(\ram[199][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n319));
   AO22CHD U5205 (.O(n3780), 
	.B2(n457), 
	.B1(\ram[199][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n319));
   AO22CHD U5206 (.O(n3781), 
	.B2(n457), 
	.B1(\ram[199][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n319));
   AO22CHD U5207 (.O(n3782), 
	.B2(n459), 
	.B1(\ram[200][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n321));
   AO22CHD U5208 (.O(n3783), 
	.B2(n459), 
	.B1(\ram[200][1] ), 
	.A2(n9), 
	.A1(n321));
   AO22CHD U5209 (.O(n3784), 
	.B2(n459), 
	.B1(\ram[200][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n321));
   AO22CHD U5210 (.O(n3785), 
	.B2(n459), 
	.B1(\ram[200][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n321));
   AO22CHD U5211 (.O(n3786), 
	.B2(n459), 
	.B1(\ram[200][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n321));
   AO22CHD U5212 (.O(n3787), 
	.B2(n459), 
	.B1(\ram[200][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n321));
   AO22CHD U5213 (.O(n3788), 
	.B2(n459), 
	.B1(\ram[200][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n321));
   AO22CHD U5214 (.O(n3789), 
	.B2(n459), 
	.B1(\ram[200][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n321));
   AO22CHD U5215 (.O(n3790), 
	.B2(n459), 
	.B1(\ram[200][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n321));
   AO22CHD U5216 (.O(n3791), 
	.B2(n459), 
	.B1(\ram[200][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n321));
   AO22CHD U5217 (.O(n3792), 
	.B2(n459), 
	.B1(\ram[200][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n321));
   AO22CHD U5218 (.O(n3793), 
	.B2(n459), 
	.B1(\ram[200][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n321));
   AO22CHD U5219 (.O(n3794), 
	.B2(n459), 
	.B1(\ram[200][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n321));
   AO22CHD U5220 (.O(n3795), 
	.B2(n459), 
	.B1(\ram[200][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n321));
   AO22CHD U5221 (.O(n3796), 
	.B2(n459), 
	.B1(\ram[200][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n321));
   AO22CHD U5222 (.O(n3797), 
	.B2(n459), 
	.B1(\ram[200][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n321));
   AO22CHD U5223 (.O(n3798), 
	.B2(n461), 
	.B1(\ram[201][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n323));
   AO22CHD U5224 (.O(n3799), 
	.B2(n461), 
	.B1(\ram[201][1] ), 
	.A2(n9), 
	.A1(n323));
   AO22CHD U5225 (.O(n3800), 
	.B2(n461), 
	.B1(\ram[201][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n323));
   AO22CHD U5226 (.O(n3801), 
	.B2(n461), 
	.B1(\ram[201][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n323));
   AO22CHD U5227 (.O(n3802), 
	.B2(n461), 
	.B1(\ram[201][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n323));
   AO22CHD U5228 (.O(n3803), 
	.B2(n461), 
	.B1(\ram[201][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n323));
   AO22CHD U5229 (.O(n3804), 
	.B2(n461), 
	.B1(\ram[201][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n323));
   AO22CHD U5230 (.O(n3805), 
	.B2(n461), 
	.B1(\ram[201][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n323));
   AO22CHD U5231 (.O(n3806), 
	.B2(n461), 
	.B1(\ram[201][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n323));
   AO22CHD U5232 (.O(n3807), 
	.B2(n461), 
	.B1(\ram[201][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n323));
   AO22CHD U5233 (.O(n3808), 
	.B2(n461), 
	.B1(\ram[201][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n323));
   AO22CHD U5234 (.O(n3809), 
	.B2(n461), 
	.B1(\ram[201][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n323));
   AO22CHD U5235 (.O(n3810), 
	.B2(n461), 
	.B1(\ram[201][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n323));
   AO22CHD U5236 (.O(n3811), 
	.B2(n461), 
	.B1(\ram[201][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n323));
   AO22CHD U5237 (.O(n3812), 
	.B2(n461), 
	.B1(\ram[201][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n323));
   AO22CHD U5238 (.O(n3813), 
	.B2(n461), 
	.B1(\ram[201][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n323));
   AO22CHD U5239 (.O(n3814), 
	.B2(n463), 
	.B1(\ram[202][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n325));
   AO22CHD U5240 (.O(n3815), 
	.B2(n463), 
	.B1(\ram[202][1] ), 
	.A2(n9), 
	.A1(n325));
   AO22CHD U5241 (.O(n3816), 
	.B2(n463), 
	.B1(\ram[202][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n325));
   AO22CHD U5242 (.O(n3817), 
	.B2(n463), 
	.B1(\ram[202][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n325));
   AO22CHD U5243 (.O(n3818), 
	.B2(n463), 
	.B1(\ram[202][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n325));
   AO22CHD U5244 (.O(n3819), 
	.B2(n463), 
	.B1(\ram[202][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n325));
   AO22CHD U5245 (.O(n3820), 
	.B2(n463), 
	.B1(\ram[202][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n325));
   AO22CHD U5246 (.O(n3821), 
	.B2(n463), 
	.B1(\ram[202][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n325));
   AO22CHD U5247 (.O(n3822), 
	.B2(n463), 
	.B1(\ram[202][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n325));
   AO22CHD U5248 (.O(n3823), 
	.B2(n463), 
	.B1(\ram[202][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n325));
   AO22CHD U5249 (.O(n3824), 
	.B2(n463), 
	.B1(\ram[202][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n325));
   AO22CHD U5250 (.O(n3825), 
	.B2(n463), 
	.B1(\ram[202][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n325));
   AO22CHD U5251 (.O(n3826), 
	.B2(n463), 
	.B1(\ram[202][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n325));
   AO22CHD U5252 (.O(n3827), 
	.B2(n463), 
	.B1(\ram[202][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n325));
   AO22CHD U5253 (.O(n3828), 
	.B2(n463), 
	.B1(\ram[202][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n325));
   AO22CHD U5254 (.O(n3829), 
	.B2(n463), 
	.B1(\ram[202][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n325));
   AO22CHD U5255 (.O(n3830), 
	.B2(n465), 
	.B1(\ram[203][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n327));
   AO22CHD U5256 (.O(n3831), 
	.B2(n465), 
	.B1(\ram[203][1] ), 
	.A2(n9), 
	.A1(n327));
   AO22CHD U5257 (.O(n3832), 
	.B2(n465), 
	.B1(\ram[203][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n327));
   AO22CHD U5258 (.O(n3833), 
	.B2(n465), 
	.B1(\ram[203][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n327));
   AO22CHD U5259 (.O(n3834), 
	.B2(n465), 
	.B1(\ram[203][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n327));
   AO22CHD U5260 (.O(n3835), 
	.B2(n465), 
	.B1(\ram[203][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n327));
   AO22CHD U5261 (.O(n3836), 
	.B2(n465), 
	.B1(\ram[203][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n327));
   AO22CHD U5262 (.O(n3837), 
	.B2(n465), 
	.B1(\ram[203][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n327));
   AO22CHD U5263 (.O(n3838), 
	.B2(n465), 
	.B1(\ram[203][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n327));
   AO22CHD U5264 (.O(n3839), 
	.B2(n465), 
	.B1(\ram[203][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n327));
   AO22CHD U5265 (.O(n3840), 
	.B2(n465), 
	.B1(\ram[203][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n327));
   AO22CHD U5266 (.O(n3841), 
	.B2(n465), 
	.B1(\ram[203][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n327));
   AO22CHD U5267 (.O(n3842), 
	.B2(n465), 
	.B1(\ram[203][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n327));
   AO22CHD U5268 (.O(n3843), 
	.B2(n465), 
	.B1(\ram[203][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n327));
   AO22CHD U5269 (.O(n3844), 
	.B2(n465), 
	.B1(\ram[203][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n327));
   AO22CHD U5270 (.O(n3845), 
	.B2(n465), 
	.B1(\ram[203][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n327));
   AO22CHD U5271 (.O(n3846), 
	.B2(n467), 
	.B1(\ram[204][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n329));
   AO22CHD U5272 (.O(n3847), 
	.B2(n467), 
	.B1(\ram[204][1] ), 
	.A2(n9), 
	.A1(n329));
   AO22CHD U5273 (.O(n3848), 
	.B2(n467), 
	.B1(\ram[204][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n329));
   AO22CHD U5274 (.O(n3849), 
	.B2(n467), 
	.B1(\ram[204][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n329));
   AO22CHD U5275 (.O(n3850), 
	.B2(n467), 
	.B1(\ram[204][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n329));
   AO22CHD U5276 (.O(n3851), 
	.B2(n467), 
	.B1(\ram[204][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n329));
   AO22CHD U5277 (.O(n3852), 
	.B2(n467), 
	.B1(\ram[204][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n329));
   AO22CHD U5278 (.O(n3853), 
	.B2(n467), 
	.B1(\ram[204][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n329));
   AO22CHD U5279 (.O(n3854), 
	.B2(n467), 
	.B1(\ram[204][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n329));
   AO22CHD U5280 (.O(n3855), 
	.B2(n467), 
	.B1(\ram[204][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n329));
   AO22CHD U5281 (.O(n3856), 
	.B2(n467), 
	.B1(\ram[204][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n329));
   AO22CHD U5282 (.O(n3857), 
	.B2(n467), 
	.B1(\ram[204][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n329));
   AO22CHD U5283 (.O(n3858), 
	.B2(n467), 
	.B1(\ram[204][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n329));
   AO22CHD U5284 (.O(n3859), 
	.B2(n467), 
	.B1(\ram[204][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n329));
   AO22CHD U5285 (.O(n3860), 
	.B2(n467), 
	.B1(\ram[204][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n329));
   AO22CHD U5286 (.O(n3861), 
	.B2(n467), 
	.B1(\ram[204][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n329));
   AO22CHD U5287 (.O(n3862), 
	.B2(n469), 
	.B1(\ram[205][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n331));
   AO22CHD U5288 (.O(n3863), 
	.B2(n469), 
	.B1(\ram[205][1] ), 
	.A2(n9), 
	.A1(n331));
   AO22CHD U5289 (.O(n3864), 
	.B2(n469), 
	.B1(\ram[205][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n331));
   AO22CHD U5290 (.O(n3865), 
	.B2(n469), 
	.B1(\ram[205][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n331));
   AO22CHD U5291 (.O(n3866), 
	.B2(n469), 
	.B1(\ram[205][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n331));
   AO22CHD U5292 (.O(n3867), 
	.B2(n469), 
	.B1(\ram[205][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n331));
   AO22CHD U5293 (.O(n3868), 
	.B2(n469), 
	.B1(\ram[205][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n331));
   AO22CHD U5294 (.O(n3869), 
	.B2(n469), 
	.B1(\ram[205][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n331));
   AO22CHD U5295 (.O(n3870), 
	.B2(n469), 
	.B1(\ram[205][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n331));
   AO22CHD U5296 (.O(n3871), 
	.B2(n469), 
	.B1(\ram[205][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n331));
   AO22CHD U5297 (.O(n3872), 
	.B2(n469), 
	.B1(\ram[205][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n331));
   AO22CHD U5298 (.O(n3873), 
	.B2(n469), 
	.B1(\ram[205][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n331));
   AO22CHD U5299 (.O(n3874), 
	.B2(n469), 
	.B1(\ram[205][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n331));
   AO22CHD U5300 (.O(n3875), 
	.B2(n469), 
	.B1(\ram[205][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n331));
   AO22CHD U5301 (.O(n3876), 
	.B2(n469), 
	.B1(\ram[205][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n331));
   AO22CHD U5302 (.O(n3877), 
	.B2(n469), 
	.B1(\ram[205][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n331));
   AO22CHD U5303 (.O(n3878), 
	.B2(n471), 
	.B1(\ram[206][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n333));
   AO22CHD U5304 (.O(n3879), 
	.B2(n471), 
	.B1(\ram[206][1] ), 
	.A2(n9), 
	.A1(n333));
   AO22CHD U5305 (.O(n3880), 
	.B2(n471), 
	.B1(\ram[206][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n333));
   AO22CHD U5306 (.O(n3881), 
	.B2(n471), 
	.B1(\ram[206][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n333));
   AO22CHD U5307 (.O(n3882), 
	.B2(n471), 
	.B1(\ram[206][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n333));
   AO22CHD U5308 (.O(n3883), 
	.B2(n471), 
	.B1(\ram[206][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n333));
   AO22CHD U5309 (.O(n3884), 
	.B2(n471), 
	.B1(\ram[206][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n333));
   AO22CHD U5310 (.O(n3885), 
	.B2(n471), 
	.B1(\ram[206][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n333));
   AO22CHD U5311 (.O(n3886), 
	.B2(n471), 
	.B1(\ram[206][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n333));
   AO22CHD U5312 (.O(n3887), 
	.B2(n471), 
	.B1(\ram[206][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n333));
   AO22CHD U5313 (.O(n3888), 
	.B2(n471), 
	.B1(\ram[206][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n333));
   AO22CHD U5314 (.O(n3889), 
	.B2(n471), 
	.B1(\ram[206][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n333));
   AO22CHD U5315 (.O(n3890), 
	.B2(n471), 
	.B1(\ram[206][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n333));
   AO22CHD U5316 (.O(n3891), 
	.B2(n471), 
	.B1(\ram[206][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n333));
   AO22CHD U5317 (.O(n3892), 
	.B2(n471), 
	.B1(\ram[206][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n333));
   AO22CHD U5318 (.O(n3893), 
	.B2(n471), 
	.B1(\ram[206][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n333));
   AO22CHD U5319 (.O(n3894), 
	.B2(n473), 
	.B1(\ram[207][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n335));
   AO22CHD U5320 (.O(n3895), 
	.B2(n473), 
	.B1(\ram[207][1] ), 
	.A2(n9), 
	.A1(n335));
   AO22CHD U5321 (.O(n3896), 
	.B2(n473), 
	.B1(\ram[207][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n335));
   AO22CHD U5322 (.O(n3897), 
	.B2(n473), 
	.B1(\ram[207][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n335));
   AO22CHD U5323 (.O(n3898), 
	.B2(n473), 
	.B1(\ram[207][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n335));
   AO22CHD U5324 (.O(n3899), 
	.B2(n473), 
	.B1(\ram[207][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n335));
   AO22CHD U5325 (.O(n3900), 
	.B2(n473), 
	.B1(\ram[207][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n335));
   AO22CHD U5326 (.O(n3901), 
	.B2(n473), 
	.B1(\ram[207][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n335));
   AO22CHD U5327 (.O(n3902), 
	.B2(n473), 
	.B1(\ram[207][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n335));
   AO22CHD U5328 (.O(n3903), 
	.B2(n473), 
	.B1(\ram[207][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n335));
   AO22CHD U5329 (.O(n3904), 
	.B2(n473), 
	.B1(\ram[207][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n335));
   AO22CHD U5330 (.O(n3905), 
	.B2(n473), 
	.B1(\ram[207][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n335));
   AO22CHD U5331 (.O(n3906), 
	.B2(n473), 
	.B1(\ram[207][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n335));
   AO22CHD U5332 (.O(n3907), 
	.B2(n473), 
	.B1(\ram[207][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n335));
   AO22CHD U5333 (.O(n3908), 
	.B2(n473), 
	.B1(\ram[207][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n335));
   AO22CHD U5334 (.O(n3909), 
	.B2(n473), 
	.B1(\ram[207][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n335));
   AO22CHD U5335 (.O(n3910), 
	.B2(n476), 
	.B1(\ram[208][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n337));
   AO22CHD U5336 (.O(n3911), 
	.B2(n476), 
	.B1(\ram[208][1] ), 
	.A2(n9), 
	.A1(n337));
   AO22CHD U5337 (.O(n3912), 
	.B2(n476), 
	.B1(\ram[208][2] ), 
	.A2(n10), 
	.A1(n337));
   AO22CHD U5338 (.O(n3913), 
	.B2(n476), 
	.B1(\ram[208][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n337));
   AO22CHD U5339 (.O(n3914), 
	.B2(n476), 
	.B1(\ram[208][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n337));
   AO22CHD U5340 (.O(n3915), 
	.B2(n476), 
	.B1(\ram[208][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n337));
   AO22CHD U5341 (.O(n3916), 
	.B2(n476), 
	.B1(\ram[208][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n337));
   AO22CHD U5342 (.O(n3917), 
	.B2(n476), 
	.B1(\ram[208][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n337));
   AO22CHD U5343 (.O(n3918), 
	.B2(n476), 
	.B1(\ram[208][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n337));
   AO22CHD U5344 (.O(n3919), 
	.B2(n476), 
	.B1(\ram[208][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n337));
   AO22CHD U5345 (.O(n3920), 
	.B2(n476), 
	.B1(\ram[208][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n337));
   AO22CHD U5346 (.O(n3921), 
	.B2(n476), 
	.B1(\ram[208][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n337));
   AO22CHD U5347 (.O(n3922), 
	.B2(n476), 
	.B1(\ram[208][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n337));
   AO22CHD U5348 (.O(n3923), 
	.B2(n476), 
	.B1(\ram[208][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n337));
   AO22CHD U5349 (.O(n3924), 
	.B2(n476), 
	.B1(\ram[208][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n337));
   AO22CHD U5350 (.O(n3925), 
	.B2(n476), 
	.B1(\ram[208][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n337));
   AO22CHD U5351 (.O(n3926), 
	.B2(n479), 
	.B1(\ram[209][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n339));
   AO22CHD U5352 (.O(n3927), 
	.B2(n479), 
	.B1(\ram[209][1] ), 
	.A2(n9), 
	.A1(n339));
   AO22CHD U5353 (.O(n3928), 
	.B2(n479), 
	.B1(\ram[209][2] ), 
	.A2(n10), 
	.A1(n339));
   AO22CHD U5354 (.O(n3929), 
	.B2(n479), 
	.B1(\ram[209][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n339));
   AO22CHD U5355 (.O(n3930), 
	.B2(n479), 
	.B1(\ram[209][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n339));
   AO22CHD U5356 (.O(n3931), 
	.B2(n479), 
	.B1(\ram[209][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n339));
   AO22CHD U5357 (.O(n3932), 
	.B2(n479), 
	.B1(\ram[209][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n339));
   AO22CHD U5358 (.O(n3933), 
	.B2(n479), 
	.B1(\ram[209][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n339));
   AO22CHD U5359 (.O(n3934), 
	.B2(n479), 
	.B1(\ram[209][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n339));
   AO22CHD U5360 (.O(n3935), 
	.B2(n479), 
	.B1(\ram[209][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n339));
   AO22CHD U5361 (.O(n3936), 
	.B2(n479), 
	.B1(\ram[209][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n339));
   AO22CHD U5362 (.O(n3937), 
	.B2(n479), 
	.B1(\ram[209][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n339));
   AO22CHD U5363 (.O(n3938), 
	.B2(n479), 
	.B1(\ram[209][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n339));
   AO22CHD U5364 (.O(n3939), 
	.B2(n479), 
	.B1(\ram[209][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n339));
   AO22CHD U5365 (.O(n3940), 
	.B2(n479), 
	.B1(\ram[209][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n339));
   AO22CHD U5366 (.O(n3941), 
	.B2(n479), 
	.B1(\ram[209][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n339));
   AO22CHD U5367 (.O(n3942), 
	.B2(n481), 
	.B1(\ram[210][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n342));
   AO22CHD U5368 (.O(n3943), 
	.B2(n481), 
	.B1(\ram[210][1] ), 
	.A2(n9), 
	.A1(n342));
   AO22CHD U5369 (.O(n3944), 
	.B2(n481), 
	.B1(\ram[210][2] ), 
	.A2(n10), 
	.A1(n342));
   AO22CHD U5370 (.O(n3945), 
	.B2(n481), 
	.B1(\ram[210][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n342));
   AO22CHD U5371 (.O(n3946), 
	.B2(n481), 
	.B1(\ram[210][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n342));
   AO22CHD U5372 (.O(n3947), 
	.B2(n481), 
	.B1(\ram[210][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n342));
   AO22CHD U5373 (.O(n3948), 
	.B2(n481), 
	.B1(\ram[210][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n342));
   AO22CHD U5374 (.O(n3949), 
	.B2(n481), 
	.B1(\ram[210][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n342));
   AO22CHD U5375 (.O(n3950), 
	.B2(n481), 
	.B1(\ram[210][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n342));
   AO22CHD U5376 (.O(n3951), 
	.B2(n481), 
	.B1(\ram[210][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n342));
   AO22CHD U5377 (.O(n3952), 
	.B2(n481), 
	.B1(\ram[210][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n342));
   AO22CHD U5378 (.O(n3953), 
	.B2(n481), 
	.B1(\ram[210][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n342));
   AO22CHD U5379 (.O(n3954), 
	.B2(n481), 
	.B1(\ram[210][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n342));
   AO22CHD U5380 (.O(n3955), 
	.B2(n481), 
	.B1(\ram[210][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n342));
   AO22CHD U5381 (.O(n3956), 
	.B2(n481), 
	.B1(\ram[210][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n342));
   AO22CHD U5382 (.O(n3957), 
	.B2(n481), 
	.B1(\ram[210][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n342));
   AO22CHD U5383 (.O(n3958), 
	.B2(n483), 
	.B1(\ram[211][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n344));
   AO22CHD U5384 (.O(n3959), 
	.B2(n483), 
	.B1(\ram[211][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n344));
   AO22CHD U5385 (.O(n3960), 
	.B2(n483), 
	.B1(\ram[211][2] ), 
	.A2(n10), 
	.A1(n344));
   AO22CHD U5386 (.O(n3961), 
	.B2(n483), 
	.B1(\ram[211][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n344));
   AO22CHD U5387 (.O(n3962), 
	.B2(n483), 
	.B1(\ram[211][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n344));
   AO22CHD U5388 (.O(n3963), 
	.B2(n483), 
	.B1(\ram[211][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n344));
   AO22CHD U5389 (.O(n3964), 
	.B2(n483), 
	.B1(\ram[211][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n344));
   AO22CHD U5390 (.O(n3965), 
	.B2(n483), 
	.B1(\ram[211][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n344));
   AO22CHD U5391 (.O(n3966), 
	.B2(n483), 
	.B1(\ram[211][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n344));
   AO22CHD U5392 (.O(n3967), 
	.B2(n483), 
	.B1(\ram[211][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n344));
   AO22CHD U5393 (.O(n3968), 
	.B2(n483), 
	.B1(\ram[211][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n344));
   AO22CHD U5394 (.O(n3969), 
	.B2(n483), 
	.B1(\ram[211][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n344));
   AO22CHD U5395 (.O(n3970), 
	.B2(n483), 
	.B1(\ram[211][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n344));
   AO22CHD U5396 (.O(n3971), 
	.B2(n483), 
	.B1(\ram[211][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n344));
   AO22CHD U5397 (.O(n3972), 
	.B2(n483), 
	.B1(\ram[211][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n344));
   AO22CHD U5398 (.O(n3973), 
	.B2(n483), 
	.B1(\ram[211][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n344));
   AO22CHD U5399 (.O(n3974), 
	.B2(n485), 
	.B1(\ram[212][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n345));
   AO22CHD U5400 (.O(n3975), 
	.B2(n485), 
	.B1(\ram[212][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n345));
   AO22CHD U5401 (.O(n3976), 
	.B2(n485), 
	.B1(\ram[212][2] ), 
	.A2(n10), 
	.A1(n345));
   AO22CHD U5402 (.O(n3977), 
	.B2(n485), 
	.B1(\ram[212][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n345));
   AO22CHD U5403 (.O(n3978), 
	.B2(n485), 
	.B1(\ram[212][4] ), 
	.A2(n12), 
	.A1(n345));
   AO22CHD U5404 (.O(n3979), 
	.B2(n485), 
	.B1(\ram[212][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n345));
   AO22CHD U5405 (.O(n3980), 
	.B2(n485), 
	.B1(\ram[212][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n345));
   AO22CHD U5406 (.O(n3981), 
	.B2(n485), 
	.B1(\ram[212][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n345));
   AO22CHD U5407 (.O(n3982), 
	.B2(n485), 
	.B1(\ram[212][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n345));
   AO22CHD U5408 (.O(n3983), 
	.B2(n485), 
	.B1(\ram[212][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n345));
   AO22CHD U5409 (.O(n3984), 
	.B2(n485), 
	.B1(\ram[212][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n345));
   AO22CHD U5410 (.O(n3985), 
	.B2(n485), 
	.B1(\ram[212][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n345));
   AO22CHD U5411 (.O(n3986), 
	.B2(n485), 
	.B1(\ram[212][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n345));
   AO22CHD U5412 (.O(n3987), 
	.B2(n485), 
	.B1(\ram[212][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n345));
   AO22CHD U5413 (.O(n3988), 
	.B2(n485), 
	.B1(\ram[212][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n345));
   AO22CHD U5414 (.O(n3989), 
	.B2(n485), 
	.B1(\ram[212][15] ), 
	.A2(n23), 
	.A1(n345));
   AO22CHD U5415 (.O(n3990), 
	.B2(n487), 
	.B1(\ram[213][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n347));
   AO22CHD U5416 (.O(n3991), 
	.B2(n487), 
	.B1(\ram[213][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n347));
   AO22CHD U5417 (.O(n3992), 
	.B2(n487), 
	.B1(\ram[213][2] ), 
	.A2(n10), 
	.A1(n347));
   AO22CHD U5418 (.O(n3993), 
	.B2(n487), 
	.B1(\ram[213][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n347));
   AO22CHD U5419 (.O(n3994), 
	.B2(n487), 
	.B1(\ram[213][4] ), 
	.A2(n12), 
	.A1(n347));
   AO22CHD U5420 (.O(n3995), 
	.B2(n487), 
	.B1(\ram[213][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n347));
   AO22CHD U5421 (.O(n3996), 
	.B2(n487), 
	.B1(\ram[213][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n347));
   AO22CHD U5422 (.O(n3997), 
	.B2(n487), 
	.B1(\ram[213][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n347));
   AO22CHD U5423 (.O(n3998), 
	.B2(n487), 
	.B1(\ram[213][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n347));
   AO22CHD U5424 (.O(n3999), 
	.B2(n487), 
	.B1(\ram[213][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n347));
   AO22CHD U5425 (.O(n4000), 
	.B2(n487), 
	.B1(\ram[213][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n347));
   AO22CHD U5426 (.O(n4001), 
	.B2(n487), 
	.B1(\ram[213][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n347));
   AO22CHD U5427 (.O(n4002), 
	.B2(n487), 
	.B1(\ram[213][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n347));
   AO22CHD U5428 (.O(n4003), 
	.B2(n487), 
	.B1(\ram[213][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n347));
   AO22CHD U5429 (.O(n4004), 
	.B2(n487), 
	.B1(\ram[213][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n347));
   AO22CHD U5430 (.O(n4005), 
	.B2(n487), 
	.B1(\ram[213][15] ), 
	.A2(n23), 
	.A1(n347));
   AO22CHD U5431 (.O(n4006), 
	.B2(n489), 
	.B1(\ram[214][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n349));
   AO22CHD U5432 (.O(n4007), 
	.B2(n489), 
	.B1(\ram[214][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n349));
   AO22CHD U5433 (.O(n4008), 
	.B2(n489), 
	.B1(\ram[214][2] ), 
	.A2(n10), 
	.A1(n349));
   AO22CHD U5434 (.O(n4009), 
	.B2(n489), 
	.B1(\ram[214][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n349));
   AO22CHD U5435 (.O(n4010), 
	.B2(n489), 
	.B1(\ram[214][4] ), 
	.A2(n12), 
	.A1(n349));
   AO22CHD U5436 (.O(n4011), 
	.B2(n489), 
	.B1(\ram[214][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n349));
   AO22CHD U5437 (.O(n4012), 
	.B2(n489), 
	.B1(\ram[214][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n349));
   AO22CHD U5438 (.O(n4013), 
	.B2(n489), 
	.B1(\ram[214][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n349));
   AO22CHD U5439 (.O(n4014), 
	.B2(n489), 
	.B1(\ram[214][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n349));
   AO22CHD U5440 (.O(n4015), 
	.B2(n489), 
	.B1(\ram[214][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n349));
   AO22CHD U5441 (.O(n4016), 
	.B2(n489), 
	.B1(\ram[214][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n349));
   AO22CHD U5442 (.O(n4017), 
	.B2(n489), 
	.B1(\ram[214][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n349));
   AO22CHD U5443 (.O(n4018), 
	.B2(n489), 
	.B1(\ram[214][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n349));
   AO22CHD U5444 (.O(n4019), 
	.B2(n489), 
	.B1(\ram[214][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n349));
   AO22CHD U5445 (.O(n4020), 
	.B2(n489), 
	.B1(\ram[214][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n349));
   AO22CHD U5446 (.O(n4021), 
	.B2(n489), 
	.B1(\ram[214][15] ), 
	.A2(n23), 
	.A1(n349));
   AO22CHD U5447 (.O(n4022), 
	.B2(n491), 
	.B1(\ram[215][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n351));
   AO22CHD U5448 (.O(n4023), 
	.B2(n491), 
	.B1(\ram[215][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n351));
   AO22CHD U5449 (.O(n4024), 
	.B2(n491), 
	.B1(\ram[215][2] ), 
	.A2(n10), 
	.A1(n351));
   AO22CHD U5450 (.O(n4025), 
	.B2(n491), 
	.B1(\ram[215][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n351));
   AO22CHD U5451 (.O(n4026), 
	.B2(n491), 
	.B1(\ram[215][4] ), 
	.A2(n12), 
	.A1(n351));
   AO22CHD U5452 (.O(n4027), 
	.B2(n491), 
	.B1(\ram[215][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n351));
   AO22CHD U5453 (.O(n4028), 
	.B2(n491), 
	.B1(\ram[215][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n351));
   AO22CHD U5454 (.O(n4029), 
	.B2(n491), 
	.B1(\ram[215][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n351));
   AO22CHD U5455 (.O(n4030), 
	.B2(n491), 
	.B1(\ram[215][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n351));
   AO22CHD U5456 (.O(n4031), 
	.B2(n491), 
	.B1(\ram[215][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n351));
   AO22CHD U5457 (.O(n4032), 
	.B2(n491), 
	.B1(\ram[215][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n351));
   AO22CHD U5458 (.O(n4033), 
	.B2(n491), 
	.B1(\ram[215][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n351));
   AO22CHD U5459 (.O(n4034), 
	.B2(n491), 
	.B1(\ram[215][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n351));
   AO22CHD U5460 (.O(n4035), 
	.B2(n491), 
	.B1(\ram[215][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n351));
   AO22CHD U5461 (.O(n4036), 
	.B2(n491), 
	.B1(\ram[215][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n351));
   AO22CHD U5462 (.O(n4037), 
	.B2(n491), 
	.B1(\ram[215][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n351));
   AO22CHD U5463 (.O(n4038), 
	.B2(n493), 
	.B1(\ram[216][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n353));
   AO22CHD U5464 (.O(n4039), 
	.B2(n493), 
	.B1(\ram[216][1] ), 
	.A2(n9), 
	.A1(n353));
   AO22CHD U5465 (.O(n4040), 
	.B2(n493), 
	.B1(\ram[216][2] ), 
	.A2(n10), 
	.A1(n353));
   AO22CHD U5466 (.O(n4041), 
	.B2(n493), 
	.B1(\ram[216][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n353));
   AO22CHD U5467 (.O(n4042), 
	.B2(n493), 
	.B1(\ram[216][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n353));
   AO22CHD U5468 (.O(n4043), 
	.B2(n493), 
	.B1(\ram[216][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n353));
   AO22CHD U5469 (.O(n4044), 
	.B2(n493), 
	.B1(\ram[216][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n353));
   AO22CHD U5470 (.O(n4045), 
	.B2(n493), 
	.B1(\ram[216][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n353));
   AO22CHD U5471 (.O(n4046), 
	.B2(n493), 
	.B1(\ram[216][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n353));
   AO22CHD U5472 (.O(n4047), 
	.B2(n493), 
	.B1(\ram[216][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n353));
   AO22CHD U5473 (.O(n4048), 
	.B2(n493), 
	.B1(\ram[216][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n353));
   AO22CHD U5474 (.O(n4049), 
	.B2(n493), 
	.B1(\ram[216][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n353));
   AO22CHD U5475 (.O(n4050), 
	.B2(n493), 
	.B1(\ram[216][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n353));
   AO22CHD U5476 (.O(n4051), 
	.B2(n493), 
	.B1(\ram[216][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n353));
   AO22CHD U5477 (.O(n4052), 
	.B2(n493), 
	.B1(\ram[216][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n353));
   AO22CHD U5478 (.O(n4053), 
	.B2(n493), 
	.B1(\ram[216][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n353));
   AO22CHD U5479 (.O(n4054), 
	.B2(n495), 
	.B1(\ram[217][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n355));
   AO22CHD U5480 (.O(n4055), 
	.B2(n495), 
	.B1(\ram[217][1] ), 
	.A2(n9), 
	.A1(n355));
   AO22CHD U5481 (.O(n4056), 
	.B2(n495), 
	.B1(\ram[217][2] ), 
	.A2(n10), 
	.A1(n355));
   AO22CHD U5482 (.O(n4057), 
	.B2(n495), 
	.B1(\ram[217][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n355));
   AO22CHD U5483 (.O(n4058), 
	.B2(n495), 
	.B1(\ram[217][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n355));
   AO22CHD U5484 (.O(n4059), 
	.B2(n495), 
	.B1(\ram[217][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n355));
   AO22CHD U5485 (.O(n4060), 
	.B2(n495), 
	.B1(\ram[217][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n355));
   AO22CHD U5486 (.O(n4061), 
	.B2(n495), 
	.B1(\ram[217][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n355));
   AO22CHD U5487 (.O(n4062), 
	.B2(n495), 
	.B1(\ram[217][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n355));
   AO22CHD U5488 (.O(n4063), 
	.B2(n495), 
	.B1(\ram[217][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n355));
   AO22CHD U5489 (.O(n4064), 
	.B2(n495), 
	.B1(\ram[217][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n355));
   AO22CHD U5490 (.O(n4065), 
	.B2(n495), 
	.B1(\ram[217][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n355));
   AO22CHD U5491 (.O(n4066), 
	.B2(n495), 
	.B1(\ram[217][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n355));
   AO22CHD U5492 (.O(n4067), 
	.B2(n495), 
	.B1(\ram[217][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n355));
   AO22CHD U5493 (.O(n4068), 
	.B2(n495), 
	.B1(\ram[217][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n355));
   AO22CHD U5494 (.O(n4069), 
	.B2(n495), 
	.B1(\ram[217][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n355));
   AO22CHD U5495 (.O(n4070), 
	.B2(n497), 
	.B1(\ram[218][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n357));
   AO22CHD U5496 (.O(n4071), 
	.B2(n497), 
	.B1(\ram[218][1] ), 
	.A2(n9), 
	.A1(n357));
   AO22CHD U5497 (.O(n4072), 
	.B2(n497), 
	.B1(\ram[218][2] ), 
	.A2(n10), 
	.A1(n357));
   AO22CHD U5498 (.O(n4073), 
	.B2(n497), 
	.B1(\ram[218][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n357));
   AO22CHD U5499 (.O(n4074), 
	.B2(n497), 
	.B1(\ram[218][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n357));
   AO22CHD U5500 (.O(n4075), 
	.B2(n497), 
	.B1(\ram[218][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n357));
   AO22CHD U5501 (.O(n4076), 
	.B2(n497), 
	.B1(\ram[218][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n357));
   AO22CHD U5502 (.O(n4077), 
	.B2(n497), 
	.B1(\ram[218][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n357));
   AO22CHD U5503 (.O(n4078), 
	.B2(n497), 
	.B1(\ram[218][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n357));
   AO22CHD U5504 (.O(n4079), 
	.B2(n497), 
	.B1(\ram[218][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n357));
   AO22CHD U5505 (.O(n4080), 
	.B2(n497), 
	.B1(\ram[218][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n357));
   AO22CHD U5506 (.O(n4081), 
	.B2(n497), 
	.B1(\ram[218][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n357));
   AO22CHD U5507 (.O(n4082), 
	.B2(n497), 
	.B1(\ram[218][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n357));
   AO22CHD U5508 (.O(n4083), 
	.B2(n497), 
	.B1(\ram[218][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n357));
   AO22CHD U5509 (.O(n4084), 
	.B2(n497), 
	.B1(\ram[218][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n357));
   AO22CHD U5510 (.O(n4085), 
	.B2(n497), 
	.B1(\ram[218][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n357));
   AO22CHD U5511 (.O(n4086), 
	.B2(n499), 
	.B1(\ram[219][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n359));
   AO22CHD U5512 (.O(n4087), 
	.B2(n499), 
	.B1(\ram[219][1] ), 
	.A2(n9), 
	.A1(n359));
   AO22CHD U5513 (.O(n4088), 
	.B2(n499), 
	.B1(\ram[219][2] ), 
	.A2(n10), 
	.A1(n359));
   AO22CHD U5514 (.O(n4089), 
	.B2(n499), 
	.B1(\ram[219][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n359));
   AO22CHD U5515 (.O(n4090), 
	.B2(n499), 
	.B1(\ram[219][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n359));
   AO22CHD U5516 (.O(n4091), 
	.B2(n499), 
	.B1(\ram[219][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n359));
   AO22CHD U5517 (.O(n4092), 
	.B2(n499), 
	.B1(\ram[219][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n359));
   AO22CHD U5518 (.O(n4093), 
	.B2(n499), 
	.B1(\ram[219][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n359));
   AO22CHD U5519 (.O(n4094), 
	.B2(n499), 
	.B1(\ram[219][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n359));
   AO22CHD U5520 (.O(n4095), 
	.B2(n499), 
	.B1(\ram[219][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n359));
   AO22CHD U5521 (.O(n4096), 
	.B2(n499), 
	.B1(\ram[219][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n359));
   AO22CHD U5522 (.O(n4097), 
	.B2(n499), 
	.B1(\ram[219][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n359));
   AO22CHD U5523 (.O(n4098), 
	.B2(n499), 
	.B1(\ram[219][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n359));
   AO22CHD U5524 (.O(n4099), 
	.B2(n499), 
	.B1(\ram[219][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n359));
   AO22CHD U5525 (.O(n4100), 
	.B2(n499), 
	.B1(\ram[219][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n359));
   AO22CHD U5526 (.O(n4101), 
	.B2(n499), 
	.B1(\ram[219][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n359));
   AO22CHD U5527 (.O(n4102), 
	.B2(n501), 
	.B1(\ram[220][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n361));
   AO22CHD U5528 (.O(n4103), 
	.B2(n501), 
	.B1(\ram[220][1] ), 
	.A2(n9), 
	.A1(n361));
   AO22CHD U5529 (.O(n4104), 
	.B2(n501), 
	.B1(\ram[220][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n361));
   AO22CHD U5530 (.O(n4105), 
	.B2(n501), 
	.B1(\ram[220][3] ), 
	.A2(n11), 
	.A1(n361));
   AO22CHD U5531 (.O(n4106), 
	.B2(n501), 
	.B1(\ram[220][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n361));
   AO22CHD U5532 (.O(n4107), 
	.B2(n501), 
	.B1(\ram[220][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n361));
   AO22CHD U5533 (.O(n4108), 
	.B2(n501), 
	.B1(\ram[220][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n361));
   AO22CHD U5534 (.O(n4109), 
	.B2(n501), 
	.B1(\ram[220][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n361));
   AO22CHD U5535 (.O(n4110), 
	.B2(n501), 
	.B1(\ram[220][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n361));
   AO22CHD U5536 (.O(n4111), 
	.B2(n501), 
	.B1(\ram[220][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n361));
   AO22CHD U5537 (.O(n4112), 
	.B2(n501), 
	.B1(\ram[220][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n361));
   AO22CHD U5538 (.O(n4113), 
	.B2(n501), 
	.B1(\ram[220][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n361));
   AO22CHD U5539 (.O(n4114), 
	.B2(n501), 
	.B1(\ram[220][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n361));
   AO22CHD U5540 (.O(n4115), 
	.B2(n501), 
	.B1(\ram[220][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n361));
   AO22CHD U5541 (.O(n4116), 
	.B2(n501), 
	.B1(\ram[220][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n361));
   AO22CHD U5542 (.O(n4117), 
	.B2(n501), 
	.B1(\ram[220][15] ), 
	.A2(n23), 
	.A1(n361));
   AO22CHD U5543 (.O(n4118), 
	.B2(n503), 
	.B1(\ram[221][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n363));
   AO22CHD U5544 (.O(n4119), 
	.B2(n503), 
	.B1(\ram[221][1] ), 
	.A2(n9), 
	.A1(n363));
   AO22CHD U5545 (.O(n4120), 
	.B2(n503), 
	.B1(\ram[221][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n363));
   AO22CHD U5546 (.O(n4121), 
	.B2(n503), 
	.B1(\ram[221][3] ), 
	.A2(n11), 
	.A1(n363));
   AO22CHD U5547 (.O(n4122), 
	.B2(n503), 
	.B1(\ram[221][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n363));
   AO22CHD U5548 (.O(n4123), 
	.B2(n503), 
	.B1(\ram[221][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n363));
   AO22CHD U5549 (.O(n4124), 
	.B2(n503), 
	.B1(\ram[221][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n363));
   AO22CHD U5550 (.O(n4125), 
	.B2(n503), 
	.B1(\ram[221][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n363));
   AO22CHD U5551 (.O(n4126), 
	.B2(n503), 
	.B1(\ram[221][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n363));
   AO22CHD U5552 (.O(n4127), 
	.B2(n503), 
	.B1(\ram[221][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n363));
   AO22CHD U5553 (.O(n4128), 
	.B2(n503), 
	.B1(\ram[221][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n363));
   AO22CHD U5554 (.O(n4129), 
	.B2(n503), 
	.B1(\ram[221][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n363));
   AO22CHD U5555 (.O(n4130), 
	.B2(n503), 
	.B1(\ram[221][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n363));
   AO22CHD U5556 (.O(n4131), 
	.B2(n503), 
	.B1(\ram[221][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n363));
   AO22CHD U5557 (.O(n4132), 
	.B2(n503), 
	.B1(\ram[221][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n363));
   AO22CHD U5558 (.O(n4133), 
	.B2(n503), 
	.B1(\ram[221][15] ), 
	.A2(n23), 
	.A1(n363));
   AO22CHD U5559 (.O(n4134), 
	.B2(n505), 
	.B1(\ram[222][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n365));
   AO22CHD U5560 (.O(n4135), 
	.B2(n505), 
	.B1(\ram[222][1] ), 
	.A2(n9), 
	.A1(n365));
   AO22CHD U5561 (.O(n4136), 
	.B2(n505), 
	.B1(\ram[222][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n365));
   AO22CHD U5562 (.O(n4137), 
	.B2(n505), 
	.B1(\ram[222][3] ), 
	.A2(n11), 
	.A1(n365));
   AO22CHD U5563 (.O(n4138), 
	.B2(n505), 
	.B1(\ram[222][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n365));
   AO22CHD U5564 (.O(n4139), 
	.B2(n505), 
	.B1(\ram[222][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n365));
   AO22CHD U5565 (.O(n4140), 
	.B2(n505), 
	.B1(\ram[222][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n365));
   AO22CHD U5566 (.O(n4141), 
	.B2(n505), 
	.B1(\ram[222][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n365));
   AO22CHD U5567 (.O(n4142), 
	.B2(n505), 
	.B1(\ram[222][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n365));
   AO22CHD U5568 (.O(n4143), 
	.B2(n505), 
	.B1(\ram[222][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n365));
   AO22CHD U5569 (.O(n4144), 
	.B2(n505), 
	.B1(\ram[222][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n365));
   AO22CHD U5570 (.O(n4145), 
	.B2(n505), 
	.B1(\ram[222][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n365));
   AO22CHD U5571 (.O(n4146), 
	.B2(n505), 
	.B1(\ram[222][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n365));
   AO22CHD U5572 (.O(n4147), 
	.B2(n505), 
	.B1(\ram[222][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n365));
   AO22CHD U5573 (.O(n4148), 
	.B2(n505), 
	.B1(\ram[222][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n365));
   AO22CHD U5574 (.O(n4149), 
	.B2(n505), 
	.B1(\ram[222][15] ), 
	.A2(n23), 
	.A1(n365));
   AO22CHD U5575 (.O(n4150), 
	.B2(n507), 
	.B1(\ram[223][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n367));
   AO22CHD U5576 (.O(n4151), 
	.B2(n507), 
	.B1(\ram[223][1] ), 
	.A2(n9), 
	.A1(n367));
   AO22CHD U5577 (.O(n4152), 
	.B2(n507), 
	.B1(\ram[223][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n367));
   AO22CHD U5578 (.O(n4153), 
	.B2(n507), 
	.B1(\ram[223][3] ), 
	.A2(n11), 
	.A1(n367));
   AO22CHD U5579 (.O(n4154), 
	.B2(n507), 
	.B1(\ram[223][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n367));
   AO22CHD U5580 (.O(n4155), 
	.B2(n507), 
	.B1(\ram[223][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n367));
   AO22CHD U5581 (.O(n4156), 
	.B2(n507), 
	.B1(\ram[223][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n367));
   AO22CHD U5582 (.O(n4157), 
	.B2(n507), 
	.B1(\ram[223][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n367));
   AO22CHD U5583 (.O(n4158), 
	.B2(n507), 
	.B1(\ram[223][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n367));
   AO22CHD U5584 (.O(n4159), 
	.B2(n507), 
	.B1(\ram[223][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n367));
   AO22CHD U5585 (.O(n4160), 
	.B2(n507), 
	.B1(\ram[223][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n367));
   AO22CHD U5586 (.O(n4161), 
	.B2(n507), 
	.B1(\ram[223][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n367));
   AO22CHD U5587 (.O(n4162), 
	.B2(n507), 
	.B1(\ram[223][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n367));
   AO22CHD U5588 (.O(n4163), 
	.B2(n507), 
	.B1(\ram[223][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n367));
   AO22CHD U5589 (.O(n4164), 
	.B2(n507), 
	.B1(\ram[223][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n367));
   AO22CHD U5590 (.O(n4165), 
	.B2(n507), 
	.B1(\ram[223][15] ), 
	.A2(n23), 
	.A1(n367));
   AO22CHD U5591 (.O(n4166), 
	.B2(n509), 
	.B1(\ram[224][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n369));
   AO22CHD U5592 (.O(n4167), 
	.B2(n509), 
	.B1(\ram[224][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n369));
   AO22CHD U5593 (.O(n4168), 
	.B2(n509), 
	.B1(\ram[224][2] ), 
	.A2(n10), 
	.A1(n369));
   AO22CHD U5594 (.O(n4169), 
	.B2(n509), 
	.B1(\ram[224][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n369));
   AO22CHD U5595 (.O(n4170), 
	.B2(n509), 
	.B1(\ram[224][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n369));
   AO22CHD U5596 (.O(n4171), 
	.B2(n509), 
	.B1(\ram[224][5] ), 
	.A2(n13), 
	.A1(n369));
   AO22CHD U5597 (.O(n4172), 
	.B2(n509), 
	.B1(\ram[224][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n369));
   AO22CHD U5598 (.O(n4173), 
	.B2(n509), 
	.B1(\ram[224][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n369));
   AO22CHD U5599 (.O(n4174), 
	.B2(n509), 
	.B1(\ram[224][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n369));
   AO22CHD U5600 (.O(n4175), 
	.B2(n509), 
	.B1(\ram[224][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n369));
   AO22CHD U5601 (.O(n4176), 
	.B2(n509), 
	.B1(\ram[224][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n369));
   AO22CHD U5602 (.O(n4177), 
	.B2(n509), 
	.B1(\ram[224][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n369));
   AO22CHD U5603 (.O(n4178), 
	.B2(n509), 
	.B1(\ram[224][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n369));
   AO22CHD U5604 (.O(n4179), 
	.B2(n509), 
	.B1(\ram[224][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n369));
   AO22CHD U5605 (.O(n4180), 
	.B2(n509), 
	.B1(\ram[224][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n369));
   AO22CHD U5606 (.O(n4181), 
	.B2(n509), 
	.B1(\ram[224][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n369));
   AO22CHD U5607 (.O(n4182), 
	.B2(n512), 
	.B1(\ram[225][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n371));
   AO22CHD U5608 (.O(n4183), 
	.B2(n512), 
	.B1(\ram[225][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n371));
   AO22CHD U5609 (.O(n4184), 
	.B2(n512), 
	.B1(\ram[225][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n371));
   AO22CHD U5610 (.O(n4185), 
	.B2(n512), 
	.B1(\ram[225][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n371));
   AO22CHD U5611 (.O(n4186), 
	.B2(n512), 
	.B1(\ram[225][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n371));
   AO22CHD U5612 (.O(n4187), 
	.B2(n512), 
	.B1(\ram[225][5] ), 
	.A2(n13), 
	.A1(n371));
   AO22CHD U5613 (.O(n4188), 
	.B2(n512), 
	.B1(\ram[225][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n371));
   AO22CHD U5614 (.O(n4189), 
	.B2(n512), 
	.B1(\ram[225][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n371));
   AO22CHD U5615 (.O(n4190), 
	.B2(n512), 
	.B1(\ram[225][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n371));
   AO22CHD U5616 (.O(n4191), 
	.B2(n512), 
	.B1(\ram[225][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n371));
   AO22CHD U5617 (.O(n4192), 
	.B2(n512), 
	.B1(\ram[225][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n371));
   AO22CHD U5618 (.O(n4193), 
	.B2(n512), 
	.B1(\ram[225][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n371));
   AO22CHD U5619 (.O(n4194), 
	.B2(n512), 
	.B1(\ram[225][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n371));
   AO22CHD U5620 (.O(n4195), 
	.B2(n512), 
	.B1(\ram[225][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n371));
   AO22CHD U5621 (.O(n4196), 
	.B2(n512), 
	.B1(\ram[225][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n371));
   AO22CHD U5622 (.O(n4197), 
	.B2(n512), 
	.B1(\ram[225][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n371));
   AO22CHD U5623 (.O(n4198), 
	.B2(n514), 
	.B1(\ram[226][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n373));
   AO22CHD U5624 (.O(n4199), 
	.B2(n514), 
	.B1(\ram[226][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n373));
   AO22CHD U5625 (.O(n4200), 
	.B2(n514), 
	.B1(\ram[226][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n373));
   AO22CHD U5626 (.O(n4201), 
	.B2(n514), 
	.B1(\ram[226][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n373));
   AO22CHD U5627 (.O(n4202), 
	.B2(n514), 
	.B1(\ram[226][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n373));
   AO22CHD U5628 (.O(n4203), 
	.B2(n514), 
	.B1(\ram[226][5] ), 
	.A2(n13), 
	.A1(n373));
   AO22CHD U5629 (.O(n4204), 
	.B2(n514), 
	.B1(\ram[226][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n373));
   AO22CHD U5630 (.O(n4205), 
	.B2(n514), 
	.B1(\ram[226][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n373));
   AO22CHD U5631 (.O(n4206), 
	.B2(n514), 
	.B1(\ram[226][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n373));
   AO22CHD U5632 (.O(n4207), 
	.B2(n514), 
	.B1(\ram[226][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n373));
   AO22CHD U5633 (.O(n4208), 
	.B2(n514), 
	.B1(\ram[226][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n373));
   AO22CHD U5634 (.O(n4209), 
	.B2(n514), 
	.B1(\ram[226][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n373));
   AO22CHD U5635 (.O(n4210), 
	.B2(n514), 
	.B1(\ram[226][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n373));
   AO22CHD U5636 (.O(n4211), 
	.B2(n514), 
	.B1(\ram[226][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n373));
   AO22CHD U5637 (.O(n4212), 
	.B2(n514), 
	.B1(\ram[226][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n373));
   AO22CHD U5638 (.O(n4213), 
	.B2(n514), 
	.B1(\ram[226][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n373));
   AO22CHD U5639 (.O(n4214), 
	.B2(n516), 
	.B1(\ram[227][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n375));
   AO22CHD U5640 (.O(n4215), 
	.B2(n516), 
	.B1(\ram[227][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n375));
   AO22CHD U5641 (.O(n4216), 
	.B2(n516), 
	.B1(\ram[227][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n375));
   AO22CHD U5642 (.O(n4217), 
	.B2(n516), 
	.B1(\ram[227][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n375));
   AO22CHD U5643 (.O(n4218), 
	.B2(n516), 
	.B1(\ram[227][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n375));
   AO22CHD U5644 (.O(n4219), 
	.B2(n516), 
	.B1(\ram[227][5] ), 
	.A2(n13), 
	.A1(n375));
   AO22CHD U5645 (.O(n4220), 
	.B2(n516), 
	.B1(\ram[227][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n375));
   AO22CHD U5646 (.O(n4221), 
	.B2(n516), 
	.B1(\ram[227][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n375));
   AO22CHD U5647 (.O(n4222), 
	.B2(n516), 
	.B1(\ram[227][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n375));
   AO22CHD U5648 (.O(n4223), 
	.B2(n516), 
	.B1(\ram[227][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n375));
   AO22CHD U5649 (.O(n4224), 
	.B2(n516), 
	.B1(\ram[227][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n375));
   AO22CHD U5650 (.O(n4225), 
	.B2(n516), 
	.B1(\ram[227][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n375));
   AO22CHD U5651 (.O(n4226), 
	.B2(n516), 
	.B1(\ram[227][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n375));
   AO22CHD U5652 (.O(n4227), 
	.B2(n516), 
	.B1(\ram[227][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n375));
   AO22CHD U5653 (.O(n4228), 
	.B2(n516), 
	.B1(\ram[227][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n375));
   AO22CHD U5654 (.O(n4229), 
	.B2(n516), 
	.B1(\ram[227][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n375));
   AO22CHD U5655 (.O(n4230), 
	.B2(n518), 
	.B1(\ram[228][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n377));
   AO22CHD U5656 (.O(n4231), 
	.B2(n518), 
	.B1(\ram[228][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n377));
   AO22CHD U5657 (.O(n4232), 
	.B2(n518), 
	.B1(\ram[228][2] ), 
	.A2(n10), 
	.A1(n377));
   AO22CHD U5658 (.O(n4233), 
	.B2(n518), 
	.B1(\ram[228][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n377));
   AO22CHD U5659 (.O(n4234), 
	.B2(n518), 
	.B1(\ram[228][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n377));
   AO22CHD U5660 (.O(n4235), 
	.B2(n518), 
	.B1(\ram[228][5] ), 
	.A2(n13), 
	.A1(n377));
   AO22CHD U5661 (.O(n4236), 
	.B2(n518), 
	.B1(\ram[228][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n377));
   AO22CHD U5662 (.O(n4237), 
	.B2(n518), 
	.B1(\ram[228][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n377));
   AO22CHD U5663 (.O(n4238), 
	.B2(n518), 
	.B1(\ram[228][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n377));
   AO22CHD U5664 (.O(n4239), 
	.B2(n518), 
	.B1(\ram[228][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n377));
   AO22CHD U5665 (.O(n4240), 
	.B2(n518), 
	.B1(\ram[228][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n377));
   AO22CHD U5666 (.O(n4241), 
	.B2(n518), 
	.B1(\ram[228][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n377));
   AO22CHD U5667 (.O(n4242), 
	.B2(n518), 
	.B1(\ram[228][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n377));
   AO22CHD U5668 (.O(n4243), 
	.B2(n518), 
	.B1(\ram[228][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n377));
   AO22CHD U5669 (.O(n4244), 
	.B2(n518), 
	.B1(\ram[228][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n377));
   AO22CHD U5670 (.O(n4245), 
	.B2(n518), 
	.B1(\ram[228][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n377));
   AO22CHD U5671 (.O(n4246), 
	.B2(n520), 
	.B1(\ram[229][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n378));
   AO22CHD U5672 (.O(n4247), 
	.B2(n520), 
	.B1(\ram[229][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n378));
   AO22CHD U5673 (.O(n4248), 
	.B2(n520), 
	.B1(\ram[229][2] ), 
	.A2(n10), 
	.A1(n378));
   AO22CHD U5674 (.O(n4249), 
	.B2(n520), 
	.B1(\ram[229][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n378));
   AO22CHD U5675 (.O(n4250), 
	.B2(n520), 
	.B1(\ram[229][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n378));
   AO22CHD U5676 (.O(n4251), 
	.B2(n520), 
	.B1(\ram[229][5] ), 
	.A2(n13), 
	.A1(n378));
   AO22CHD U5677 (.O(n4252), 
	.B2(n520), 
	.B1(\ram[229][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n378));
   AO22CHD U5678 (.O(n4253), 
	.B2(n520), 
	.B1(\ram[229][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n378));
   AO22CHD U5679 (.O(n4254), 
	.B2(n520), 
	.B1(\ram[229][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n378));
   AO22CHD U5680 (.O(n4255), 
	.B2(n520), 
	.B1(\ram[229][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n378));
   AO22CHD U5681 (.O(n4256), 
	.B2(n520), 
	.B1(\ram[229][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n378));
   AO22CHD U5682 (.O(n4257), 
	.B2(n520), 
	.B1(\ram[229][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n378));
   AO22CHD U5683 (.O(n4258), 
	.B2(n520), 
	.B1(\ram[229][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n378));
   AO22CHD U5684 (.O(n4259), 
	.B2(n520), 
	.B1(\ram[229][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n378));
   AO22CHD U5685 (.O(n4260), 
	.B2(n520), 
	.B1(\ram[229][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n378));
   AO22CHD U5686 (.O(n4261), 
	.B2(n520), 
	.B1(\ram[229][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n378));
   AO22CHD U5687 (.O(n4262), 
	.B2(n522), 
	.B1(\ram[230][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n380));
   AO22CHD U5688 (.O(n4263), 
	.B2(n522), 
	.B1(\ram[230][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n380));
   AO22CHD U5689 (.O(n4264), 
	.B2(n522), 
	.B1(\ram[230][2] ), 
	.A2(n10), 
	.A1(n380));
   AO22CHD U5690 (.O(n4265), 
	.B2(n522), 
	.B1(\ram[230][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n380));
   AO22CHD U5691 (.O(n4266), 
	.B2(n522), 
	.B1(\ram[230][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n380));
   AO22CHD U5692 (.O(n4267), 
	.B2(n522), 
	.B1(\ram[230][5] ), 
	.A2(n13), 
	.A1(n380));
   AO22CHD U5693 (.O(n4268), 
	.B2(n522), 
	.B1(\ram[230][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n380));
   AO22CHD U5694 (.O(n4269), 
	.B2(n522), 
	.B1(\ram[230][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n380));
   AO22CHD U5695 (.O(n4270), 
	.B2(n522), 
	.B1(\ram[230][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n380));
   AO22CHD U5696 (.O(n4271), 
	.B2(n522), 
	.B1(\ram[230][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n380));
   AO22CHD U5697 (.O(n4272), 
	.B2(n522), 
	.B1(\ram[230][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n380));
   AO22CHD U5698 (.O(n4273), 
	.B2(n522), 
	.B1(\ram[230][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n380));
   AO22CHD U5699 (.O(n4274), 
	.B2(n522), 
	.B1(\ram[230][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n380));
   AO22CHD U5700 (.O(n4275), 
	.B2(n522), 
	.B1(\ram[230][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n380));
   AO22CHD U5701 (.O(n4276), 
	.B2(n522), 
	.B1(\ram[230][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n380));
   AO22CHD U5702 (.O(n4277), 
	.B2(n522), 
	.B1(\ram[230][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n380));
   AO22CHD U5703 (.O(n4278), 
	.B2(n524), 
	.B1(\ram[231][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n382));
   AO22CHD U5704 (.O(n4279), 
	.B2(n524), 
	.B1(\ram[231][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n382));
   AO22CHD U5705 (.O(n4280), 
	.B2(n524), 
	.B1(\ram[231][2] ), 
	.A2(n10), 
	.A1(n382));
   AO22CHD U5706 (.O(n4281), 
	.B2(n524), 
	.B1(\ram[231][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n382));
   AO22CHD U5707 (.O(n4282), 
	.B2(n524), 
	.B1(\ram[231][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n382));
   AO22CHD U5708 (.O(n4283), 
	.B2(n524), 
	.B1(\ram[231][5] ), 
	.A2(n13), 
	.A1(n382));
   AO22CHD U5709 (.O(n4284), 
	.B2(n524), 
	.B1(\ram[231][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n382));
   AO22CHD U5710 (.O(n4285), 
	.B2(n524), 
	.B1(\ram[231][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n382));
   AO22CHD U5711 (.O(n4286), 
	.B2(n524), 
	.B1(\ram[231][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n382));
   AO22CHD U5712 (.O(n4287), 
	.B2(n524), 
	.B1(\ram[231][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n382));
   AO22CHD U5713 (.O(n4288), 
	.B2(n524), 
	.B1(\ram[231][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n382));
   AO22CHD U5714 (.O(n4289), 
	.B2(n524), 
	.B1(\ram[231][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n382));
   AO22CHD U5715 (.O(n4290), 
	.B2(n524), 
	.B1(\ram[231][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n382));
   AO22CHD U5716 (.O(n4291), 
	.B2(n524), 
	.B1(\ram[231][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n382));
   AO22CHD U5717 (.O(n4292), 
	.B2(n524), 
	.B1(\ram[231][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n382));
   AO22CHD U5718 (.O(n4293), 
	.B2(n524), 
	.B1(\ram[231][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n382));
   AO22CHD U5719 (.O(n4294), 
	.B2(n526), 
	.B1(\ram[232][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n384));
   AO22CHD U5720 (.O(n4295), 
	.B2(n526), 
	.B1(\ram[232][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n384));
   AO22CHD U5721 (.O(n4296), 
	.B2(n526), 
	.B1(\ram[232][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n384));
   AO22CHD U5722 (.O(n4297), 
	.B2(n526), 
	.B1(\ram[232][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n384));
   AO22CHD U5723 (.O(n4298), 
	.B2(n526), 
	.B1(\ram[232][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n384));
   AO22CHD U5724 (.O(n4299), 
	.B2(n526), 
	.B1(\ram[232][5] ), 
	.A2(n13), 
	.A1(n384));
   AO22CHD U5725 (.O(n4300), 
	.B2(n526), 
	.B1(\ram[232][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n384));
   AO22CHD U5726 (.O(n4301), 
	.B2(n526), 
	.B1(\ram[232][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n384));
   AO22CHD U5727 (.O(n4302), 
	.B2(n526), 
	.B1(\ram[232][8] ), 
	.A2(n16), 
	.A1(n384));
   AO22CHD U5728 (.O(n4303), 
	.B2(n526), 
	.B1(\ram[232][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n384));
   AO22CHD U5729 (.O(n4304), 
	.B2(n526), 
	.B1(\ram[232][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n384));
   AO22CHD U5730 (.O(n4305), 
	.B2(n526), 
	.B1(\ram[232][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n384));
   AO22CHD U5731 (.O(n4306), 
	.B2(n526), 
	.B1(\ram[232][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n384));
   AO22CHD U5732 (.O(n4307), 
	.B2(n526), 
	.B1(\ram[232][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n384));
   AO22CHD U5733 (.O(n4308), 
	.B2(n526), 
	.B1(\ram[232][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n384));
   AO22CHD U5734 (.O(n4309), 
	.B2(n526), 
	.B1(\ram[232][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n384));
   AO22CHD U5735 (.O(n4310), 
	.B2(n528), 
	.B1(\ram[233][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n386));
   AO22CHD U5736 (.O(n4311), 
	.B2(n528), 
	.B1(\ram[233][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n386));
   AO22CHD U5737 (.O(n4312), 
	.B2(n528), 
	.B1(\ram[233][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n386));
   AO22CHD U5738 (.O(n4313), 
	.B2(n528), 
	.B1(\ram[233][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n386));
   AO22CHD U5739 (.O(n4314), 
	.B2(n528), 
	.B1(\ram[233][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n386));
   AO22CHD U5740 (.O(n4315), 
	.B2(n528), 
	.B1(\ram[233][5] ), 
	.A2(n13), 
	.A1(n386));
   AO22CHD U5741 (.O(n4316), 
	.B2(n528), 
	.B1(\ram[233][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n386));
   AO22CHD U5742 (.O(n4317), 
	.B2(n528), 
	.B1(\ram[233][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n386));
   AO22CHD U5743 (.O(n4318), 
	.B2(n528), 
	.B1(\ram[233][8] ), 
	.A2(n16), 
	.A1(n386));
   AO22CHD U5744 (.O(n4319), 
	.B2(n528), 
	.B1(\ram[233][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n386));
   AO22CHD U5745 (.O(n4320), 
	.B2(n528), 
	.B1(\ram[233][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n386));
   AO22CHD U5746 (.O(n4321), 
	.B2(n528), 
	.B1(\ram[233][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n386));
   AO22CHD U5747 (.O(n4322), 
	.B2(n528), 
	.B1(\ram[233][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n386));
   AO22CHD U5748 (.O(n4323), 
	.B2(n528), 
	.B1(\ram[233][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n386));
   AO22CHD U5749 (.O(n4324), 
	.B2(n528), 
	.B1(\ram[233][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n386));
   AO22CHD U5750 (.O(n4325), 
	.B2(n528), 
	.B1(\ram[233][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n386));
   AO22CHD U5751 (.O(n4326), 
	.B2(n530), 
	.B1(\ram[234][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n388));
   AO22CHD U5752 (.O(n4327), 
	.B2(n530), 
	.B1(\ram[234][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n388));
   AO22CHD U5753 (.O(n4328), 
	.B2(n530), 
	.B1(\ram[234][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n388));
   AO22CHD U5754 (.O(n4329), 
	.B2(n530), 
	.B1(\ram[234][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n388));
   AO22CHD U5755 (.O(n4330), 
	.B2(n530), 
	.B1(\ram[234][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n388));
   AO22CHD U5756 (.O(n4331), 
	.B2(n530), 
	.B1(\ram[234][5] ), 
	.A2(n13), 
	.A1(n388));
   AO22CHD U5757 (.O(n4332), 
	.B2(n530), 
	.B1(\ram[234][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n388));
   AO22CHD U5758 (.O(n4333), 
	.B2(n530), 
	.B1(\ram[234][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n388));
   AO22CHD U5759 (.O(n4334), 
	.B2(n530), 
	.B1(\ram[234][8] ), 
	.A2(n16), 
	.A1(n388));
   AO22CHD U5760 (.O(n4335), 
	.B2(n530), 
	.B1(\ram[234][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n388));
   AO22CHD U5761 (.O(n4336), 
	.B2(n530), 
	.B1(\ram[234][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n388));
   AO22CHD U5762 (.O(n4337), 
	.B2(n530), 
	.B1(\ram[234][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n388));
   AO22CHD U5763 (.O(n4338), 
	.B2(n530), 
	.B1(\ram[234][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n388));
   AO22CHD U5764 (.O(n4339), 
	.B2(n530), 
	.B1(\ram[234][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n388));
   AO22CHD U5765 (.O(n4340), 
	.B2(n530), 
	.B1(\ram[234][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n388));
   AO22CHD U5766 (.O(n4341), 
	.B2(n530), 
	.B1(\ram[234][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n388));
   AO22CHD U5767 (.O(n4342), 
	.B2(n532), 
	.B1(\ram[235][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n390));
   AO22CHD U5768 (.O(n4343), 
	.B2(n532), 
	.B1(\ram[235][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n390));
   AO22CHD U5769 (.O(n4344), 
	.B2(n532), 
	.B1(\ram[235][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n390));
   AO22CHD U5770 (.O(n4345), 
	.B2(n532), 
	.B1(\ram[235][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n390));
   AO22CHD U5771 (.O(n4346), 
	.B2(n532), 
	.B1(\ram[235][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n390));
   AO22CHD U5772 (.O(n4347), 
	.B2(n532), 
	.B1(\ram[235][5] ), 
	.A2(n13), 
	.A1(n390));
   AO22CHD U5773 (.O(n4348), 
	.B2(n532), 
	.B1(\ram[235][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n390));
   AO22CHD U5774 (.O(n4349), 
	.B2(n532), 
	.B1(\ram[235][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n390));
   AO22CHD U5775 (.O(n4350), 
	.B2(n532), 
	.B1(\ram[235][8] ), 
	.A2(n16), 
	.A1(n390));
   AO22CHD U5776 (.O(n4351), 
	.B2(n532), 
	.B1(\ram[235][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n390));
   AO22CHD U5777 (.O(n4352), 
	.B2(n532), 
	.B1(\ram[235][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n390));
   AO22CHD U5778 (.O(n4353), 
	.B2(n532), 
	.B1(\ram[235][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n390));
   AO22CHD U5779 (.O(n4354), 
	.B2(n532), 
	.B1(\ram[235][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n390));
   AO22CHD U5780 (.O(n4355), 
	.B2(n532), 
	.B1(\ram[235][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n390));
   AO22CHD U5781 (.O(n4356), 
	.B2(n532), 
	.B1(\ram[235][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n390));
   AO22CHD U5782 (.O(n4357), 
	.B2(n532), 
	.B1(\ram[235][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n390));
   AO22CHD U5783 (.O(n4358), 
	.B2(n534), 
	.B1(\ram[236][0] ), 
	.A2(n6), 
	.A1(n392));
   AO22CHD U5784 (.O(n4359), 
	.B2(n534), 
	.B1(\ram[236][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n392));
   AO22CHD U5785 (.O(n4360), 
	.B2(n534), 
	.B1(\ram[236][2] ), 
	.A2(n10), 
	.A1(n392));
   AO22CHD U5786 (.O(n4361), 
	.B2(n534), 
	.B1(\ram[236][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n392));
   AO22CHD U5787 (.O(n4362), 
	.B2(n534), 
	.B1(\ram[236][4] ), 
	.A2(n12), 
	.A1(n392));
   AO22CHD U5788 (.O(n4363), 
	.B2(n534), 
	.B1(\ram[236][5] ), 
	.A2(n13), 
	.A1(n392));
   AO22CHD U5789 (.O(n4364), 
	.B2(n534), 
	.B1(\ram[236][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n392));
   AO22CHD U5790 (.O(n4365), 
	.B2(n534), 
	.B1(\ram[236][7] ), 
	.A2(n15), 
	.A1(n392));
   AO22CHD U5791 (.O(n4366), 
	.B2(n534), 
	.B1(\ram[236][8] ), 
	.A2(n16), 
	.A1(n392));
   AO22CHD U5792 (.O(n4367), 
	.B2(n534), 
	.B1(\ram[236][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n392));
   AO22CHD U5793 (.O(n4368), 
	.B2(n534), 
	.B1(\ram[236][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n392));
   AO22CHD U5794 (.O(n4369), 
	.B2(n534), 
	.B1(\ram[236][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n392));
   AO22CHD U5795 (.O(n4370), 
	.B2(n534), 
	.B1(\ram[236][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n392));
   AO22CHD U5796 (.O(n4371), 
	.B2(n534), 
	.B1(\ram[236][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n392));
   AO22CHD U5797 (.O(n4372), 
	.B2(n534), 
	.B1(\ram[236][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n392));
   AO22CHD U5798 (.O(n4373), 
	.B2(n534), 
	.B1(\ram[236][15] ), 
	.A2(n23), 
	.A1(n392));
   AO22CHD U5799 (.O(n4374), 
	.B2(n536), 
	.B1(\ram[237][0] ), 
	.A2(n6), 
	.A1(n394));
   AO22CHD U5800 (.O(n4375), 
	.B2(n536), 
	.B1(\ram[237][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n394));
   AO22CHD U5801 (.O(n4376), 
	.B2(n536), 
	.B1(\ram[237][2] ), 
	.A2(n10), 
	.A1(n394));
   AO22CHD U5802 (.O(n4377), 
	.B2(n536), 
	.B1(\ram[237][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n394));
   AO22CHD U5803 (.O(n4378), 
	.B2(n536), 
	.B1(\ram[237][4] ), 
	.A2(n12), 
	.A1(n394));
   AO22CHD U5804 (.O(n4379), 
	.B2(n536), 
	.B1(\ram[237][5] ), 
	.A2(n13), 
	.A1(n394));
   AO22CHD U5805 (.O(n4380), 
	.B2(n536), 
	.B1(\ram[237][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n394));
   AO22CHD U5806 (.O(n4381), 
	.B2(n536), 
	.B1(\ram[237][7] ), 
	.A2(n15), 
	.A1(n394));
   AO22CHD U5807 (.O(n4382), 
	.B2(n536), 
	.B1(\ram[237][8] ), 
	.A2(n16), 
	.A1(n394));
   AO22CHD U5808 (.O(n4383), 
	.B2(n536), 
	.B1(\ram[237][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n394));
   AO22CHD U5809 (.O(n4384), 
	.B2(n536), 
	.B1(\ram[237][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n394));
   AO22CHD U5810 (.O(n4385), 
	.B2(n536), 
	.B1(\ram[237][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n394));
   AO22CHD U5811 (.O(n4386), 
	.B2(n536), 
	.B1(\ram[237][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n394));
   AO22CHD U5812 (.O(n4387), 
	.B2(n536), 
	.B1(\ram[237][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n394));
   AO22CHD U5813 (.O(n4388), 
	.B2(n536), 
	.B1(\ram[237][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n394));
   AO22CHD U5814 (.O(n4389), 
	.B2(n536), 
	.B1(\ram[237][15] ), 
	.A2(n23), 
	.A1(n394));
   AO22CHD U5815 (.O(n4390), 
	.B2(n538), 
	.B1(\ram[238][0] ), 
	.A2(n6), 
	.A1(n396));
   AO22CHD U5816 (.O(n4391), 
	.B2(n538), 
	.B1(\ram[238][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n396));
   AO22CHD U5817 (.O(n4392), 
	.B2(n538), 
	.B1(\ram[238][2] ), 
	.A2(n10), 
	.A1(n396));
   AO22CHD U5818 (.O(n4393), 
	.B2(n538), 
	.B1(\ram[238][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n396));
   AO22CHD U5819 (.O(n4394), 
	.B2(n538), 
	.B1(\ram[238][4] ), 
	.A2(n12), 
	.A1(n396));
   AO22CHD U5820 (.O(n4395), 
	.B2(n538), 
	.B1(\ram[238][5] ), 
	.A2(n13), 
	.A1(n396));
   AO22CHD U5821 (.O(n4396), 
	.B2(n538), 
	.B1(\ram[238][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n396));
   AO22CHD U5822 (.O(n4397), 
	.B2(n538), 
	.B1(\ram[238][7] ), 
	.A2(n15), 
	.A1(n396));
   AO22CHD U5823 (.O(n4398), 
	.B2(n538), 
	.B1(\ram[238][8] ), 
	.A2(n16), 
	.A1(n396));
   AO22CHD U5824 (.O(n4399), 
	.B2(n538), 
	.B1(\ram[238][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n396));
   AO22CHD U5825 (.O(n4400), 
	.B2(n538), 
	.B1(\ram[238][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n396));
   AO22CHD U5826 (.O(n4401), 
	.B2(n538), 
	.B1(\ram[238][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n396));
   AO22CHD U5827 (.O(n4402), 
	.B2(n538), 
	.B1(\ram[238][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n396));
   AO22CHD U5828 (.O(n4403), 
	.B2(n538), 
	.B1(\ram[238][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n396));
   AO22CHD U5829 (.O(n4404), 
	.B2(n538), 
	.B1(\ram[238][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n396));
   AO22CHD U5830 (.O(n4405), 
	.B2(n538), 
	.B1(\ram[238][15] ), 
	.A2(n23), 
	.A1(n396));
   AO22CHD U5831 (.O(n4406), 
	.B2(n540), 
	.B1(\ram[239][0] ), 
	.A2(n6), 
	.A1(n398));
   AO22CHD U5832 (.O(n4407), 
	.B2(n540), 
	.B1(\ram[239][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n398));
   AO22CHD U5833 (.O(n4408), 
	.B2(n540), 
	.B1(\ram[239][2] ), 
	.A2(n10), 
	.A1(n398));
   AO22CHD U5834 (.O(n4409), 
	.B2(n540), 
	.B1(\ram[239][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n398));
   AO22CHD U5835 (.O(n4410), 
	.B2(n540), 
	.B1(\ram[239][4] ), 
	.A2(n12), 
	.A1(n398));
   AO22CHD U5836 (.O(n4411), 
	.B2(n540), 
	.B1(\ram[239][5] ), 
	.A2(n13), 
	.A1(n398));
   AO22CHD U5837 (.O(n4412), 
	.B2(n540), 
	.B1(\ram[239][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n398));
   AO22CHD U5838 (.O(n4413), 
	.B2(n540), 
	.B1(\ram[239][7] ), 
	.A2(n15), 
	.A1(n398));
   AO22CHD U5839 (.O(n4414), 
	.B2(n540), 
	.B1(\ram[239][8] ), 
	.A2(n16), 
	.A1(n398));
   AO22CHD U5840 (.O(n4415), 
	.B2(n540), 
	.B1(\ram[239][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n398));
   AO22CHD U5841 (.O(n4416), 
	.B2(n540), 
	.B1(\ram[239][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n398));
   AO22CHD U5842 (.O(n4417), 
	.B2(n540), 
	.B1(\ram[239][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n398));
   AO22CHD U5843 (.O(n4418), 
	.B2(n540), 
	.B1(\ram[239][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n398));
   AO22CHD U5844 (.O(n4419), 
	.B2(n540), 
	.B1(\ram[239][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n398));
   AO22CHD U5845 (.O(n4420), 
	.B2(n540), 
	.B1(\ram[239][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n398));
   AO22CHD U5846 (.O(n4421), 
	.B2(n540), 
	.B1(\ram[239][15] ), 
	.A2(n23), 
	.A1(n398));
   AO22CHD U5847 (.O(n4422), 
	.B2(n542), 
	.B1(\ram[240][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n400));
   AO22CHD U5848 (.O(n4423), 
	.B2(n542), 
	.B1(\ram[240][1] ), 
	.A2(n9), 
	.A1(n400));
   AO22CHD U5849 (.O(n4424), 
	.B2(n542), 
	.B1(\ram[240][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n400));
   AO22CHD U5850 (.O(n4425), 
	.B2(n542), 
	.B1(\ram[240][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n400));
   AO22CHD U5851 (.O(n4426), 
	.B2(n542), 
	.B1(\ram[240][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n400));
   AO22CHD U5852 (.O(n4427), 
	.B2(n542), 
	.B1(\ram[240][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n400));
   AO22CHD U5853 (.O(n4428), 
	.B2(n542), 
	.B1(\ram[240][6] ), 
	.A2(n14), 
	.A1(n400));
   AO22CHD U5854 (.O(n4429), 
	.B2(n542), 
	.B1(\ram[240][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n400));
   AO22CHD U5855 (.O(n4430), 
	.B2(n542), 
	.B1(\ram[240][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n400));
   AO22CHD U5856 (.O(n4431), 
	.B2(n542), 
	.B1(\ram[240][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n400));
   AO22CHD U5857 (.O(n4432), 
	.B2(n542), 
	.B1(\ram[240][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n400));
   AO22CHD U5858 (.O(n4433), 
	.B2(n542), 
	.B1(\ram[240][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n400));
   AO22CHD U5859 (.O(n4434), 
	.B2(n542), 
	.B1(\ram[240][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n400));
   AO22CHD U5860 (.O(n4435), 
	.B2(n542), 
	.B1(\ram[240][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n400));
   AO22CHD U5861 (.O(n4436), 
	.B2(n542), 
	.B1(\ram[240][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n400));
   AO22CHD U5862 (.O(n4437), 
	.B2(n542), 
	.B1(\ram[240][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n400));
   AO22CHD U5863 (.O(n4438), 
	.B2(n547), 
	.B1(\ram[241][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n402));
   AO22CHD U5864 (.O(n4439), 
	.B2(n547), 
	.B1(\ram[241][1] ), 
	.A2(n9), 
	.A1(n402));
   AO22CHD U5865 (.O(n4440), 
	.B2(n547), 
	.B1(\ram[241][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n402));
   AO22CHD U5866 (.O(n4441), 
	.B2(n547), 
	.B1(\ram[241][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n402));
   AO22CHD U5867 (.O(n4442), 
	.B2(n547), 
	.B1(\ram[241][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n402));
   AO22CHD U5868 (.O(n4443), 
	.B2(n547), 
	.B1(\ram[241][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n402));
   AO22CHD U5869 (.O(n4444), 
	.B2(n547), 
	.B1(\ram[241][6] ), 
	.A2(n14), 
	.A1(n402));
   AO22CHD U5870 (.O(n4445), 
	.B2(n547), 
	.B1(\ram[241][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n402));
   AO22CHD U5871 (.O(n4446), 
	.B2(n547), 
	.B1(\ram[241][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n402));
   AO22CHD U5872 (.O(n4447), 
	.B2(n547), 
	.B1(\ram[241][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n402));
   AO22CHD U5873 (.O(n4448), 
	.B2(n547), 
	.B1(\ram[241][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n402));
   AO22CHD U5874 (.O(n4449), 
	.B2(n547), 
	.B1(\ram[241][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n402));
   AO22CHD U5875 (.O(n4450), 
	.B2(n547), 
	.B1(\ram[241][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n402));
   AO22CHD U5876 (.O(n4451), 
	.B2(n547), 
	.B1(\ram[241][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n402));
   AO22CHD U5877 (.O(n4452), 
	.B2(n547), 
	.B1(\ram[241][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n402));
   AO22CHD U5878 (.O(n4453), 
	.B2(n547), 
	.B1(\ram[241][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n402));
   AO22CHD U5879 (.O(n4454), 
	.B2(n550), 
	.B1(\ram[242][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n404));
   AO22CHD U5880 (.O(n4455), 
	.B2(n550), 
	.B1(\ram[242][1] ), 
	.A2(n9), 
	.A1(n404));
   AO22CHD U5881 (.O(n4456), 
	.B2(n550), 
	.B1(\ram[242][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n404));
   AO22CHD U5882 (.O(n4457), 
	.B2(n550), 
	.B1(\ram[242][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n404));
   AO22CHD U5883 (.O(n4458), 
	.B2(n550), 
	.B1(\ram[242][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n404));
   AO22CHD U5884 (.O(n4459), 
	.B2(n550), 
	.B1(\ram[242][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n404));
   AO22CHD U5885 (.O(n4460), 
	.B2(n550), 
	.B1(\ram[242][6] ), 
	.A2(n14), 
	.A1(n404));
   AO22CHD U5886 (.O(n4461), 
	.B2(n550), 
	.B1(\ram[242][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n404));
   AO22CHD U5887 (.O(n4462), 
	.B2(n550), 
	.B1(\ram[242][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n404));
   AO22CHD U5888 (.O(n4463), 
	.B2(n550), 
	.B1(\ram[242][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n404));
   AO22CHD U5889 (.O(n4464), 
	.B2(n550), 
	.B1(\ram[242][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n404));
   AO22CHD U5890 (.O(n4465), 
	.B2(n550), 
	.B1(\ram[242][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n404));
   AO22CHD U5891 (.O(n4466), 
	.B2(n550), 
	.B1(\ram[242][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n404));
   AO22CHD U5892 (.O(n4467), 
	.B2(n550), 
	.B1(\ram[242][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n404));
   AO22CHD U5893 (.O(n4468), 
	.B2(n550), 
	.B1(\ram[242][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n404));
   AO22CHD U5894 (.O(n4469), 
	.B2(n550), 
	.B1(\ram[242][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n404));
   AO22CHD U5895 (.O(n4470), 
	.B2(n553), 
	.B1(\ram[243][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n406));
   AO22CHD U5896 (.O(n4471), 
	.B2(n553), 
	.B1(\ram[243][1] ), 
	.A2(n9), 
	.A1(n406));
   AO22CHD U5897 (.O(n4472), 
	.B2(n553), 
	.B1(\ram[243][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n406));
   AO22CHD U5898 (.O(n4473), 
	.B2(n553), 
	.B1(\ram[243][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n406));
   AO22CHD U5899 (.O(n4474), 
	.B2(n553), 
	.B1(\ram[243][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n406));
   AO22CHD U5900 (.O(n4475), 
	.B2(n553), 
	.B1(\ram[243][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n406));
   AO22CHD U5901 (.O(n4476), 
	.B2(n553), 
	.B1(\ram[243][6] ), 
	.A2(n14), 
	.A1(n406));
   AO22CHD U5902 (.O(n4477), 
	.B2(n553), 
	.B1(\ram[243][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n406));
   AO22CHD U5903 (.O(n4478), 
	.B2(n553), 
	.B1(\ram[243][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n406));
   AO22CHD U5904 (.O(n4479), 
	.B2(n553), 
	.B1(\ram[243][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n406));
   AO22CHD U5905 (.O(n4480), 
	.B2(n553), 
	.B1(\ram[243][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n406));
   AO22CHD U5906 (.O(n4481), 
	.B2(n553), 
	.B1(\ram[243][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n406));
   AO22CHD U5907 (.O(n4482), 
	.B2(n553), 
	.B1(\ram[243][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n406));
   AO22CHD U5908 (.O(n4483), 
	.B2(n553), 
	.B1(\ram[243][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n406));
   AO22CHD U5909 (.O(n4484), 
	.B2(n553), 
	.B1(\ram[243][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n406));
   AO22CHD U5910 (.O(n4485), 
	.B2(n553), 
	.B1(\ram[243][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n406));
   AO22CHD U5911 (.O(n4486), 
	.B2(n556), 
	.B1(\ram[244][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n408));
   AO22CHD U5912 (.O(n4487), 
	.B2(n556), 
	.B1(\ram[244][1] ), 
	.A2(n9), 
	.A1(n408));
   AO22CHD U5913 (.O(n4488), 
	.B2(n556), 
	.B1(\ram[244][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n408));
   AO22CHD U5914 (.O(n4489), 
	.B2(n556), 
	.B1(\ram[244][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n408));
   AO22CHD U5915 (.O(n4490), 
	.B2(n556), 
	.B1(\ram[244][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n408));
   AO22CHD U5916 (.O(n4491), 
	.B2(n556), 
	.B1(\ram[244][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n408));
   AO22CHD U5917 (.O(n4492), 
	.B2(n556), 
	.B1(\ram[244][6] ), 
	.A2(n14), 
	.A1(n408));
   AO22CHD U5918 (.O(n4493), 
	.B2(n556), 
	.B1(\ram[244][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n408));
   AO22CHD U5919 (.O(n4494), 
	.B2(n556), 
	.B1(\ram[244][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n408));
   AO22CHD U5920 (.O(n4495), 
	.B2(n556), 
	.B1(\ram[244][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n408));
   AO22CHD U5921 (.O(n4496), 
	.B2(n556), 
	.B1(\ram[244][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n408));
   AO22CHD U5922 (.O(n4497), 
	.B2(n556), 
	.B1(\ram[244][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n408));
   AO22CHD U5923 (.O(n4498), 
	.B2(n556), 
	.B1(\ram[244][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n408));
   AO22CHD U5924 (.O(n4499), 
	.B2(n556), 
	.B1(\ram[244][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n408));
   AO22CHD U5925 (.O(n4500), 
	.B2(n556), 
	.B1(\ram[244][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n408));
   AO22CHD U5926 (.O(n4501), 
	.B2(n556), 
	.B1(\ram[244][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n408));
   AO22CHD U5927 (.O(n4502), 
	.B2(n559), 
	.B1(\ram[245][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n410));
   AO22CHD U5928 (.O(n4503), 
	.B2(n559), 
	.B1(\ram[245][1] ), 
	.A2(n9), 
	.A1(n410));
   AO22CHD U5929 (.O(n4504), 
	.B2(n559), 
	.B1(\ram[245][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n410));
   AO22CHD U5930 (.O(n4505), 
	.B2(n559), 
	.B1(\ram[245][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n410));
   AO22CHD U5931 (.O(n4506), 
	.B2(n559), 
	.B1(\ram[245][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n410));
   AO22CHD U5932 (.O(n4507), 
	.B2(n559), 
	.B1(\ram[245][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n410));
   AO22CHD U5933 (.O(n4508), 
	.B2(n559), 
	.B1(\ram[245][6] ), 
	.A2(n14), 
	.A1(n410));
   AO22CHD U5934 (.O(n4509), 
	.B2(n559), 
	.B1(\ram[245][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n410));
   AO22CHD U5935 (.O(n4510), 
	.B2(n559), 
	.B1(\ram[245][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n410));
   AO22CHD U5936 (.O(n4511), 
	.B2(n559), 
	.B1(\ram[245][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n410));
   AO22CHD U5937 (.O(n4512), 
	.B2(n559), 
	.B1(\ram[245][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n410));
   AO22CHD U5938 (.O(n4513), 
	.B2(n559), 
	.B1(\ram[245][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n410));
   AO22CHD U5939 (.O(n4514), 
	.B2(n559), 
	.B1(\ram[245][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n410));
   AO22CHD U5940 (.O(n4515), 
	.B2(n559), 
	.B1(\ram[245][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n410));
   AO22CHD U5941 (.O(n4516), 
	.B2(n559), 
	.B1(\ram[245][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n410));
   AO22CHD U5942 (.O(n4517), 
	.B2(n559), 
	.B1(\ram[245][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n410));
   AO22CHD U5943 (.O(n4518), 
	.B2(n561), 
	.B1(\ram[246][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n411));
   AO22CHD U5944 (.O(n4519), 
	.B2(n561), 
	.B1(\ram[246][1] ), 
	.A2(n9), 
	.A1(n411));
   AO22CHD U5945 (.O(n4520), 
	.B2(n561), 
	.B1(\ram[246][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n411));
   AO22CHD U5946 (.O(n4521), 
	.B2(n561), 
	.B1(\ram[246][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n411));
   AO22CHD U5947 (.O(n4522), 
	.B2(n561), 
	.B1(\ram[246][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n411));
   AO22CHD U5948 (.O(n4523), 
	.B2(n561), 
	.B1(\ram[246][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n411));
   AO22CHD U5949 (.O(n4524), 
	.B2(n561), 
	.B1(\ram[246][6] ), 
	.A2(n14), 
	.A1(n411));
   AO22CHD U5950 (.O(n4525), 
	.B2(n561), 
	.B1(\ram[246][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n411));
   AO22CHD U5951 (.O(n4526), 
	.B2(n561), 
	.B1(\ram[246][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n411));
   AO22CHD U5952 (.O(n4527), 
	.B2(n561), 
	.B1(\ram[246][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n411));
   AO22CHD U5953 (.O(n4528), 
	.B2(n561), 
	.B1(\ram[246][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n411));
   AO22CHD U5954 (.O(n4529), 
	.B2(n561), 
	.B1(\ram[246][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n411));
   AO22CHD U5955 (.O(n4530), 
	.B2(n561), 
	.B1(\ram[246][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n411));
   AO22CHD U5956 (.O(n4531), 
	.B2(n561), 
	.B1(\ram[246][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n411));
   AO22CHD U5957 (.O(n4532), 
	.B2(n561), 
	.B1(\ram[246][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n411));
   AO22CHD U5958 (.O(n4533), 
	.B2(n561), 
	.B1(\ram[246][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n411));
   AO22CHD U5959 (.O(n4534), 
	.B2(n563), 
	.B1(\ram[247][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n413));
   AO22CHD U5960 (.O(n4535), 
	.B2(n563), 
	.B1(\ram[247][1] ), 
	.A2(n9), 
	.A1(n413));
   AO22CHD U5961 (.O(n4536), 
	.B2(n563), 
	.B1(\ram[247][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n413));
   AO22CHD U5962 (.O(n4537), 
	.B2(n563), 
	.B1(\ram[247][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n413));
   AO22CHD U5963 (.O(n4538), 
	.B2(n563), 
	.B1(\ram[247][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n413));
   AO22CHD U5964 (.O(n4539), 
	.B2(n563), 
	.B1(\ram[247][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n413));
   AO22CHD U5965 (.O(n4540), 
	.B2(n563), 
	.B1(\ram[247][6] ), 
	.A2(n14), 
	.A1(n413));
   AO22CHD U5966 (.O(n4541), 
	.B2(n563), 
	.B1(\ram[247][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n413));
   AO22CHD U5967 (.O(n4542), 
	.B2(n563), 
	.B1(\ram[247][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n413));
   AO22CHD U5968 (.O(n4543), 
	.B2(n563), 
	.B1(\ram[247][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n413));
   AO22CHD U5969 (.O(n4544), 
	.B2(n563), 
	.B1(\ram[247][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n413));
   AO22CHD U5970 (.O(n4545), 
	.B2(n563), 
	.B1(\ram[247][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n413));
   AO22CHD U5971 (.O(n4546), 
	.B2(n563), 
	.B1(\ram[247][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n413));
   AO22CHD U5972 (.O(n4547), 
	.B2(n563), 
	.B1(\ram[247][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n413));
   AO22CHD U5973 (.O(n4548), 
	.B2(n563), 
	.B1(\ram[247][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n413));
   AO22CHD U5974 (.O(n4549), 
	.B2(n563), 
	.B1(\ram[247][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n413));
   AO22CHD U5975 (.O(n4550), 
	.B2(n565), 
	.B1(\ram[248][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n415));
   AO22CHD U5976 (.O(n4551), 
	.B2(n565), 
	.B1(\ram[248][1] ), 
	.A2(n9), 
	.A1(n415));
   AO22CHD U5977 (.O(n4552), 
	.B2(n565), 
	.B1(\ram[248][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n415));
   AO22CHD U5978 (.O(n4553), 
	.B2(n565), 
	.B1(\ram[248][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n415));
   AO22CHD U5979 (.O(n4554), 
	.B2(n565), 
	.B1(\ram[248][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n415));
   AO22CHD U5980 (.O(n4555), 
	.B2(n565), 
	.B1(\ram[248][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n415));
   AO22CHD U5981 (.O(n4556), 
	.B2(n565), 
	.B1(\ram[248][6] ), 
	.A2(n14), 
	.A1(n415));
   AO22CHD U5982 (.O(n4557), 
	.B2(n565), 
	.B1(\ram[248][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n415));
   AO22CHD U5983 (.O(n4558), 
	.B2(n565), 
	.B1(\ram[248][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n415));
   AO22CHD U5984 (.O(n4559), 
	.B2(n565), 
	.B1(\ram[248][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n415));
   AO22CHD U5985 (.O(n4560), 
	.B2(n565), 
	.B1(\ram[248][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n415));
   AO22CHD U5986 (.O(n4561), 
	.B2(n565), 
	.B1(\ram[248][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n415));
   AO22CHD U5987 (.O(n4562), 
	.B2(n565), 
	.B1(\ram[248][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n415));
   AO22CHD U5988 (.O(n4563), 
	.B2(n565), 
	.B1(\ram[248][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n415));
   AO22CHD U5989 (.O(n4564), 
	.B2(n565), 
	.B1(\ram[248][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n415));
   AO22CHD U5990 (.O(n4565), 
	.B2(n565), 
	.B1(\ram[248][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n415));
   AO22CHD U5991 (.O(n4566), 
	.B2(n568), 
	.B1(\ram[249][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n417));
   AO22CHD U5992 (.O(n4567), 
	.B2(n568), 
	.B1(\ram[249][1] ), 
	.A2(n9), 
	.A1(n417));
   AO22CHD U5993 (.O(n4568), 
	.B2(n568), 
	.B1(\ram[249][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n417));
   AO22CHD U5994 (.O(n4569), 
	.B2(n568), 
	.B1(\ram[249][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n417));
   AO22CHD U5995 (.O(n4570), 
	.B2(n568), 
	.B1(\ram[249][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n417));
   AO22CHD U5996 (.O(n4571), 
	.B2(n568), 
	.B1(\ram[249][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n417));
   AO22CHD U5997 (.O(n4572), 
	.B2(n568), 
	.B1(\ram[249][6] ), 
	.A2(n14), 
	.A1(n417));
   AO22CHD U5998 (.O(n4573), 
	.B2(n568), 
	.B1(\ram[249][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n417));
   AO22CHD U5999 (.O(n4574), 
	.B2(n568), 
	.B1(\ram[249][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n417));
   AO22CHD U6000 (.O(n4575), 
	.B2(n568), 
	.B1(\ram[249][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n417));
   AO22CHD U6001 (.O(n4576), 
	.B2(n568), 
	.B1(\ram[249][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n417));
   AO22CHD U6002 (.O(n4577), 
	.B2(n568), 
	.B1(\ram[249][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n417));
   AO22CHD U6003 (.O(n4578), 
	.B2(n568), 
	.B1(\ram[249][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n417));
   AO22CHD U6004 (.O(n4579), 
	.B2(n568), 
	.B1(\ram[249][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n417));
   AO22CHD U6005 (.O(n4580), 
	.B2(n568), 
	.B1(\ram[249][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n417));
   AO22CHD U6006 (.O(n4581), 
	.B2(n568), 
	.B1(\ram[249][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n417));
   AO22CHD U6007 (.O(n4582), 
	.B2(n570), 
	.B1(\ram[250][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n419));
   AO22CHD U6008 (.O(n4583), 
	.B2(n570), 
	.B1(\ram[250][1] ), 
	.A2(n9), 
	.A1(n419));
   AO22CHD U6009 (.O(n4584), 
	.B2(n570), 
	.B1(\ram[250][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n419));
   AO22CHD U6010 (.O(n4585), 
	.B2(n570), 
	.B1(\ram[250][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n419));
   AO22CHD U6011 (.O(n4586), 
	.B2(n570), 
	.B1(\ram[250][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n419));
   AO22CHD U6012 (.O(n4587), 
	.B2(n570), 
	.B1(\ram[250][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n419));
   AO22CHD U6013 (.O(n4588), 
	.B2(n570), 
	.B1(\ram[250][6] ), 
	.A2(n14), 
	.A1(n419));
   AO22CHD U6014 (.O(n4589), 
	.B2(n570), 
	.B1(\ram[250][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n419));
   AO22CHD U6015 (.O(n4590), 
	.B2(n570), 
	.B1(\ram[250][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n419));
   AO22CHD U6016 (.O(n4591), 
	.B2(n570), 
	.B1(\ram[250][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n419));
   AO22CHD U6017 (.O(n4592), 
	.B2(n570), 
	.B1(\ram[250][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n419));
   AO22CHD U6018 (.O(n4593), 
	.B2(n570), 
	.B1(\ram[250][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n419));
   AO22CHD U6019 (.O(n4594), 
	.B2(n570), 
	.B1(\ram[250][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n419));
   AO22CHD U6020 (.O(n4595), 
	.B2(n570), 
	.B1(\ram[250][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n419));
   AO22CHD U6021 (.O(n4596), 
	.B2(n570), 
	.B1(\ram[250][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n419));
   AO22CHD U6022 (.O(n4597), 
	.B2(n570), 
	.B1(\ram[250][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n419));
   AO22CHD U6023 (.O(n4598), 
	.B2(n572), 
	.B1(\ram[251][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n421));
   AO22CHD U6024 (.O(n4599), 
	.B2(n572), 
	.B1(\ram[251][1] ), 
	.A2(n9), 
	.A1(n421));
   AO22CHD U6025 (.O(n4600), 
	.B2(n572), 
	.B1(\ram[251][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n421));
   AO22CHD U6026 (.O(n4601), 
	.B2(n572), 
	.B1(\ram[251][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n421));
   AO22CHD U6027 (.O(n4602), 
	.B2(n572), 
	.B1(\ram[251][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n421));
   AO22CHD U6028 (.O(n4603), 
	.B2(n572), 
	.B1(\ram[251][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n421));
   AO22CHD U6029 (.O(n4604), 
	.B2(n572), 
	.B1(\ram[251][6] ), 
	.A2(n14), 
	.A1(n421));
   AO22CHD U6030 (.O(n4605), 
	.B2(n572), 
	.B1(\ram[251][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n421));
   AO22CHD U6031 (.O(n4606), 
	.B2(n572), 
	.B1(\ram[251][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n421));
   AO22CHD U6032 (.O(n4607), 
	.B2(n572), 
	.B1(\ram[251][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n421));
   AO22CHD U6033 (.O(n4608), 
	.B2(n572), 
	.B1(\ram[251][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n421));
   AO22CHD U6034 (.O(n4609), 
	.B2(n572), 
	.B1(\ram[251][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n421));
   AO22CHD U6035 (.O(n4610), 
	.B2(n572), 
	.B1(\ram[251][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n421));
   AO22CHD U6036 (.O(n4611), 
	.B2(n572), 
	.B1(\ram[251][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n421));
   AO22CHD U6037 (.O(n4612), 
	.B2(n572), 
	.B1(\ram[251][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n421));
   AO22CHD U6038 (.O(n4613), 
	.B2(n572), 
	.B1(\ram[251][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n421));
   AO22CHD U6039 (.O(n4614), 
	.B2(n574), 
	.B1(\ram[252][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n423));
   AO22CHD U6040 (.O(n4615), 
	.B2(n574), 
	.B1(\ram[252][1] ), 
	.A2(n9), 
	.A1(n423));
   AO22CHD U6041 (.O(n4616), 
	.B2(n574), 
	.B1(\ram[252][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n423));
   AO22CHD U6042 (.O(n4617), 
	.B2(n574), 
	.B1(\ram[252][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n423));
   AO22CHD U6043 (.O(n4618), 
	.B2(n574), 
	.B1(\ram[252][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n423));
   AO22CHD U6044 (.O(n4619), 
	.B2(n574), 
	.B1(\ram[252][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n423));
   AO22CHD U6045 (.O(n4620), 
	.B2(n574), 
	.B1(\ram[252][6] ), 
	.A2(n14), 
	.A1(n423));
   AO22CHD U6046 (.O(n4621), 
	.B2(n574), 
	.B1(\ram[252][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n423));
   AO22CHD U6047 (.O(n4622), 
	.B2(n574), 
	.B1(\ram[252][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n423));
   AO22CHD U6048 (.O(n4623), 
	.B2(n574), 
	.B1(\ram[252][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n423));
   AO22CHD U6049 (.O(n4624), 
	.B2(n574), 
	.B1(\ram[252][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n423));
   AO22CHD U6050 (.O(n4625), 
	.B2(n574), 
	.B1(\ram[252][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n423));
   AO22CHD U6051 (.O(n4626), 
	.B2(n574), 
	.B1(\ram[252][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n423));
   AO22CHD U6052 (.O(n4627), 
	.B2(n574), 
	.B1(\ram[252][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n423));
   AO22CHD U6053 (.O(n4628), 
	.B2(n574), 
	.B1(\ram[252][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n423));
   AO22CHD U6054 (.O(n4629), 
	.B2(n574), 
	.B1(\ram[252][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n423));
   AO22CHD U6055 (.O(n4630), 
	.B2(n577), 
	.B1(\ram[253][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n425));
   AO22CHD U6056 (.O(n4631), 
	.B2(n577), 
	.B1(\ram[253][1] ), 
	.A2(n9), 
	.A1(n425));
   AO22CHD U6057 (.O(n4632), 
	.B2(n577), 
	.B1(\ram[253][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n425));
   AO22CHD U6058 (.O(n4633), 
	.B2(n577), 
	.B1(\ram[253][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n425));
   AO22CHD U6059 (.O(n4634), 
	.B2(n577), 
	.B1(\ram[253][4] ), 
	.A2(n12), 
	.A1(n425));
   AO22CHD U6060 (.O(n4635), 
	.B2(n577), 
	.B1(\ram[253][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n425));
   AO22CHD U6061 (.O(n4636), 
	.B2(n577), 
	.B1(\ram[253][6] ), 
	.A2(n14), 
	.A1(n425));
   AO22CHD U6062 (.O(n4637), 
	.B2(n577), 
	.B1(\ram[253][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n425));
   AO22CHD U6063 (.O(n4638), 
	.B2(n577), 
	.B1(\ram[253][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n425));
   AO22CHD U6064 (.O(n4639), 
	.B2(n577), 
	.B1(\ram[253][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n425));
   AO22CHD U6065 (.O(n4640), 
	.B2(n577), 
	.B1(\ram[253][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n425));
   AO22CHD U6066 (.O(n4641), 
	.B2(n577), 
	.B1(\ram[253][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n425));
   AO22CHD U6067 (.O(n4642), 
	.B2(n577), 
	.B1(\ram[253][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n425));
   AO22CHD U6068 (.O(n4643), 
	.B2(n577), 
	.B1(\ram[253][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n425));
   AO22CHD U6069 (.O(n4644), 
	.B2(n577), 
	.B1(\ram[253][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n425));
   AO22CHD U6070 (.O(n4645), 
	.B2(n577), 
	.B1(\ram[253][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n425));
   AO22CHD U6071 (.O(n4646), 
	.B2(n579), 
	.B1(\ram[254][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n427));
   AO22CHD U6072 (.O(n4647), 
	.B2(n579), 
	.B1(\ram[254][1] ), 
	.A2(n9), 
	.A1(n427));
   AO22CHD U6073 (.O(n4648), 
	.B2(n579), 
	.B1(\ram[254][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n427));
   AO22CHD U6074 (.O(n4649), 
	.B2(n579), 
	.B1(\ram[254][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n427));
   AO22CHD U6075 (.O(n4650), 
	.B2(n579), 
	.B1(\ram[254][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n427));
   AO22CHD U6076 (.O(n4651), 
	.B2(n579), 
	.B1(\ram[254][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n427));
   AO22CHD U6077 (.O(n4652), 
	.B2(n579), 
	.B1(\ram[254][6] ), 
	.A2(n14), 
	.A1(n427));
   AO22CHD U6078 (.O(n4653), 
	.B2(n579), 
	.B1(\ram[254][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n427));
   AO22CHD U6079 (.O(n4654), 
	.B2(n579), 
	.B1(\ram[254][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n427));
   AO22CHD U6080 (.O(n4655), 
	.B2(n579), 
	.B1(\ram[254][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n427));
   AO22CHD U6081 (.O(n4656), 
	.B2(n579), 
	.B1(\ram[254][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n427));
   AO22CHD U6082 (.O(n4657), 
	.B2(n579), 
	.B1(\ram[254][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n427));
   AO22CHD U6083 (.O(n4658), 
	.B2(n579), 
	.B1(\ram[254][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n427));
   AO22CHD U6084 (.O(n4659), 
	.B2(n579), 
	.B1(\ram[254][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n427));
   AO22CHD U6085 (.O(n4660), 
	.B2(n579), 
	.B1(\ram[254][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n427));
   AO22CHD U6086 (.O(n4661), 
	.B2(n579), 
	.B1(\ram[254][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n427));
   AO22CHD U6087 (.O(n4662), 
	.B2(n581), 
	.B1(\ram[255][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n429));
   AO22CHD U6088 (.O(n4663), 
	.B2(n581), 
	.B1(\ram[255][1] ), 
	.A2(n9), 
	.A1(n429));
   AO22CHD U6089 (.O(n4664), 
	.B2(n581), 
	.B1(\ram[255][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n429));
   AO22CHD U6090 (.O(n4665), 
	.B2(n581), 
	.B1(\ram[255][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n429));
   AO22CHD U6091 (.O(n4666), 
	.B2(n581), 
	.B1(\ram[255][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n429));
   AO22CHD U6092 (.O(n4667), 
	.B2(n581), 
	.B1(\ram[255][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n429));
   AO22CHD U6093 (.O(n4668), 
	.B2(n581), 
	.B1(\ram[255][6] ), 
	.A2(n14), 
	.A1(n429));
   AO22CHD U6094 (.O(n4669), 
	.B2(n581), 
	.B1(\ram[255][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n429));
   AO22CHD U6095 (.O(n4670), 
	.B2(n581), 
	.B1(\ram[255][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n429));
   AO22CHD U6096 (.O(n4671), 
	.B2(n581), 
	.B1(\ram[255][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n429));
   AO22CHD U6097 (.O(n4672), 
	.B2(n581), 
	.B1(\ram[255][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n429));
   AO22CHD U6098 (.O(n4673), 
	.B2(n581), 
	.B1(\ram[255][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n429));
   AO22CHD U6099 (.O(n4674), 
	.B2(n581), 
	.B1(\ram[255][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n429));
   AO22CHD U6100 (.O(n4675), 
	.B2(n581), 
	.B1(\ram[255][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n429));
   AO22CHD U6101 (.O(n4676), 
	.B2(n581), 
	.B1(\ram[255][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n429));
   AO22CHD U6102 (.O(n4677), 
	.B2(n581), 
	.B1(\ram[255][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n429));
   AO22CHD U6103 (.O(n582), 
	.B2(n8), 
	.B1(\ram[0][0] ), 
	.A2(n433), 
	.A1(n6));
   AO22CHD U6104 (.O(n583), 
	.B2(n8), 
	.B1(\ram[0][1] ), 
	.A2(n433), 
	.A1(FE_OFN46_n9));
   AO22CHD U6105 (.O(n584), 
	.B2(n8), 
	.B1(\ram[0][2] ), 
	.A2(n433), 
	.A1(FE_OFN49_n10));
   AO22CHD U6106 (.O(n585), 
	.B2(n8), 
	.B1(\ram[0][3] ), 
	.A2(n433), 
	.A1(FE_OFN52_n11));
   AO22CHD U6107 (.O(n586), 
	.B2(n8), 
	.B1(\ram[0][4] ), 
	.A2(n433), 
	.A1(FE_OFN55_n12));
   AO22CHD U6108 (.O(n587), 
	.B2(n8), 
	.B1(\ram[0][5] ), 
	.A2(n433), 
	.A1(FE_OFN58_n13));
   AO22CHD U6109 (.O(n588), 
	.B2(n8), 
	.B1(\ram[0][6] ), 
	.A2(n433), 
	.A1(FE_OFN62_n14));
   AO22CHD U6110 (.O(n589), 
	.B2(n8), 
	.B1(\ram[0][7] ), 
	.A2(n433), 
	.A1(FE_OFN63_n15));
   AO22CHD U6111 (.O(n590), 
	.B2(n8), 
	.B1(\ram[0][8] ), 
	.A2(n433), 
	.A1(FE_OFN68_n16));
   AO22CHD U6112 (.O(n591), 
	.B2(n8), 
	.B1(\ram[0][9] ), 
	.A2(n433), 
	.A1(FE_OFN70_n17));
   AO22CHD U6113 (.O(n592), 
	.B2(n8), 
	.B1(\ram[0][10] ), 
	.A2(n433), 
	.A1(FE_OFN73_n18));
   AO22CHD U6114 (.O(n593), 
	.B2(n8), 
	.B1(\ram[0][11] ), 
	.A2(n433), 
	.A1(FE_OFN76_n19));
   AO22CHD U6115 (.O(n594), 
	.B2(n8), 
	.B1(\ram[0][12] ), 
	.A2(n433), 
	.A1(FE_OFN80_n20));
   AO22CHD U6116 (.O(n595), 
	.B2(n8), 
	.B1(\ram[0][13] ), 
	.A2(n433), 
	.A1(FE_OFN85_n21));
   AO22CHD U6117 (.O(n596), 
	.B2(n8), 
	.B1(\ram[0][14] ), 
	.A2(n433), 
	.A1(n22));
   AO22CHD U6118 (.O(n597), 
	.B2(n8), 
	.B1(\ram[0][15] ), 
	.A2(n433), 
	.A1(FE_OFN91_n23));
   MUX4EHD U6119 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n571), 
	.D(\ram[255][0] ), 
	.C(\ram[253][0] ), 
	.B(\ram[254][0] ), 
	.A(\ram[252][0] ));
   MUX4EHD U6120 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n573), 
	.D(\ram[251][0] ), 
	.C(\ram[249][0] ), 
	.B(\ram[250][0] ), 
	.A(\ram[248][0] ));
   MUX4EHD U6121 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n576), 
	.D(\ram[247][0] ), 
	.C(\ram[245][0] ), 
	.B(\ram[246][0] ), 
	.A(\ram[244][0] ));
   MUX4EHD U6122 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n578), 
	.D(\ram[243][0] ), 
	.C(\ram[241][0] ), 
	.B(\ram[242][0] ), 
	.A(\ram[240][0] ));
   MUX4EHD U6123 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n580), 
	.D(n571), 
	.C(n576), 
	.B(n573), 
	.A(n578));
   MUX4EHD U6124 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4678), 
	.D(\ram[239][0] ), 
	.C(\ram[237][0] ), 
	.B(\ram[238][0] ), 
	.A(\ram[236][0] ));
   MUX4EHD U6125 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4679), 
	.D(\ram[235][0] ), 
	.C(\ram[233][0] ), 
	.B(\ram[234][0] ), 
	.A(\ram[232][0] ));
   MUX4EHD U6126 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4680), 
	.D(\ram[231][0] ), 
	.C(\ram[229][0] ), 
	.B(\ram[230][0] ), 
	.A(\ram[228][0] ));
   MUX4EHD U6127 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4681), 
	.D(\ram[227][0] ), 
	.C(\ram[225][0] ), 
	.B(\ram[226][0] ), 
	.A(\ram[224][0] ));
   MUX4EHD U6128 (.S1(n6136), 
	.S0(n7442), 
	.O(n4682), 
	.D(n4678), 
	.C(n4680), 
	.B(n4679), 
	.A(n4681));
   MUX4EHD U6129 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4683), 
	.D(\ram[223][0] ), 
	.C(\ram[221][0] ), 
	.B(\ram[222][0] ), 
	.A(\ram[220][0] ));
   MUX4EHD U6130 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4684), 
	.D(\ram[219][0] ), 
	.C(\ram[217][0] ), 
	.B(\ram[218][0] ), 
	.A(\ram[216][0] ));
   MUX4EHD U6131 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4685), 
	.D(\ram[215][0] ), 
	.C(\ram[213][0] ), 
	.B(\ram[214][0] ), 
	.A(\ram[212][0] ));
   MUX4EHD U6132 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4686), 
	.D(\ram[211][0] ), 
	.C(\ram[209][0] ), 
	.B(\ram[210][0] ), 
	.A(\ram[208][0] ));
   MUX4EHD U6133 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4687), 
	.D(n4683), 
	.C(n4685), 
	.B(n4684), 
	.A(n4686));
   MUX4EHD U6134 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4688), 
	.D(\ram[207][0] ), 
	.C(\ram[205][0] ), 
	.B(\ram[206][0] ), 
	.A(\ram[204][0] ));
   MUX4EHD U6135 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4689), 
	.D(\ram[203][0] ), 
	.C(\ram[201][0] ), 
	.B(\ram[202][0] ), 
	.A(\ram[200][0] ));
   MUX4EHD U6136 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4690), 
	.D(\ram[199][0] ), 
	.C(\ram[197][0] ), 
	.B(\ram[198][0] ), 
	.A(\ram[196][0] ));
   MUX4EHD U6137 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4691), 
	.D(\ram[195][0] ), 
	.C(\ram[193][0] ), 
	.B(\ram[194][0] ), 
	.A(\ram[192][0] ));
   MUX4EHD U6138 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4692), 
	.D(n4688), 
	.C(n4690), 
	.B(n4689), 
	.A(n4691));
   MUX4EHD U6139 (.S1(n6038), 
	.S0(n7444), 
	.O(n4693), 
	.D(n580), 
	.C(n4687), 
	.B(n4682), 
	.A(n4692));
   MUX4EHD U6140 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4694), 
	.D(\ram[191][0] ), 
	.C(\ram[189][0] ), 
	.B(\ram[190][0] ), 
	.A(\ram[188][0] ));
   MUX4EHD U6141 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4695), 
	.D(\ram[187][0] ), 
	.C(\ram[185][0] ), 
	.B(\ram[186][0] ), 
	.A(\ram[184][0] ));
   MUX4EHD U6142 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4696), 
	.D(\ram[183][0] ), 
	.C(\ram[181][0] ), 
	.B(\ram[182][0] ), 
	.A(\ram[180][0] ));
   MUX4EHD U6143 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4697), 
	.D(\ram[179][0] ), 
	.C(\ram[177][0] ), 
	.B(\ram[178][0] ), 
	.A(\ram[176][0] ));
   MUX4EHD U6144 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4698), 
	.D(n4694), 
	.C(n4696), 
	.B(n4695), 
	.A(n4697));
   MUX4EHD U6145 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4699), 
	.D(\ram[175][0] ), 
	.C(\ram[173][0] ), 
	.B(\ram[174][0] ), 
	.A(\ram[172][0] ));
   MUX4EHD U6146 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4700), 
	.D(\ram[171][0] ), 
	.C(\ram[169][0] ), 
	.B(\ram[170][0] ), 
	.A(\ram[168][0] ));
   MUX4EHD U6147 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4701), 
	.D(\ram[167][0] ), 
	.C(\ram[165][0] ), 
	.B(\ram[166][0] ), 
	.A(\ram[164][0] ));
   MUX4EHD U6148 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4702), 
	.D(\ram[163][0] ), 
	.C(\ram[161][0] ), 
	.B(\ram[162][0] ), 
	.A(\ram[160][0] ));
   MUX4EHD U6149 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4703), 
	.D(n4699), 
	.C(n4701), 
	.B(n4700), 
	.A(n4702));
   MUX4EHD U6150 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4704), 
	.D(\ram[159][0] ), 
	.C(\ram[157][0] ), 
	.B(\ram[158][0] ), 
	.A(\ram[156][0] ));
   MUX4EHD U6151 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4705), 
	.D(\ram[155][0] ), 
	.C(\ram[153][0] ), 
	.B(\ram[154][0] ), 
	.A(\ram[152][0] ));
   MUX4EHD U6152 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4706), 
	.D(\ram[151][0] ), 
	.C(\ram[149][0] ), 
	.B(\ram[150][0] ), 
	.A(\ram[148][0] ));
   MUX4EHD U6153 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4707), 
	.D(\ram[147][0] ), 
	.C(\ram[145][0] ), 
	.B(\ram[146][0] ), 
	.A(\ram[144][0] ));
   MUX4EHD U6154 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4708), 
	.D(n4704), 
	.C(n4706), 
	.B(n4705), 
	.A(n4707));
   MUX4EHD U6155 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4709), 
	.D(\ram[143][0] ), 
	.C(\ram[141][0] ), 
	.B(\ram[142][0] ), 
	.A(\ram[140][0] ));
   MUX4EHD U6156 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4710), 
	.D(\ram[139][0] ), 
	.C(\ram[137][0] ), 
	.B(\ram[138][0] ), 
	.A(\ram[136][0] ));
   MUX4EHD U6157 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4711), 
	.D(\ram[135][0] ), 
	.C(\ram[133][0] ), 
	.B(\ram[134][0] ), 
	.A(\ram[132][0] ));
   MUX4EHD U6158 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4712), 
	.D(\ram[131][0] ), 
	.C(\ram[129][0] ), 
	.B(\ram[130][0] ), 
	.A(\ram[128][0] ));
   MUX4EHD U6159 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4713), 
	.D(n4709), 
	.C(n4711), 
	.B(n4710), 
	.A(n4712));
   MUX4EHD U6160 (.S1(n6038), 
	.S0(n7444), 
	.O(n4714), 
	.D(n4698), 
	.C(n4708), 
	.B(n4703), 
	.A(n4713));
   MUX4EHD U6161 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4715), 
	.D(\ram[127][0] ), 
	.C(\ram[125][0] ), 
	.B(\ram[126][0] ), 
	.A(\ram[124][0] ));
   MUX4EHD U6162 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4716), 
	.D(\ram[123][0] ), 
	.C(\ram[121][0] ), 
	.B(\ram[122][0] ), 
	.A(\ram[120][0] ));
   MUX4EHD U6163 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4717), 
	.D(\ram[119][0] ), 
	.C(\ram[117][0] ), 
	.B(\ram[118][0] ), 
	.A(\ram[116][0] ));
   MUX4EHD U6164 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4718), 
	.D(\ram[115][0] ), 
	.C(\ram[113][0] ), 
	.B(\ram[114][0] ), 
	.A(\ram[112][0] ));
   MUX4EHD U6165 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4719), 
	.D(n4715), 
	.C(n4717), 
	.B(n4716), 
	.A(n4718));
   MUX4EHD U6166 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4720), 
	.D(\ram[111][0] ), 
	.C(\ram[109][0] ), 
	.B(\ram[110][0] ), 
	.A(\ram[108][0] ));
   MUX4EHD U6167 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4721), 
	.D(\ram[107][0] ), 
	.C(\ram[105][0] ), 
	.B(\ram[106][0] ), 
	.A(\ram[104][0] ));
   MUX4EHD U6168 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4722), 
	.D(\ram[103][0] ), 
	.C(\ram[101][0] ), 
	.B(\ram[102][0] ), 
	.A(\ram[100][0] ));
   MUX4EHD U6169 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4723), 
	.D(\ram[99][0] ), 
	.C(\ram[97][0] ), 
	.B(\ram[98][0] ), 
	.A(\ram[96][0] ));
   MUX4EHD U6170 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4724), 
	.D(n4720), 
	.C(n4722), 
	.B(n4721), 
	.A(n4723));
   MUX4EHD U6171 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4725), 
	.D(\ram[95][0] ), 
	.C(\ram[93][0] ), 
	.B(\ram[94][0] ), 
	.A(\ram[92][0] ));
   MUX4EHD U6172 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4726), 
	.D(\ram[91][0] ), 
	.C(\ram[89][0] ), 
	.B(\ram[90][0] ), 
	.A(\ram[88][0] ));
   MUX4EHD U6173 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4727), 
	.D(\ram[87][0] ), 
	.C(\ram[85][0] ), 
	.B(\ram[86][0] ), 
	.A(\ram[84][0] ));
   MUX4EHD U6174 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4728), 
	.D(\ram[83][0] ), 
	.C(\ram[81][0] ), 
	.B(\ram[82][0] ), 
	.A(\ram[80][0] ));
   MUX4EHD U6175 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4729), 
	.D(n4725), 
	.C(n4727), 
	.B(n4726), 
	.A(n4728));
   MUX4EHD U6176 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4730), 
	.D(\ram[79][0] ), 
	.C(\ram[77][0] ), 
	.B(\ram[78][0] ), 
	.A(\ram[76][0] ));
   MUX4EHD U6177 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4731), 
	.D(\ram[75][0] ), 
	.C(\ram[73][0] ), 
	.B(\ram[74][0] ), 
	.A(\ram[72][0] ));
   MUX4EHD U6178 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4732), 
	.D(\ram[71][0] ), 
	.C(\ram[69][0] ), 
	.B(\ram[70][0] ), 
	.A(\ram[68][0] ));
   MUX4EHD U6179 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4733), 
	.D(\ram[67][0] ), 
	.C(\ram[65][0] ), 
	.B(\ram[66][0] ), 
	.A(\ram[64][0] ));
   MUX4EHD U6180 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4734), 
	.D(n4730), 
	.C(n4732), 
	.B(n4731), 
	.A(n4733));
   MUX4EHD U6181 (.S1(n6038), 
	.S0(n7444), 
	.O(n4735), 
	.D(n4719), 
	.C(n4729), 
	.B(n4724), 
	.A(n4734));
   MUX4EHD U6182 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4736), 
	.D(\ram[63][0] ), 
	.C(\ram[61][0] ), 
	.B(\ram[62][0] ), 
	.A(\ram[60][0] ));
   MUX4EHD U6183 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4737), 
	.D(\ram[59][0] ), 
	.C(\ram[57][0] ), 
	.B(\ram[58][0] ), 
	.A(\ram[56][0] ));
   MUX4EHD U6184 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4738), 
	.D(\ram[55][0] ), 
	.C(\ram[53][0] ), 
	.B(\ram[54][0] ), 
	.A(\ram[52][0] ));
   MUX4EHD U6185 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4739), 
	.D(\ram[51][0] ), 
	.C(\ram[49][0] ), 
	.B(\ram[50][0] ), 
	.A(\ram[48][0] ));
   MUX4EHD U6186 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4740), 
	.D(n4736), 
	.C(n4738), 
	.B(n4737), 
	.A(n4739));
   MUX4EHD U6187 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4741), 
	.D(\ram[47][0] ), 
	.C(\ram[45][0] ), 
	.B(\ram[46][0] ), 
	.A(\ram[44][0] ));
   MUX4EHD U6188 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4742), 
	.D(\ram[43][0] ), 
	.C(\ram[41][0] ), 
	.B(\ram[42][0] ), 
	.A(\ram[40][0] ));
   MUX4EHD U6189 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4743), 
	.D(\ram[39][0] ), 
	.C(\ram[37][0] ), 
	.B(\ram[38][0] ), 
	.A(\ram[36][0] ));
   MUX4EHD U6190 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4744), 
	.D(\ram[35][0] ), 
	.C(\ram[33][0] ), 
	.B(\ram[34][0] ), 
	.A(\ram[32][0] ));
   MUX4EHD U6191 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4745), 
	.D(n4741), 
	.C(n4743), 
	.B(n4742), 
	.A(n4744));
   MUX4EHD U6192 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4746), 
	.D(\ram[31][0] ), 
	.C(\ram[29][0] ), 
	.B(\ram[30][0] ), 
	.A(\ram[28][0] ));
   MUX4EHD U6193 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4747), 
	.D(\ram[27][0] ), 
	.C(\ram[25][0] ), 
	.B(\ram[26][0] ), 
	.A(\ram[24][0] ));
   MUX4EHD U6194 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4748), 
	.D(\ram[23][0] ), 
	.C(\ram[21][0] ), 
	.B(\ram[22][0] ), 
	.A(\ram[20][0] ));
   MUX4EHD U6195 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4749), 
	.D(\ram[19][0] ), 
	.C(\ram[17][0] ), 
	.B(\ram[18][0] ), 
	.A(\ram[16][0] ));
   MUX4EHD U6196 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4750), 
	.D(n4746), 
	.C(n4748), 
	.B(n4747), 
	.A(n4749));
   MUX4EHD U6197 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4751), 
	.D(\ram[15][0] ), 
	.C(\ram[13][0] ), 
	.B(\ram[14][0] ), 
	.A(\ram[12][0] ));
   MUX4EHD U6198 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4752), 
	.D(\ram[11][0] ), 
	.C(\ram[9][0] ), 
	.B(\ram[10][0] ), 
	.A(\ram[8][0] ));
   MUX4EHD U6199 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4753), 
	.D(\ram[7][0] ), 
	.C(\ram[5][0] ), 
	.B(\ram[6][0] ), 
	.A(\ram[4][0] ));
   MUX4EHD U6200 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4754), 
	.D(\ram[3][0] ), 
	.C(\ram[1][0] ), 
	.B(\ram[2][0] ), 
	.A(\ram[0][0] ));
   MUX4EHD U6201 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4755), 
	.D(n4751), 
	.C(n4753), 
	.B(n4752), 
	.A(n4754));
   MUX4EHD U6202 (.S1(n6038), 
	.S0(n7444), 
	.O(n4756), 
	.D(n4740), 
	.C(n4750), 
	.B(n4745), 
	.A(n4755));
   MUX4EHD U6203 (.S1(n6469), 
	.S0(n6470), 
	.O(N4141), 
	.D(n4693), 
	.C(n4735), 
	.B(n4714), 
	.A(n4756));
   MUX4EHD U6204 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4757), 
	.D(\ram[255][1] ), 
	.C(\ram[253][1] ), 
	.B(\ram[254][1] ), 
	.A(\ram[252][1] ));
   MUX4EHD U6205 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4758), 
	.D(\ram[251][1] ), 
	.C(\ram[249][1] ), 
	.B(\ram[250][1] ), 
	.A(\ram[248][1] ));
   MUX4EHD U6206 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4759), 
	.D(\ram[247][1] ), 
	.C(\ram[245][1] ), 
	.B(\ram[246][1] ), 
	.A(\ram[244][1] ));
   MUX4EHD U6207 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4760), 
	.D(\ram[243][1] ), 
	.C(\ram[241][1] ), 
	.B(\ram[242][1] ), 
	.A(\ram[240][1] ));
   MUX4EHD U6208 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4761), 
	.D(n4757), 
	.C(n4759), 
	.B(n4758), 
	.A(n4760));
   MUX4EHD U6209 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4762), 
	.D(\ram[239][1] ), 
	.C(\ram[237][1] ), 
	.B(\ram[238][1] ), 
	.A(\ram[236][1] ));
   MUX4EHD U6210 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4763), 
	.D(\ram[235][1] ), 
	.C(\ram[233][1] ), 
	.B(\ram[234][1] ), 
	.A(\ram[232][1] ));
   MUX4EHD U6211 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4764), 
	.D(\ram[231][1] ), 
	.C(\ram[229][1] ), 
	.B(\ram[230][1] ), 
	.A(\ram[228][1] ));
   MUX4EHD U6212 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4765), 
	.D(\ram[227][1] ), 
	.C(\ram[225][1] ), 
	.B(\ram[226][1] ), 
	.A(\ram[224][1] ));
   MUX4EHD U6213 (.S1(n6136), 
	.S0(n7442), 
	.O(n4766), 
	.D(n4762), 
	.C(n4764), 
	.B(n4763), 
	.A(n4765));
   MUX4EHD U6214 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4767), 
	.D(\ram[223][1] ), 
	.C(\ram[221][1] ), 
	.B(\ram[222][1] ), 
	.A(\ram[220][1] ));
   MUX4EHD U6215 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4768), 
	.D(\ram[219][1] ), 
	.C(\ram[217][1] ), 
	.B(\ram[218][1] ), 
	.A(\ram[216][1] ));
   MUX4EHD U6216 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4769), 
	.D(\ram[215][1] ), 
	.C(\ram[213][1] ), 
	.B(\ram[214][1] ), 
	.A(\ram[212][1] ));
   MUX4EHD U6217 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4770), 
	.D(\ram[211][1] ), 
	.C(\ram[209][1] ), 
	.B(\ram[210][1] ), 
	.A(\ram[208][1] ));
   MUX4EHD U6218 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4771), 
	.D(n4767), 
	.C(n4769), 
	.B(n4768), 
	.A(n4770));
   MUX4EHD U6219 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4772), 
	.D(\ram[207][1] ), 
	.C(\ram[205][1] ), 
	.B(\ram[206][1] ), 
	.A(\ram[204][1] ));
   MUX4EHD U6220 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4773), 
	.D(\ram[203][1] ), 
	.C(\ram[201][1] ), 
	.B(\ram[202][1] ), 
	.A(\ram[200][1] ));
   MUX4EHD U6221 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4774), 
	.D(\ram[199][1] ), 
	.C(\ram[197][1] ), 
	.B(\ram[198][1] ), 
	.A(\ram[196][1] ));
   MUX4EHD U6222 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4775), 
	.D(\ram[195][1] ), 
	.C(\ram[193][1] ), 
	.B(\ram[194][1] ), 
	.A(\ram[192][1] ));
   MUX4EHD U6223 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4776), 
	.D(n4772), 
	.C(n4774), 
	.B(n4773), 
	.A(n4775));
   MUX4EHD U6224 (.S1(n6038), 
	.S0(n7444), 
	.O(n4777), 
	.D(n4761), 
	.C(n4771), 
	.B(n4766), 
	.A(n4776));
   MUX4EHD U6225 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4778), 
	.D(\ram[191][1] ), 
	.C(\ram[189][1] ), 
	.B(\ram[190][1] ), 
	.A(\ram[188][1] ));
   MUX4EHD U6226 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4779), 
	.D(\ram[187][1] ), 
	.C(\ram[185][1] ), 
	.B(\ram[186][1] ), 
	.A(\ram[184][1] ));
   MUX4EHD U6227 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4780), 
	.D(\ram[183][1] ), 
	.C(\ram[181][1] ), 
	.B(\ram[182][1] ), 
	.A(\ram[180][1] ));
   MUX4EHD U6228 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4781), 
	.D(\ram[179][1] ), 
	.C(\ram[177][1] ), 
	.B(\ram[178][1] ), 
	.A(\ram[176][1] ));
   MUX4EHD U6229 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4782), 
	.D(n4778), 
	.C(n4780), 
	.B(n4779), 
	.A(n4781));
   MUX4EHD U6230 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4783), 
	.D(\ram[175][1] ), 
	.C(\ram[173][1] ), 
	.B(\ram[174][1] ), 
	.A(\ram[172][1] ));
   MUX4EHD U6231 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4784), 
	.D(\ram[171][1] ), 
	.C(\ram[169][1] ), 
	.B(\ram[170][1] ), 
	.A(\ram[168][1] ));
   MUX4EHD U6232 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4785), 
	.D(\ram[167][1] ), 
	.C(\ram[165][1] ), 
	.B(\ram[166][1] ), 
	.A(\ram[164][1] ));
   MUX4EHD U6233 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4786), 
	.D(\ram[163][1] ), 
	.C(\ram[161][1] ), 
	.B(\ram[162][1] ), 
	.A(\ram[160][1] ));
   MUX4EHD U6234 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4787), 
	.D(n4783), 
	.C(n4785), 
	.B(n4784), 
	.A(n4786));
   MUX4EHD U6235 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4788), 
	.D(\ram[159][1] ), 
	.C(\ram[157][1] ), 
	.B(\ram[158][1] ), 
	.A(\ram[156][1] ));
   MUX4EHD U6236 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4789), 
	.D(\ram[155][1] ), 
	.C(\ram[153][1] ), 
	.B(\ram[154][1] ), 
	.A(\ram[152][1] ));
   MUX4EHD U6237 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4790), 
	.D(\ram[151][1] ), 
	.C(\ram[149][1] ), 
	.B(\ram[150][1] ), 
	.A(\ram[148][1] ));
   MUX4EHD U6238 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4791), 
	.D(\ram[147][1] ), 
	.C(\ram[145][1] ), 
	.B(\ram[146][1] ), 
	.A(\ram[144][1] ));
   MUX4EHD U6239 (.S1(n6136), 
	.S0(n7442), 
	.O(n4792), 
	.D(n4788), 
	.C(n4790), 
	.B(n4789), 
	.A(n4791));
   MUX4EHD U6240 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4793), 
	.D(\ram[143][1] ), 
	.C(\ram[141][1] ), 
	.B(\ram[142][1] ), 
	.A(\ram[140][1] ));
   MUX4EHD U6241 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4794), 
	.D(\ram[139][1] ), 
	.C(\ram[137][1] ), 
	.B(\ram[138][1] ), 
	.A(\ram[136][1] ));
   MUX4EHD U6242 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4795), 
	.D(\ram[135][1] ), 
	.C(\ram[133][1] ), 
	.B(\ram[134][1] ), 
	.A(\ram[132][1] ));
   MUX4EHD U6243 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4796), 
	.D(\ram[131][1] ), 
	.C(\ram[129][1] ), 
	.B(\ram[130][1] ), 
	.A(\ram[128][1] ));
   MUX4EHD U6244 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4797), 
	.D(n4793), 
	.C(n4795), 
	.B(n4794), 
	.A(n4796));
   MUX4EHD U6245 (.S1(n6038), 
	.S0(n7444), 
	.O(n4798), 
	.D(n4782), 
	.C(n4792), 
	.B(n4787), 
	.A(n4797));
   MUX4EHD U6246 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4799), 
	.D(\ram[127][1] ), 
	.C(\ram[125][1] ), 
	.B(\ram[126][1] ), 
	.A(\ram[124][1] ));
   MUX4EHD U6247 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4800), 
	.D(\ram[123][1] ), 
	.C(\ram[121][1] ), 
	.B(\ram[122][1] ), 
	.A(\ram[120][1] ));
   MUX4EHD U6248 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4801), 
	.D(\ram[119][1] ), 
	.C(\ram[117][1] ), 
	.B(\ram[118][1] ), 
	.A(\ram[116][1] ));
   MUX4EHD U6249 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4802), 
	.D(\ram[115][1] ), 
	.C(\ram[113][1] ), 
	.B(\ram[114][1] ), 
	.A(\ram[112][1] ));
   MUX4EHD U6250 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4803), 
	.D(n4799), 
	.C(n4801), 
	.B(n4800), 
	.A(n4802));
   MUX4EHD U6251 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4804), 
	.D(\ram[111][1] ), 
	.C(\ram[109][1] ), 
	.B(\ram[110][1] ), 
	.A(\ram[108][1] ));
   MUX4EHD U6252 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4805), 
	.D(\ram[107][1] ), 
	.C(\ram[105][1] ), 
	.B(\ram[106][1] ), 
	.A(\ram[104][1] ));
   MUX4EHD U6253 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4806), 
	.D(\ram[103][1] ), 
	.C(\ram[101][1] ), 
	.B(\ram[102][1] ), 
	.A(\ram[100][1] ));
   MUX4EHD U6254 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4807), 
	.D(\ram[99][1] ), 
	.C(\ram[97][1] ), 
	.B(\ram[98][1] ), 
	.A(\ram[96][1] ));
   MUX4EHD U6255 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4808), 
	.D(n4804), 
	.C(n4806), 
	.B(n4805), 
	.A(n4807));
   MUX4EHD U6256 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4809), 
	.D(\ram[95][1] ), 
	.C(\ram[93][1] ), 
	.B(\ram[94][1] ), 
	.A(\ram[92][1] ));
   MUX4EHD U6257 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4810), 
	.D(\ram[91][1] ), 
	.C(\ram[89][1] ), 
	.B(\ram[90][1] ), 
	.A(\ram[88][1] ));
   MUX4EHD U6258 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4811), 
	.D(\ram[87][1] ), 
	.C(\ram[85][1] ), 
	.B(\ram[86][1] ), 
	.A(\ram[84][1] ));
   MUX4EHD U6259 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4812), 
	.D(\ram[83][1] ), 
	.C(\ram[81][1] ), 
	.B(\ram[82][1] ), 
	.A(\ram[80][1] ));
   MUX4EHD U6260 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4813), 
	.D(n4809), 
	.C(n4811), 
	.B(n4810), 
	.A(n4812));
   MUX4EHD U6261 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4814), 
	.D(\ram[79][1] ), 
	.C(\ram[77][1] ), 
	.B(\ram[78][1] ), 
	.A(\ram[76][1] ));
   MUX4EHD U6262 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4815), 
	.D(\ram[75][1] ), 
	.C(\ram[73][1] ), 
	.B(\ram[74][1] ), 
	.A(\ram[72][1] ));
   MUX4EHD U6263 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4816), 
	.D(\ram[71][1] ), 
	.C(\ram[69][1] ), 
	.B(\ram[70][1] ), 
	.A(\ram[68][1] ));
   MUX4EHD U6264 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4817), 
	.D(\ram[67][1] ), 
	.C(\ram[65][1] ), 
	.B(\ram[66][1] ), 
	.A(\ram[64][1] ));
   MUX4EHD U6265 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4818), 
	.D(n4814), 
	.C(n4816), 
	.B(n4815), 
	.A(n4817));
   MUX4EHD U6266 (.S1(n6038), 
	.S0(n7444), 
	.O(n4819), 
	.D(n4803), 
	.C(n4813), 
	.B(n4808), 
	.A(n4818));
   MUX4EHD U6267 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4820), 
	.D(\ram[63][1] ), 
	.C(\ram[61][1] ), 
	.B(\ram[62][1] ), 
	.A(\ram[60][1] ));
   MUX4EHD U6268 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4821), 
	.D(\ram[59][1] ), 
	.C(\ram[57][1] ), 
	.B(\ram[58][1] ), 
	.A(\ram[56][1] ));
   MUX4EHD U6269 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4822), 
	.D(\ram[55][1] ), 
	.C(\ram[53][1] ), 
	.B(\ram[54][1] ), 
	.A(\ram[52][1] ));
   MUX4EHD U6270 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4823), 
	.D(\ram[51][1] ), 
	.C(\ram[49][1] ), 
	.B(\ram[50][1] ), 
	.A(\ram[48][1] ));
   MUX4EHD U6271 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4824), 
	.D(n4820), 
	.C(n4822), 
	.B(n4821), 
	.A(n4823));
   MUX4EHD U6272 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4825), 
	.D(\ram[47][1] ), 
	.C(\ram[45][1] ), 
	.B(\ram[46][1] ), 
	.A(\ram[44][1] ));
   MUX4EHD U6273 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4826), 
	.D(\ram[43][1] ), 
	.C(\ram[41][1] ), 
	.B(\ram[42][1] ), 
	.A(\ram[40][1] ));
   MUX4EHD U6274 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4827), 
	.D(\ram[39][1] ), 
	.C(\ram[37][1] ), 
	.B(\ram[38][1] ), 
	.A(\ram[36][1] ));
   MUX4EHD U6275 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4828), 
	.D(\ram[35][1] ), 
	.C(\ram[33][1] ), 
	.B(\ram[34][1] ), 
	.A(\ram[32][1] ));
   MUX4EHD U6276 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4829), 
	.D(n4825), 
	.C(n4827), 
	.B(n4826), 
	.A(n4828));
   MUX4EHD U6277 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4830), 
	.D(\ram[31][1] ), 
	.C(\ram[29][1] ), 
	.B(\ram[30][1] ), 
	.A(\ram[28][1] ));
   MUX4EHD U6278 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4831), 
	.D(\ram[27][1] ), 
	.C(\ram[25][1] ), 
	.B(\ram[26][1] ), 
	.A(\ram[24][1] ));
   MUX4EHD U6279 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4832), 
	.D(\ram[23][1] ), 
	.C(\ram[21][1] ), 
	.B(\ram[22][1] ), 
	.A(\ram[20][1] ));
   MUX4EHD U6280 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4833), 
	.D(\ram[19][1] ), 
	.C(\ram[17][1] ), 
	.B(\ram[18][1] ), 
	.A(\ram[16][1] ));
   MUX4EHD U6281 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4834), 
	.D(n4830), 
	.C(n4832), 
	.B(n4831), 
	.A(n4833));
   MUX4EHD U6282 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n4835), 
	.D(\ram[15][1] ), 
	.C(\ram[13][1] ), 
	.B(\ram[14][1] ), 
	.A(\ram[12][1] ));
   MUX4EHD U6283 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4836), 
	.D(\ram[11][1] ), 
	.C(\ram[9][1] ), 
	.B(\ram[10][1] ), 
	.A(\ram[8][1] ));
   MUX4EHD U6284 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4837), 
	.D(\ram[7][1] ), 
	.C(\ram[5][1] ), 
	.B(\ram[6][1] ), 
	.A(\ram[4][1] ));
   MUX4EHD U6285 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n4838), 
	.D(\ram[3][1] ), 
	.C(\ram[1][1] ), 
	.B(\ram[2][1] ), 
	.A(\ram[0][1] ));
   MUX4EHD U6286 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4839), 
	.D(n4835), 
	.C(n4837), 
	.B(n4836), 
	.A(n4838));
   MUX4EHD U6287 (.S1(n6038), 
	.S0(n7444), 
	.O(n4840), 
	.D(n4824), 
	.C(n4834), 
	.B(n4829), 
	.A(n4839));
   MUX4EHD U6288 (.S1(n6469), 
	.S0(n6470), 
	.O(N4140), 
	.D(n4777), 
	.C(n4819), 
	.B(n4798), 
	.A(n4840));
   MUX4EHD U6289 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4841), 
	.D(\ram[255][2] ), 
	.C(\ram[253][2] ), 
	.B(\ram[254][2] ), 
	.A(\ram[252][2] ));
   MUX4EHD U6290 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4842), 
	.D(\ram[251][2] ), 
	.C(\ram[249][2] ), 
	.B(\ram[250][2] ), 
	.A(\ram[248][2] ));
   MUX4EHD U6291 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4843), 
	.D(\ram[247][2] ), 
	.C(\ram[245][2] ), 
	.B(\ram[246][2] ), 
	.A(\ram[244][2] ));
   MUX4EHD U6292 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4844), 
	.D(\ram[243][2] ), 
	.C(\ram[241][2] ), 
	.B(\ram[242][2] ), 
	.A(\ram[240][2] ));
   MUX4EHD U6293 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4845), 
	.D(n4841), 
	.C(n4843), 
	.B(n4842), 
	.A(n4844));
   MUX4EHD U6294 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4846), 
	.D(\ram[239][2] ), 
	.C(\ram[237][2] ), 
	.B(\ram[238][2] ), 
	.A(\ram[236][2] ));
   MUX4EHD U6295 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4847), 
	.D(\ram[235][2] ), 
	.C(\ram[233][2] ), 
	.B(\ram[234][2] ), 
	.A(\ram[232][2] ));
   MUX4EHD U6296 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4848), 
	.D(\ram[231][2] ), 
	.C(\ram[229][2] ), 
	.B(\ram[230][2] ), 
	.A(\ram[228][2] ));
   MUX4EHD U6297 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4849), 
	.D(\ram[227][2] ), 
	.C(\ram[225][2] ), 
	.B(\ram[226][2] ), 
	.A(\ram[224][2] ));
   MUX4EHD U6298 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4850), 
	.D(n4846), 
	.C(n4848), 
	.B(n4847), 
	.A(n4849));
   MUX4EHD U6299 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4851), 
	.D(\ram[223][2] ), 
	.C(\ram[221][2] ), 
	.B(\ram[222][2] ), 
	.A(\ram[220][2] ));
   MUX4EHD U6300 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4852), 
	.D(\ram[219][2] ), 
	.C(\ram[217][2] ), 
	.B(\ram[218][2] ), 
	.A(\ram[216][2] ));
   MUX4EHD U6301 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4853), 
	.D(\ram[215][2] ), 
	.C(\ram[213][2] ), 
	.B(\ram[214][2] ), 
	.A(\ram[212][2] ));
   MUX4EHD U6302 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4854), 
	.D(\ram[211][2] ), 
	.C(\ram[209][2] ), 
	.B(\ram[210][2] ), 
	.A(\ram[208][2] ));
   MUX4EHD U6303 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4855), 
	.D(n4851), 
	.C(n4853), 
	.B(n4852), 
	.A(n4854));
   MUX4EHD U6304 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4856), 
	.D(\ram[207][2] ), 
	.C(\ram[205][2] ), 
	.B(\ram[206][2] ), 
	.A(\ram[204][2] ));
   MUX4EHD U6305 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4857), 
	.D(\ram[203][2] ), 
	.C(\ram[201][2] ), 
	.B(\ram[202][2] ), 
	.A(\ram[200][2] ));
   MUX4EHD U6306 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4858), 
	.D(\ram[199][2] ), 
	.C(\ram[197][2] ), 
	.B(\ram[198][2] ), 
	.A(\ram[196][2] ));
   MUX4EHD U6307 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4859), 
	.D(\ram[195][2] ), 
	.C(\ram[193][2] ), 
	.B(\ram[194][2] ), 
	.A(\ram[192][2] ));
   MUX4EHD U6308 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4860), 
	.D(n4856), 
	.C(n4858), 
	.B(n4857), 
	.A(n4859));
   MUX4EHD U6309 (.S1(n6038), 
	.S0(n7444), 
	.O(n4861), 
	.D(n4845), 
	.C(n4855), 
	.B(n4850), 
	.A(n4860));
   MUX4EHD U6310 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4862), 
	.D(\ram[191][2] ), 
	.C(\ram[189][2] ), 
	.B(\ram[190][2] ), 
	.A(\ram[188][2] ));
   MUX4EHD U6311 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4863), 
	.D(\ram[187][2] ), 
	.C(\ram[185][2] ), 
	.B(\ram[186][2] ), 
	.A(\ram[184][2] ));
   MUX4EHD U6312 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4864), 
	.D(\ram[183][2] ), 
	.C(\ram[181][2] ), 
	.B(\ram[182][2] ), 
	.A(\ram[180][2] ));
   MUX4EHD U6313 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4865), 
	.D(\ram[179][2] ), 
	.C(\ram[177][2] ), 
	.B(\ram[178][2] ), 
	.A(\ram[176][2] ));
   MUX4EHD U6314 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4866), 
	.D(n4862), 
	.C(n4864), 
	.B(n4863), 
	.A(n4865));
   MUX4EHD U6315 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4867), 
	.D(\ram[175][2] ), 
	.C(\ram[173][2] ), 
	.B(\ram[174][2] ), 
	.A(\ram[172][2] ));
   MUX4EHD U6316 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4868), 
	.D(\ram[171][2] ), 
	.C(\ram[169][2] ), 
	.B(\ram[170][2] ), 
	.A(\ram[168][2] ));
   MUX4EHD U6317 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4869), 
	.D(\ram[167][2] ), 
	.C(\ram[165][2] ), 
	.B(\ram[166][2] ), 
	.A(\ram[164][2] ));
   MUX4EHD U6318 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4870), 
	.D(\ram[163][2] ), 
	.C(\ram[161][2] ), 
	.B(\ram[162][2] ), 
	.A(\ram[160][2] ));
   MUX4EHD U6319 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4871), 
	.D(n4867), 
	.C(n4869), 
	.B(n4868), 
	.A(n4870));
   MUX4EHD U6320 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4872), 
	.D(\ram[159][2] ), 
	.C(\ram[157][2] ), 
	.B(\ram[158][2] ), 
	.A(\ram[156][2] ));
   MUX4EHD U6321 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4873), 
	.D(\ram[155][2] ), 
	.C(\ram[153][2] ), 
	.B(\ram[154][2] ), 
	.A(\ram[152][2] ));
   MUX4EHD U6322 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4874), 
	.D(\ram[151][2] ), 
	.C(\ram[149][2] ), 
	.B(\ram[150][2] ), 
	.A(\ram[148][2] ));
   MUX4EHD U6323 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4875), 
	.D(\ram[147][2] ), 
	.C(\ram[145][2] ), 
	.B(\ram[146][2] ), 
	.A(\ram[144][2] ));
   MUX4EHD U6324 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4876), 
	.D(n4872), 
	.C(n4874), 
	.B(n4873), 
	.A(n4875));
   MUX4EHD U6325 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4877), 
	.D(\ram[143][2] ), 
	.C(\ram[141][2] ), 
	.B(\ram[142][2] ), 
	.A(\ram[140][2] ));
   MUX4EHD U6326 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4878), 
	.D(\ram[139][2] ), 
	.C(\ram[137][2] ), 
	.B(\ram[138][2] ), 
	.A(\ram[136][2] ));
   MUX4EHD U6327 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4879), 
	.D(\ram[135][2] ), 
	.C(\ram[133][2] ), 
	.B(\ram[134][2] ), 
	.A(\ram[132][2] ));
   MUX4EHD U6328 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4880), 
	.D(\ram[131][2] ), 
	.C(\ram[129][2] ), 
	.B(\ram[130][2] ), 
	.A(\ram[128][2] ));
   MUX4EHD U6329 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4881), 
	.D(n4877), 
	.C(n4879), 
	.B(n4878), 
	.A(n4880));
   MUX4EHD U6330 (.S1(n6038), 
	.S0(n7444), 
	.O(n4882), 
	.D(n4866), 
	.C(n4876), 
	.B(n4871), 
	.A(n4881));
   MUX4EHD U6331 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4883), 
	.D(\ram[127][2] ), 
	.C(\ram[125][2] ), 
	.B(\ram[126][2] ), 
	.A(\ram[124][2] ));
   MUX4EHD U6332 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4884), 
	.D(\ram[123][2] ), 
	.C(\ram[121][2] ), 
	.B(\ram[122][2] ), 
	.A(\ram[120][2] ));
   MUX4EHD U6333 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4885), 
	.D(\ram[119][2] ), 
	.C(\ram[117][2] ), 
	.B(\ram[118][2] ), 
	.A(\ram[116][2] ));
   MUX4EHD U6334 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4886), 
	.D(\ram[115][2] ), 
	.C(\ram[113][2] ), 
	.B(\ram[114][2] ), 
	.A(\ram[112][2] ));
   MUX4EHD U6335 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4887), 
	.D(n4883), 
	.C(n4885), 
	.B(n4884), 
	.A(n4886));
   MUX4EHD U6336 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4888), 
	.D(\ram[111][2] ), 
	.C(\ram[109][2] ), 
	.B(\ram[110][2] ), 
	.A(\ram[108][2] ));
   MUX4EHD U6337 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4889), 
	.D(\ram[107][2] ), 
	.C(\ram[105][2] ), 
	.B(\ram[106][2] ), 
	.A(\ram[104][2] ));
   MUX4EHD U6338 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4890), 
	.D(\ram[103][2] ), 
	.C(\ram[101][2] ), 
	.B(\ram[102][2] ), 
	.A(\ram[100][2] ));
   MUX4EHD U6339 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4891), 
	.D(\ram[99][2] ), 
	.C(\ram[97][2] ), 
	.B(\ram[98][2] ), 
	.A(\ram[96][2] ));
   MUX4EHD U6340 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4892), 
	.D(n4888), 
	.C(n4890), 
	.B(n4889), 
	.A(n4891));
   MUX4EHD U6341 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4893), 
	.D(\ram[95][2] ), 
	.C(\ram[93][2] ), 
	.B(\ram[94][2] ), 
	.A(\ram[92][2] ));
   MUX4EHD U6342 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4894), 
	.D(\ram[91][2] ), 
	.C(\ram[89][2] ), 
	.B(\ram[90][2] ), 
	.A(\ram[88][2] ));
   MUX4EHD U6343 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4895), 
	.D(\ram[87][2] ), 
	.C(\ram[85][2] ), 
	.B(\ram[86][2] ), 
	.A(\ram[84][2] ));
   MUX4EHD U6344 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4896), 
	.D(\ram[83][2] ), 
	.C(\ram[81][2] ), 
	.B(\ram[82][2] ), 
	.A(\ram[80][2] ));
   MUX4EHD U6345 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4897), 
	.D(n4893), 
	.C(n4895), 
	.B(n4894), 
	.A(n4896));
   MUX4EHD U6346 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4898), 
	.D(\ram[79][2] ), 
	.C(\ram[77][2] ), 
	.B(\ram[78][2] ), 
	.A(\ram[76][2] ));
   MUX4EHD U6347 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4899), 
	.D(\ram[75][2] ), 
	.C(\ram[73][2] ), 
	.B(\ram[74][2] ), 
	.A(\ram[72][2] ));
   MUX4EHD U6348 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4900), 
	.D(\ram[71][2] ), 
	.C(\ram[69][2] ), 
	.B(\ram[70][2] ), 
	.A(\ram[68][2] ));
   MUX4EHD U6349 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4901), 
	.D(\ram[67][2] ), 
	.C(\ram[65][2] ), 
	.B(\ram[66][2] ), 
	.A(\ram[64][2] ));
   MUX4EHD U6350 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4902), 
	.D(n4898), 
	.C(n4900), 
	.B(n4899), 
	.A(n4901));
   MUX4EHD U6351 (.S1(n6038), 
	.S0(n7444), 
	.O(n4903), 
	.D(n4887), 
	.C(n4897), 
	.B(n4892), 
	.A(n4902));
   MUX4EHD U6352 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4904), 
	.D(\ram[63][2] ), 
	.C(\ram[61][2] ), 
	.B(\ram[62][2] ), 
	.A(\ram[60][2] ));
   MUX4EHD U6353 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4905), 
	.D(\ram[59][2] ), 
	.C(\ram[57][2] ), 
	.B(\ram[58][2] ), 
	.A(\ram[56][2] ));
   MUX4EHD U6354 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4906), 
	.D(\ram[55][2] ), 
	.C(\ram[53][2] ), 
	.B(\ram[54][2] ), 
	.A(\ram[52][2] ));
   MUX4EHD U6355 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4907), 
	.D(\ram[51][2] ), 
	.C(\ram[49][2] ), 
	.B(\ram[50][2] ), 
	.A(\ram[48][2] ));
   MUX4EHD U6356 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4908), 
	.D(n4904), 
	.C(n4906), 
	.B(n4905), 
	.A(n4907));
   MUX4EHD U6357 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4909), 
	.D(\ram[47][2] ), 
	.C(\ram[45][2] ), 
	.B(\ram[46][2] ), 
	.A(\ram[44][2] ));
   MUX4EHD U6358 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4910), 
	.D(\ram[43][2] ), 
	.C(\ram[41][2] ), 
	.B(\ram[42][2] ), 
	.A(\ram[40][2] ));
   MUX4EHD U6359 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4911), 
	.D(\ram[39][2] ), 
	.C(\ram[37][2] ), 
	.B(\ram[38][2] ), 
	.A(\ram[36][2] ));
   MUX4EHD U6360 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4912), 
	.D(\ram[35][2] ), 
	.C(\ram[33][2] ), 
	.B(\ram[34][2] ), 
	.A(\ram[32][2] ));
   MUX4EHD U6361 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4913), 
	.D(n4909), 
	.C(n4911), 
	.B(n4910), 
	.A(n4912));
   MUX4EHD U6362 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4914), 
	.D(\ram[31][2] ), 
	.C(\ram[29][2] ), 
	.B(\ram[30][2] ), 
	.A(\ram[28][2] ));
   MUX4EHD U6363 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4915), 
	.D(\ram[27][2] ), 
	.C(\ram[25][2] ), 
	.B(\ram[26][2] ), 
	.A(\ram[24][2] ));
   MUX4EHD U6364 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4916), 
	.D(\ram[23][2] ), 
	.C(\ram[21][2] ), 
	.B(\ram[22][2] ), 
	.A(\ram[20][2] ));
   MUX4EHD U6365 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4917), 
	.D(\ram[19][2] ), 
	.C(\ram[17][2] ), 
	.B(\ram[18][2] ), 
	.A(\ram[16][2] ));
   MUX4EHD U6366 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4918), 
	.D(n4914), 
	.C(n4916), 
	.B(n4915), 
	.A(n4917));
   MUX4EHD U6367 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4919), 
	.D(\ram[15][2] ), 
	.C(\ram[13][2] ), 
	.B(\ram[14][2] ), 
	.A(\ram[12][2] ));
   MUX4EHD U6368 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4920), 
	.D(\ram[11][2] ), 
	.C(\ram[9][2] ), 
	.B(\ram[10][2] ), 
	.A(\ram[8][2] ));
   MUX4EHD U6369 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4921), 
	.D(\ram[7][2] ), 
	.C(\ram[5][2] ), 
	.B(\ram[6][2] ), 
	.A(\ram[4][2] ));
   MUX4EHD U6370 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4922), 
	.D(\ram[3][2] ), 
	.C(\ram[1][2] ), 
	.B(\ram[2][2] ), 
	.A(\ram[0][2] ));
   MUX4EHD U6371 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4923), 
	.D(n4919), 
	.C(n4921), 
	.B(n4920), 
	.A(n4922));
   MUX4EHD U6372 (.S1(n6038), 
	.S0(n7444), 
	.O(n4924), 
	.D(n4908), 
	.C(n4918), 
	.B(n4913), 
	.A(n4923));
   MUX4EHD U6373 (.S1(n6469), 
	.S0(n6470), 
	.O(N4139), 
	.D(n4861), 
	.C(n4903), 
	.B(n4882), 
	.A(n4924));
   MUX4EHD U6374 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4925), 
	.D(\ram[255][3] ), 
	.C(\ram[253][3] ), 
	.B(\ram[254][3] ), 
	.A(\ram[252][3] ));
   MUX4EHD U6375 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4926), 
	.D(\ram[251][3] ), 
	.C(\ram[249][3] ), 
	.B(\ram[250][3] ), 
	.A(\ram[248][3] ));
   MUX4EHD U6376 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4927), 
	.D(\ram[247][3] ), 
	.C(\ram[245][3] ), 
	.B(\ram[246][3] ), 
	.A(\ram[244][3] ));
   MUX4EHD U6377 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4928), 
	.D(\ram[243][3] ), 
	.C(\ram[241][3] ), 
	.B(\ram[242][3] ), 
	.A(\ram[240][3] ));
   MUX4EHD U6378 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4929), 
	.D(n4925), 
	.C(n4927), 
	.B(n4926), 
	.A(n4928));
   MUX4EHD U6379 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4930), 
	.D(\ram[239][3] ), 
	.C(\ram[237][3] ), 
	.B(\ram[238][3] ), 
	.A(\ram[236][3] ));
   MUX4EHD U6380 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4931), 
	.D(\ram[235][3] ), 
	.C(\ram[233][3] ), 
	.B(\ram[234][3] ), 
	.A(\ram[232][3] ));
   MUX4EHD U6381 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4932), 
	.D(\ram[231][3] ), 
	.C(\ram[229][3] ), 
	.B(\ram[230][3] ), 
	.A(\ram[228][3] ));
   MUX4EHD U6382 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4933), 
	.D(\ram[227][3] ), 
	.C(\ram[225][3] ), 
	.B(\ram[226][3] ), 
	.A(\ram[224][3] ));
   MUX4EHD U6383 (.S1(n6136), 
	.S0(n7442), 
	.O(n4934), 
	.D(n4930), 
	.C(n4932), 
	.B(n4931), 
	.A(n4933));
   MUX4EHD U6384 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4935), 
	.D(\ram[223][3] ), 
	.C(\ram[221][3] ), 
	.B(\ram[222][3] ), 
	.A(\ram[220][3] ));
   MUX4EHD U6385 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4936), 
	.D(\ram[219][3] ), 
	.C(\ram[217][3] ), 
	.B(\ram[218][3] ), 
	.A(\ram[216][3] ));
   MUX4EHD U6386 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4937), 
	.D(\ram[215][3] ), 
	.C(\ram[213][3] ), 
	.B(\ram[214][3] ), 
	.A(\ram[212][3] ));
   MUX4EHD U6387 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4938), 
	.D(\ram[211][3] ), 
	.C(\ram[209][3] ), 
	.B(\ram[210][3] ), 
	.A(\ram[208][3] ));
   MUX4EHD U6388 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4939), 
	.D(n4935), 
	.C(n4937), 
	.B(n4936), 
	.A(n4938));
   MUX4EHD U6389 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4940), 
	.D(\ram[207][3] ), 
	.C(\ram[205][3] ), 
	.B(\ram[206][3] ), 
	.A(\ram[204][3] ));
   MUX4EHD U6390 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4941), 
	.D(\ram[203][3] ), 
	.C(\ram[201][3] ), 
	.B(\ram[202][3] ), 
	.A(\ram[200][3] ));
   MUX4EHD U6391 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4942), 
	.D(\ram[199][3] ), 
	.C(\ram[197][3] ), 
	.B(\ram[198][3] ), 
	.A(\ram[196][3] ));
   MUX4EHD U6392 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4943), 
	.D(\ram[195][3] ), 
	.C(\ram[193][3] ), 
	.B(\ram[194][3] ), 
	.A(\ram[192][3] ));
   MUX4EHD U6393 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4944), 
	.D(n4940), 
	.C(n4942), 
	.B(n4941), 
	.A(n4943));
   MUX4EHD U6394 (.S1(n6038), 
	.S0(n7444), 
	.O(n4945), 
	.D(n4929), 
	.C(n4939), 
	.B(n4934), 
	.A(n4944));
   MUX4EHD U6395 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4946), 
	.D(\ram[191][3] ), 
	.C(\ram[189][3] ), 
	.B(\ram[190][3] ), 
	.A(\ram[188][3] ));
   MUX4EHD U6396 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4947), 
	.D(\ram[187][3] ), 
	.C(\ram[185][3] ), 
	.B(\ram[186][3] ), 
	.A(\ram[184][3] ));
   MUX4EHD U6397 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4948), 
	.D(\ram[183][3] ), 
	.C(\ram[181][3] ), 
	.B(\ram[182][3] ), 
	.A(\ram[180][3] ));
   MUX4EHD U6398 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4949), 
	.D(\ram[179][3] ), 
	.C(\ram[177][3] ), 
	.B(\ram[178][3] ), 
	.A(\ram[176][3] ));
   MUX4EHD U6399 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4950), 
	.D(n4946), 
	.C(n4948), 
	.B(n4947), 
	.A(n4949));
   MUX4EHD U6400 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4951), 
	.D(\ram[175][3] ), 
	.C(\ram[173][3] ), 
	.B(\ram[174][3] ), 
	.A(\ram[172][3] ));
   MUX4EHD U6401 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4952), 
	.D(\ram[171][3] ), 
	.C(\ram[169][3] ), 
	.B(\ram[170][3] ), 
	.A(\ram[168][3] ));
   MUX4EHD U6402 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4953), 
	.D(\ram[167][3] ), 
	.C(\ram[165][3] ), 
	.B(\ram[166][3] ), 
	.A(\ram[164][3] ));
   MUX4EHD U6403 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4954), 
	.D(\ram[163][3] ), 
	.C(\ram[161][3] ), 
	.B(\ram[162][3] ), 
	.A(\ram[160][3] ));
   MUX4EHD U6404 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4955), 
	.D(n4951), 
	.C(n4953), 
	.B(n4952), 
	.A(n4954));
   MUX4EHD U6405 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4956), 
	.D(\ram[159][3] ), 
	.C(\ram[157][3] ), 
	.B(\ram[158][3] ), 
	.A(\ram[156][3] ));
   MUX4EHD U6406 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4957), 
	.D(\ram[155][3] ), 
	.C(\ram[153][3] ), 
	.B(\ram[154][3] ), 
	.A(\ram[152][3] ));
   MUX4EHD U6407 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4958), 
	.D(\ram[151][3] ), 
	.C(\ram[149][3] ), 
	.B(\ram[150][3] ), 
	.A(\ram[148][3] ));
   MUX4EHD U6408 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4959), 
	.D(\ram[147][3] ), 
	.C(\ram[145][3] ), 
	.B(\ram[146][3] ), 
	.A(\ram[144][3] ));
   MUX4EHD U6409 (.S1(n6136), 
	.S0(n7442), 
	.O(n4960), 
	.D(n4956), 
	.C(n4958), 
	.B(n4957), 
	.A(n4959));
   MUX4EHD U6410 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4961), 
	.D(\ram[143][3] ), 
	.C(\ram[141][3] ), 
	.B(\ram[142][3] ), 
	.A(\ram[140][3] ));
   MUX4EHD U6411 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4962), 
	.D(\ram[139][3] ), 
	.C(\ram[137][3] ), 
	.B(\ram[138][3] ), 
	.A(\ram[136][3] ));
   MUX4EHD U6412 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4963), 
	.D(\ram[135][3] ), 
	.C(\ram[133][3] ), 
	.B(\ram[134][3] ), 
	.A(\ram[132][3] ));
   MUX4EHD U6413 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4964), 
	.D(\ram[131][3] ), 
	.C(\ram[129][3] ), 
	.B(\ram[130][3] ), 
	.A(\ram[128][3] ));
   MUX4EHD U6414 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4965), 
	.D(n4961), 
	.C(n4963), 
	.B(n4962), 
	.A(n4964));
   MUX4EHD U6415 (.S1(n6038), 
	.S0(n7444), 
	.O(n4966), 
	.D(n4950), 
	.C(n4960), 
	.B(n4955), 
	.A(n4965));
   MUX4EHD U6416 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4967), 
	.D(\ram[127][3] ), 
	.C(\ram[125][3] ), 
	.B(\ram[126][3] ), 
	.A(\ram[124][3] ));
   MUX4EHD U6417 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4968), 
	.D(\ram[123][3] ), 
	.C(\ram[121][3] ), 
	.B(\ram[122][3] ), 
	.A(\ram[120][3] ));
   MUX4EHD U6418 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4969), 
	.D(\ram[119][3] ), 
	.C(\ram[117][3] ), 
	.B(\ram[118][3] ), 
	.A(\ram[116][3] ));
   MUX4EHD U6419 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4970), 
	.D(\ram[115][3] ), 
	.C(\ram[113][3] ), 
	.B(\ram[114][3] ), 
	.A(\ram[112][3] ));
   MUX4EHD U6420 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4971), 
	.D(n4967), 
	.C(n4969), 
	.B(n4968), 
	.A(n4970));
   MUX4EHD U6421 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4972), 
	.D(\ram[111][3] ), 
	.C(\ram[109][3] ), 
	.B(\ram[110][3] ), 
	.A(\ram[108][3] ));
   MUX4EHD U6422 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4973), 
	.D(\ram[107][3] ), 
	.C(\ram[105][3] ), 
	.B(\ram[106][3] ), 
	.A(\ram[104][3] ));
   MUX4EHD U6423 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4974), 
	.D(\ram[103][3] ), 
	.C(\ram[101][3] ), 
	.B(\ram[102][3] ), 
	.A(\ram[100][3] ));
   MUX4EHD U6424 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4975), 
	.D(\ram[99][3] ), 
	.C(\ram[97][3] ), 
	.B(\ram[98][3] ), 
	.A(\ram[96][3] ));
   MUX4EHD U6425 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4976), 
	.D(n4972), 
	.C(n4974), 
	.B(n4973), 
	.A(n4975));
   MUX4EHD U6426 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4977), 
	.D(\ram[95][3] ), 
	.C(\ram[93][3] ), 
	.B(\ram[94][3] ), 
	.A(\ram[92][3] ));
   MUX4EHD U6427 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4978), 
	.D(\ram[91][3] ), 
	.C(\ram[89][3] ), 
	.B(\ram[90][3] ), 
	.A(\ram[88][3] ));
   MUX4EHD U6428 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4979), 
	.D(\ram[87][3] ), 
	.C(\ram[85][3] ), 
	.B(\ram[86][3] ), 
	.A(\ram[84][3] ));
   MUX4EHD U6429 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4980), 
	.D(\ram[83][3] ), 
	.C(\ram[81][3] ), 
	.B(\ram[82][3] ), 
	.A(\ram[80][3] ));
   MUX4EHD U6430 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4981), 
	.D(n4977), 
	.C(n4979), 
	.B(n4978), 
	.A(n4980));
   MUX4EHD U6431 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4982), 
	.D(\ram[79][3] ), 
	.C(\ram[77][3] ), 
	.B(\ram[78][3] ), 
	.A(\ram[76][3] ));
   MUX4EHD U6432 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4983), 
	.D(\ram[75][3] ), 
	.C(\ram[73][3] ), 
	.B(\ram[74][3] ), 
	.A(\ram[72][3] ));
   MUX4EHD U6433 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4984), 
	.D(\ram[71][3] ), 
	.C(\ram[69][3] ), 
	.B(\ram[70][3] ), 
	.A(\ram[68][3] ));
   MUX4EHD U6434 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4985), 
	.D(\ram[67][3] ), 
	.C(\ram[65][3] ), 
	.B(\ram[66][3] ), 
	.A(\ram[64][3] ));
   MUX4EHD U6435 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4986), 
	.D(n4982), 
	.C(n4984), 
	.B(n4983), 
	.A(n4985));
   MUX4EHD U6436 (.S1(n6038), 
	.S0(n7444), 
	.O(n4987), 
	.D(n4971), 
	.C(n4981), 
	.B(n4976), 
	.A(n4986));
   MUX4EHD U6437 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4988), 
	.D(\ram[63][3] ), 
	.C(\ram[61][3] ), 
	.B(\ram[62][3] ), 
	.A(\ram[60][3] ));
   MUX4EHD U6438 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4989), 
	.D(\ram[59][3] ), 
	.C(\ram[57][3] ), 
	.B(\ram[58][3] ), 
	.A(\ram[56][3] ));
   MUX4EHD U6439 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4990), 
	.D(\ram[55][3] ), 
	.C(\ram[53][3] ), 
	.B(\ram[54][3] ), 
	.A(\ram[52][3] ));
   MUX4EHD U6440 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4991), 
	.D(\ram[51][3] ), 
	.C(\ram[49][3] ), 
	.B(\ram[50][3] ), 
	.A(\ram[48][3] ));
   MUX4EHD U6441 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4992), 
	.D(n4988), 
	.C(n4990), 
	.B(n4989), 
	.A(n4991));
   MUX4EHD U6442 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4993), 
	.D(\ram[47][3] ), 
	.C(\ram[45][3] ), 
	.B(\ram[46][3] ), 
	.A(\ram[44][3] ));
   MUX4EHD U6443 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4994), 
	.D(\ram[43][3] ), 
	.C(\ram[41][3] ), 
	.B(\ram[42][3] ), 
	.A(\ram[40][3] ));
   MUX4EHD U6444 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4995), 
	.D(\ram[39][3] ), 
	.C(\ram[37][3] ), 
	.B(\ram[38][3] ), 
	.A(\ram[36][3] ));
   MUX4EHD U6445 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4996), 
	.D(\ram[35][3] ), 
	.C(\ram[33][3] ), 
	.B(\ram[34][3] ), 
	.A(\ram[32][3] ));
   MUX4EHD U6446 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4997), 
	.D(n4993), 
	.C(n4995), 
	.B(n4994), 
	.A(n4996));
   MUX4EHD U6447 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4998), 
	.D(\ram[31][3] ), 
	.C(\ram[29][3] ), 
	.B(\ram[30][3] ), 
	.A(\ram[28][3] ));
   MUX4EHD U6448 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4999), 
	.D(\ram[27][3] ), 
	.C(\ram[25][3] ), 
	.B(\ram[26][3] ), 
	.A(\ram[24][3] ));
   MUX4EHD U6449 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5000), 
	.D(\ram[23][3] ), 
	.C(\ram[21][3] ), 
	.B(\ram[22][3] ), 
	.A(\ram[20][3] ));
   MUX4EHD U6450 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5001), 
	.D(\ram[19][3] ), 
	.C(\ram[17][3] ), 
	.B(\ram[18][3] ), 
	.A(\ram[16][3] ));
   MUX4EHD U6451 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5002), 
	.D(n4998), 
	.C(n5000), 
	.B(n4999), 
	.A(n5001));
   MUX4EHD U6452 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5003), 
	.D(\ram[15][3] ), 
	.C(\ram[13][3] ), 
	.B(\ram[14][3] ), 
	.A(\ram[12][3] ));
   MUX4EHD U6453 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5004), 
	.D(\ram[11][3] ), 
	.C(\ram[9][3] ), 
	.B(\ram[10][3] ), 
	.A(\ram[8][3] ));
   MUX4EHD U6454 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5005), 
	.D(\ram[7][3] ), 
	.C(\ram[5][3] ), 
	.B(\ram[6][3] ), 
	.A(\ram[4][3] ));
   MUX4EHD U6455 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5006), 
	.D(\ram[3][3] ), 
	.C(\ram[1][3] ), 
	.B(\ram[2][3] ), 
	.A(\ram[0][3] ));
   MUX4EHD U6456 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5007), 
	.D(n5003), 
	.C(n5005), 
	.B(n5004), 
	.A(n5006));
   MUX4EHD U6457 (.S1(n6038), 
	.S0(n7444), 
	.O(n5008), 
	.D(n4992), 
	.C(n5002), 
	.B(n4997), 
	.A(n5007));
   MUX4EHD U6458 (.S1(n6469), 
	.S0(n6470), 
	.O(N4138), 
	.D(n4945), 
	.C(n4987), 
	.B(n4966), 
	.A(n5008));
   MUX4EHD U6459 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5009), 
	.D(\ram[255][4] ), 
	.C(\ram[253][4] ), 
	.B(\ram[254][4] ), 
	.A(\ram[252][4] ));
   MUX4EHD U6460 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5010), 
	.D(\ram[251][4] ), 
	.C(\ram[249][4] ), 
	.B(\ram[250][4] ), 
	.A(\ram[248][4] ));
   MUX4EHD U6461 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5011), 
	.D(\ram[247][4] ), 
	.C(\ram[245][4] ), 
	.B(\ram[246][4] ), 
	.A(\ram[244][4] ));
   MUX4EHD U6462 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5012), 
	.D(\ram[243][4] ), 
	.C(\ram[241][4] ), 
	.B(\ram[242][4] ), 
	.A(\ram[240][4] ));
   MUX4EHD U6463 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5013), 
	.D(n5009), 
	.C(n5011), 
	.B(n5010), 
	.A(n5012));
   MUX4EHD U6464 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5014), 
	.D(\ram[239][4] ), 
	.C(\ram[237][4] ), 
	.B(\ram[238][4] ), 
	.A(\ram[236][4] ));
   MUX4EHD U6465 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5015), 
	.D(\ram[235][4] ), 
	.C(\ram[233][4] ), 
	.B(\ram[234][4] ), 
	.A(\ram[232][4] ));
   MUX4EHD U6466 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5016), 
	.D(\ram[231][4] ), 
	.C(\ram[229][4] ), 
	.B(\ram[230][4] ), 
	.A(\ram[228][4] ));
   MUX4EHD U6467 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5017), 
	.D(\ram[227][4] ), 
	.C(\ram[225][4] ), 
	.B(\ram[226][4] ), 
	.A(\ram[224][4] ));
   MUX4EHD U6468 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5018), 
	.D(n5014), 
	.C(n5016), 
	.B(n5015), 
	.A(n5017));
   MUX4EHD U6469 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5019), 
	.D(\ram[223][4] ), 
	.C(\ram[221][4] ), 
	.B(\ram[222][4] ), 
	.A(\ram[220][4] ));
   MUX4EHD U6470 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5020), 
	.D(\ram[219][4] ), 
	.C(\ram[217][4] ), 
	.B(\ram[218][4] ), 
	.A(\ram[216][4] ));
   MUX4EHD U6471 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5021), 
	.D(\ram[215][4] ), 
	.C(\ram[213][4] ), 
	.B(\ram[214][4] ), 
	.A(\ram[212][4] ));
   MUX4EHD U6472 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5022), 
	.D(\ram[211][4] ), 
	.C(\ram[209][4] ), 
	.B(\ram[210][4] ), 
	.A(\ram[208][4] ));
   MUX4EHD U6473 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5023), 
	.D(n5019), 
	.C(n5021), 
	.B(n5020), 
	.A(n5022));
   MUX4EHD U6474 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5024), 
	.D(\ram[207][4] ), 
	.C(\ram[205][4] ), 
	.B(\ram[206][4] ), 
	.A(\ram[204][4] ));
   MUX4EHD U6475 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5025), 
	.D(\ram[203][4] ), 
	.C(\ram[201][4] ), 
	.B(\ram[202][4] ), 
	.A(\ram[200][4] ));
   MUX4EHD U6476 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5026), 
	.D(\ram[199][4] ), 
	.C(\ram[197][4] ), 
	.B(\ram[198][4] ), 
	.A(\ram[196][4] ));
   MUX4EHD U6477 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5027), 
	.D(\ram[195][4] ), 
	.C(\ram[193][4] ), 
	.B(\ram[194][4] ), 
	.A(\ram[192][4] ));
   MUX4EHD U6478 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5028), 
	.D(n5024), 
	.C(n5026), 
	.B(n5025), 
	.A(n5027));
   MUX4EHD U6479 (.S1(n6038), 
	.S0(n7444), 
	.O(n5029), 
	.D(n5013), 
	.C(n5023), 
	.B(n5018), 
	.A(n5028));
   MUX4EHD U6480 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5030), 
	.D(\ram[191][4] ), 
	.C(\ram[189][4] ), 
	.B(\ram[190][4] ), 
	.A(\ram[188][4] ));
   MUX4EHD U6481 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5031), 
	.D(\ram[187][4] ), 
	.C(\ram[185][4] ), 
	.B(\ram[186][4] ), 
	.A(\ram[184][4] ));
   MUX4EHD U6482 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5032), 
	.D(\ram[183][4] ), 
	.C(\ram[181][4] ), 
	.B(\ram[182][4] ), 
	.A(\ram[180][4] ));
   MUX4EHD U6483 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5033), 
	.D(\ram[179][4] ), 
	.C(\ram[177][4] ), 
	.B(\ram[178][4] ), 
	.A(\ram[176][4] ));
   MUX4EHD U6484 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5034), 
	.D(n5030), 
	.C(n5032), 
	.B(n5031), 
	.A(n5033));
   MUX4EHD U6485 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5035), 
	.D(\ram[175][4] ), 
	.C(\ram[173][4] ), 
	.B(\ram[174][4] ), 
	.A(\ram[172][4] ));
   MUX4EHD U6486 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5036), 
	.D(\ram[171][4] ), 
	.C(\ram[169][4] ), 
	.B(\ram[170][4] ), 
	.A(\ram[168][4] ));
   MUX4EHD U6487 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5037), 
	.D(\ram[167][4] ), 
	.C(\ram[165][4] ), 
	.B(\ram[166][4] ), 
	.A(\ram[164][4] ));
   MUX4EHD U6488 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5038), 
	.D(\ram[163][4] ), 
	.C(\ram[161][4] ), 
	.B(\ram[162][4] ), 
	.A(\ram[160][4] ));
   MUX4EHD U6489 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5039), 
	.D(n5035), 
	.C(n5037), 
	.B(n5036), 
	.A(n5038));
   MUX4EHD U6490 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5040), 
	.D(\ram[159][4] ), 
	.C(\ram[157][4] ), 
	.B(\ram[158][4] ), 
	.A(\ram[156][4] ));
   MUX4EHD U6491 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5041), 
	.D(\ram[155][4] ), 
	.C(\ram[153][4] ), 
	.B(\ram[154][4] ), 
	.A(\ram[152][4] ));
   MUX4EHD U6492 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5042), 
	.D(\ram[151][4] ), 
	.C(\ram[149][4] ), 
	.B(\ram[150][4] ), 
	.A(\ram[148][4] ));
   MUX4EHD U6493 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5043), 
	.D(\ram[147][4] ), 
	.C(\ram[145][4] ), 
	.B(\ram[146][4] ), 
	.A(\ram[144][4] ));
   MUX4EHD U6494 (.S1(n6136), 
	.S0(n7442), 
	.O(n5044), 
	.D(n5040), 
	.C(n5042), 
	.B(n5041), 
	.A(n5043));
   MUX4EHD U6495 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5045), 
	.D(\ram[143][4] ), 
	.C(\ram[141][4] ), 
	.B(\ram[142][4] ), 
	.A(\ram[140][4] ));
   MUX4EHD U6496 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5046), 
	.D(\ram[139][4] ), 
	.C(\ram[137][4] ), 
	.B(\ram[138][4] ), 
	.A(\ram[136][4] ));
   MUX4EHD U6497 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5047), 
	.D(\ram[135][4] ), 
	.C(\ram[133][4] ), 
	.B(\ram[134][4] ), 
	.A(\ram[132][4] ));
   MUX4EHD U6498 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5048), 
	.D(\ram[131][4] ), 
	.C(\ram[129][4] ), 
	.B(\ram[130][4] ), 
	.A(\ram[128][4] ));
   MUX4EHD U6499 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5049), 
	.D(n5045), 
	.C(n5047), 
	.B(n5046), 
	.A(n5048));
   MUX4EHD U6500 (.S1(n6038), 
	.S0(n7444), 
	.O(n5050), 
	.D(n5034), 
	.C(n5044), 
	.B(n5039), 
	.A(n5049));
   MUX4EHD U6501 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5051), 
	.D(\ram[127][4] ), 
	.C(\ram[125][4] ), 
	.B(\ram[126][4] ), 
	.A(\ram[124][4] ));
   MUX4EHD U6502 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5052), 
	.D(\ram[123][4] ), 
	.C(\ram[121][4] ), 
	.B(\ram[122][4] ), 
	.A(\ram[120][4] ));
   MUX4EHD U6503 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5053), 
	.D(\ram[119][4] ), 
	.C(\ram[117][4] ), 
	.B(\ram[118][4] ), 
	.A(\ram[116][4] ));
   MUX4EHD U6504 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5054), 
	.D(\ram[115][4] ), 
	.C(\ram[113][4] ), 
	.B(\ram[114][4] ), 
	.A(\ram[112][4] ));
   MUX4EHD U6505 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5055), 
	.D(n5051), 
	.C(n5053), 
	.B(n5052), 
	.A(n5054));
   MUX4EHD U6506 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5056), 
	.D(\ram[111][4] ), 
	.C(\ram[109][4] ), 
	.B(\ram[110][4] ), 
	.A(\ram[108][4] ));
   MUX4EHD U6507 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5057), 
	.D(\ram[107][4] ), 
	.C(\ram[105][4] ), 
	.B(\ram[106][4] ), 
	.A(\ram[104][4] ));
   MUX4EHD U6508 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5058), 
	.D(\ram[103][4] ), 
	.C(\ram[101][4] ), 
	.B(\ram[102][4] ), 
	.A(\ram[100][4] ));
   MUX4EHD U6509 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5059), 
	.D(\ram[99][4] ), 
	.C(\ram[97][4] ), 
	.B(\ram[98][4] ), 
	.A(\ram[96][4] ));
   MUX4EHD U6510 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5060), 
	.D(n5056), 
	.C(n5058), 
	.B(n5057), 
	.A(n5059));
   MUX4EHD U6511 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5061), 
	.D(\ram[95][4] ), 
	.C(\ram[93][4] ), 
	.B(\ram[94][4] ), 
	.A(\ram[92][4] ));
   MUX4EHD U6512 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5062), 
	.D(\ram[91][4] ), 
	.C(\ram[89][4] ), 
	.B(\ram[90][4] ), 
	.A(\ram[88][4] ));
   MUX4EHD U6513 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5063), 
	.D(\ram[87][4] ), 
	.C(\ram[85][4] ), 
	.B(\ram[86][4] ), 
	.A(\ram[84][4] ));
   MUX4EHD U6514 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5064), 
	.D(\ram[83][4] ), 
	.C(\ram[81][4] ), 
	.B(\ram[82][4] ), 
	.A(\ram[80][4] ));
   MUX4EHD U6515 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5065), 
	.D(n5061), 
	.C(n5063), 
	.B(n5062), 
	.A(n5064));
   MUX4EHD U6516 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5066), 
	.D(\ram[79][4] ), 
	.C(\ram[77][4] ), 
	.B(\ram[78][4] ), 
	.A(\ram[76][4] ));
   MUX4EHD U6517 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5067), 
	.D(\ram[75][4] ), 
	.C(\ram[73][4] ), 
	.B(\ram[74][4] ), 
	.A(\ram[72][4] ));
   MUX4EHD U6518 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5068), 
	.D(\ram[71][4] ), 
	.C(\ram[69][4] ), 
	.B(\ram[70][4] ), 
	.A(\ram[68][4] ));
   MUX4EHD U6519 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5069), 
	.D(\ram[67][4] ), 
	.C(\ram[65][4] ), 
	.B(\ram[66][4] ), 
	.A(\ram[64][4] ));
   MUX4EHD U6520 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5070), 
	.D(n5066), 
	.C(n5068), 
	.B(n5067), 
	.A(n5069));
   MUX4EHD U6521 (.S1(n6038), 
	.S0(n7444), 
	.O(n5071), 
	.D(n5055), 
	.C(n5065), 
	.B(n5060), 
	.A(n5070));
   MUX4EHD U6522 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5072), 
	.D(\ram[63][4] ), 
	.C(\ram[61][4] ), 
	.B(\ram[62][4] ), 
	.A(\ram[60][4] ));
   MUX4EHD U6523 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5073), 
	.D(\ram[59][4] ), 
	.C(\ram[57][4] ), 
	.B(\ram[58][4] ), 
	.A(\ram[56][4] ));
   MUX4EHD U6524 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5074), 
	.D(\ram[55][4] ), 
	.C(\ram[53][4] ), 
	.B(\ram[54][4] ), 
	.A(\ram[52][4] ));
   MUX4EHD U6525 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5075), 
	.D(\ram[51][4] ), 
	.C(\ram[49][4] ), 
	.B(\ram[50][4] ), 
	.A(\ram[48][4] ));
   MUX4EHD U6526 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5076), 
	.D(n5072), 
	.C(n5074), 
	.B(n5073), 
	.A(n5075));
   MUX4EHD U6527 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5077), 
	.D(\ram[47][4] ), 
	.C(\ram[45][4] ), 
	.B(\ram[46][4] ), 
	.A(\ram[44][4] ));
   MUX4EHD U6528 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5078), 
	.D(\ram[43][4] ), 
	.C(\ram[41][4] ), 
	.B(\ram[42][4] ), 
	.A(\ram[40][4] ));
   MUX4EHD U6529 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5079), 
	.D(\ram[39][4] ), 
	.C(\ram[37][4] ), 
	.B(\ram[38][4] ), 
	.A(\ram[36][4] ));
   MUX4EHD U6530 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5080), 
	.D(\ram[35][4] ), 
	.C(\ram[33][4] ), 
	.B(\ram[34][4] ), 
	.A(\ram[32][4] ));
   MUX4EHD U6531 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5081), 
	.D(n5077), 
	.C(n5079), 
	.B(n5078), 
	.A(n5080));
   MUX4EHD U6532 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5082), 
	.D(\ram[31][4] ), 
	.C(\ram[29][4] ), 
	.B(\ram[30][4] ), 
	.A(\ram[28][4] ));
   MUX4EHD U6533 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5083), 
	.D(\ram[27][4] ), 
	.C(\ram[25][4] ), 
	.B(\ram[26][4] ), 
	.A(\ram[24][4] ));
   MUX4EHD U6534 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5084), 
	.D(\ram[23][4] ), 
	.C(\ram[21][4] ), 
	.B(\ram[22][4] ), 
	.A(\ram[20][4] ));
   MUX4EHD U6535 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5085), 
	.D(\ram[19][4] ), 
	.C(\ram[17][4] ), 
	.B(\ram[18][4] ), 
	.A(\ram[16][4] ));
   MUX4EHD U6536 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5086), 
	.D(n5082), 
	.C(n5084), 
	.B(n5083), 
	.A(n5085));
   MUX4EHD U6537 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5087), 
	.D(\ram[15][4] ), 
	.C(\ram[13][4] ), 
	.B(\ram[14][4] ), 
	.A(\ram[12][4] ));
   MUX4EHD U6538 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5088), 
	.D(\ram[11][4] ), 
	.C(\ram[9][4] ), 
	.B(\ram[10][4] ), 
	.A(\ram[8][4] ));
   MUX4EHD U6539 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5089), 
	.D(\ram[7][4] ), 
	.C(\ram[5][4] ), 
	.B(\ram[6][4] ), 
	.A(\ram[4][4] ));
   MUX4EHD U6540 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5090), 
	.D(\ram[3][4] ), 
	.C(\ram[1][4] ), 
	.B(\ram[2][4] ), 
	.A(\ram[0][4] ));
   MUX4EHD U6541 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5091), 
	.D(n5087), 
	.C(n5089), 
	.B(n5088), 
	.A(n5090));
   MUX4EHD U6542 (.S1(n6038), 
	.S0(n7444), 
	.O(n5092), 
	.D(n5076), 
	.C(n5086), 
	.B(n5081), 
	.A(n5091));
   MUX4EHD U6543 (.S1(n6469), 
	.S0(n6470), 
	.O(N4137), 
	.D(n5029), 
	.C(n5071), 
	.B(n5050), 
	.A(n5092));
   MUX4EHD U6544 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5093), 
	.D(\ram[255][5] ), 
	.C(\ram[253][5] ), 
	.B(\ram[254][5] ), 
	.A(\ram[252][5] ));
   MUX4EHD U6545 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5094), 
	.D(\ram[251][5] ), 
	.C(\ram[249][5] ), 
	.B(\ram[250][5] ), 
	.A(\ram[248][5] ));
   MUX4EHD U6546 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5095), 
	.D(\ram[247][5] ), 
	.C(\ram[245][5] ), 
	.B(\ram[246][5] ), 
	.A(\ram[244][5] ));
   MUX4EHD U6547 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5096), 
	.D(\ram[243][5] ), 
	.C(\ram[241][5] ), 
	.B(\ram[242][5] ), 
	.A(\ram[240][5] ));
   MUX4EHD U6548 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5097), 
	.D(n5093), 
	.C(n5095), 
	.B(n5094), 
	.A(n5096));
   MUX4EHD U6549 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5098), 
	.D(\ram[239][5] ), 
	.C(\ram[237][5] ), 
	.B(\ram[238][5] ), 
	.A(\ram[236][5] ));
   MUX4EHD U6550 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5099), 
	.D(\ram[235][5] ), 
	.C(\ram[233][5] ), 
	.B(\ram[234][5] ), 
	.A(\ram[232][5] ));
   MUX4EHD U6551 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5100), 
	.D(\ram[231][5] ), 
	.C(\ram[229][5] ), 
	.B(\ram[230][5] ), 
	.A(\ram[228][5] ));
   MUX4EHD U6552 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5101), 
	.D(\ram[227][5] ), 
	.C(\ram[225][5] ), 
	.B(\ram[226][5] ), 
	.A(\ram[224][5] ));
   MUX4EHD U6553 (.S1(n6136), 
	.S0(n7442), 
	.O(n5102), 
	.D(n5098), 
	.C(n5100), 
	.B(n5099), 
	.A(n5101));
   MUX4EHD U6554 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5103), 
	.D(\ram[223][5] ), 
	.C(\ram[221][5] ), 
	.B(\ram[222][5] ), 
	.A(\ram[220][5] ));
   MUX4EHD U6555 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5104), 
	.D(\ram[219][5] ), 
	.C(\ram[217][5] ), 
	.B(\ram[218][5] ), 
	.A(\ram[216][5] ));
   MUX4EHD U6556 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5105), 
	.D(\ram[215][5] ), 
	.C(\ram[213][5] ), 
	.B(\ram[214][5] ), 
	.A(\ram[212][5] ));
   MUX4EHD U6557 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5106), 
	.D(\ram[211][5] ), 
	.C(\ram[209][5] ), 
	.B(\ram[210][5] ), 
	.A(\ram[208][5] ));
   MUX4EHD U6558 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5107), 
	.D(n5103), 
	.C(n5105), 
	.B(n5104), 
	.A(n5106));
   MUX4EHD U6559 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5108), 
	.D(\ram[207][5] ), 
	.C(\ram[205][5] ), 
	.B(\ram[206][5] ), 
	.A(\ram[204][5] ));
   MUX4EHD U6560 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5109), 
	.D(\ram[203][5] ), 
	.C(\ram[201][5] ), 
	.B(\ram[202][5] ), 
	.A(\ram[200][5] ));
   MUX4EHD U6561 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5110), 
	.D(\ram[199][5] ), 
	.C(\ram[197][5] ), 
	.B(\ram[198][5] ), 
	.A(\ram[196][5] ));
   MUX4EHD U6562 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5111), 
	.D(\ram[195][5] ), 
	.C(\ram[193][5] ), 
	.B(\ram[194][5] ), 
	.A(\ram[192][5] ));
   MUX4EHD U6563 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5112), 
	.D(n5108), 
	.C(n5110), 
	.B(n5109), 
	.A(n5111));
   MUX4EHD U6564 (.S1(n6038), 
	.S0(n7444), 
	.O(n5113), 
	.D(n5097), 
	.C(n5107), 
	.B(n5102), 
	.A(n5112));
   MUX4EHD U6565 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5114), 
	.D(\ram[191][5] ), 
	.C(\ram[189][5] ), 
	.B(\ram[190][5] ), 
	.A(\ram[188][5] ));
   MUX4EHD U6566 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5115), 
	.D(\ram[187][5] ), 
	.C(\ram[185][5] ), 
	.B(\ram[186][5] ), 
	.A(\ram[184][5] ));
   MUX4EHD U6567 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5116), 
	.D(\ram[183][5] ), 
	.C(\ram[181][5] ), 
	.B(\ram[182][5] ), 
	.A(\ram[180][5] ));
   MUX4EHD U6568 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5117), 
	.D(\ram[179][5] ), 
	.C(\ram[177][5] ), 
	.B(\ram[178][5] ), 
	.A(\ram[176][5] ));
   MUX4EHD U6569 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5118), 
	.D(n5114), 
	.C(n5116), 
	.B(n5115), 
	.A(n5117));
   MUX4EHD U6570 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5119), 
	.D(\ram[175][5] ), 
	.C(\ram[173][5] ), 
	.B(\ram[174][5] ), 
	.A(\ram[172][5] ));
   MUX4EHD U6571 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5120), 
	.D(\ram[171][5] ), 
	.C(\ram[169][5] ), 
	.B(\ram[170][5] ), 
	.A(\ram[168][5] ));
   MUX4EHD U6572 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5121), 
	.D(\ram[167][5] ), 
	.C(\ram[165][5] ), 
	.B(\ram[166][5] ), 
	.A(\ram[164][5] ));
   MUX4EHD U6573 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5122), 
	.D(\ram[163][5] ), 
	.C(\ram[161][5] ), 
	.B(\ram[162][5] ), 
	.A(\ram[160][5] ));
   MUX4EHD U6574 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5123), 
	.D(n5119), 
	.C(n5121), 
	.B(n5120), 
	.A(n5122));
   MUX4EHD U6575 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5124), 
	.D(\ram[159][5] ), 
	.C(\ram[157][5] ), 
	.B(\ram[158][5] ), 
	.A(\ram[156][5] ));
   MUX4EHD U6576 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5125), 
	.D(\ram[155][5] ), 
	.C(\ram[153][5] ), 
	.B(\ram[154][5] ), 
	.A(\ram[152][5] ));
   MUX4EHD U6577 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5126), 
	.D(\ram[151][5] ), 
	.C(\ram[149][5] ), 
	.B(\ram[150][5] ), 
	.A(\ram[148][5] ));
   MUX4EHD U6578 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5127), 
	.D(\ram[147][5] ), 
	.C(\ram[145][5] ), 
	.B(\ram[146][5] ), 
	.A(\ram[144][5] ));
   MUX4EHD U6579 (.S1(n6136), 
	.S0(n7442), 
	.O(n5128), 
	.D(n5124), 
	.C(n5126), 
	.B(n5125), 
	.A(n5127));
   MUX4EHD U6580 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5129), 
	.D(\ram[143][5] ), 
	.C(\ram[141][5] ), 
	.B(\ram[142][5] ), 
	.A(\ram[140][5] ));
   MUX4EHD U6581 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5130), 
	.D(\ram[139][5] ), 
	.C(\ram[137][5] ), 
	.B(\ram[138][5] ), 
	.A(\ram[136][5] ));
   MUX4EHD U6582 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5131), 
	.D(\ram[135][5] ), 
	.C(\ram[133][5] ), 
	.B(\ram[134][5] ), 
	.A(\ram[132][5] ));
   MUX4EHD U6583 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5132), 
	.D(\ram[131][5] ), 
	.C(\ram[129][5] ), 
	.B(\ram[130][5] ), 
	.A(\ram[128][5] ));
   MUX4EHD U6584 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5133), 
	.D(n5129), 
	.C(n5131), 
	.B(n5130), 
	.A(n5132));
   MUX4EHD U6585 (.S1(n6038), 
	.S0(n7444), 
	.O(n5134), 
	.D(n5118), 
	.C(n5128), 
	.B(n5123), 
	.A(n5133));
   MUX4EHD U6586 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5135), 
	.D(\ram[127][5] ), 
	.C(\ram[125][5] ), 
	.B(\ram[126][5] ), 
	.A(\ram[124][5] ));
   MUX4EHD U6587 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5136), 
	.D(\ram[123][5] ), 
	.C(\ram[121][5] ), 
	.B(\ram[122][5] ), 
	.A(\ram[120][5] ));
   MUX4EHD U6588 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5137), 
	.D(\ram[119][5] ), 
	.C(\ram[117][5] ), 
	.B(\ram[118][5] ), 
	.A(\ram[116][5] ));
   MUX4EHD U6589 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5138), 
	.D(\ram[115][5] ), 
	.C(\ram[113][5] ), 
	.B(\ram[114][5] ), 
	.A(\ram[112][5] ));
   MUX4EHD U6590 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5139), 
	.D(n5135), 
	.C(n5137), 
	.B(n5136), 
	.A(n5138));
   MUX4EHD U6591 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5140), 
	.D(\ram[111][5] ), 
	.C(\ram[109][5] ), 
	.B(\ram[110][5] ), 
	.A(\ram[108][5] ));
   MUX4EHD U6592 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5141), 
	.D(\ram[107][5] ), 
	.C(\ram[105][5] ), 
	.B(\ram[106][5] ), 
	.A(\ram[104][5] ));
   MUX4EHD U6593 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5142), 
	.D(\ram[103][5] ), 
	.C(\ram[101][5] ), 
	.B(\ram[102][5] ), 
	.A(\ram[100][5] ));
   MUX4EHD U6594 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5143), 
	.D(\ram[99][5] ), 
	.C(\ram[97][5] ), 
	.B(\ram[98][5] ), 
	.A(\ram[96][5] ));
   MUX4EHD U6595 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5144), 
	.D(n5140), 
	.C(n5142), 
	.B(n5141), 
	.A(n5143));
   MUX4EHD U6596 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5145), 
	.D(\ram[95][5] ), 
	.C(\ram[93][5] ), 
	.B(\ram[94][5] ), 
	.A(\ram[92][5] ));
   MUX4EHD U6597 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5146), 
	.D(\ram[91][5] ), 
	.C(\ram[89][5] ), 
	.B(\ram[90][5] ), 
	.A(\ram[88][5] ));
   MUX4EHD U6598 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5147), 
	.D(\ram[87][5] ), 
	.C(\ram[85][5] ), 
	.B(\ram[86][5] ), 
	.A(\ram[84][5] ));
   MUX4EHD U6599 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5148), 
	.D(\ram[83][5] ), 
	.C(\ram[81][5] ), 
	.B(\ram[82][5] ), 
	.A(\ram[80][5] ));
   MUX4EHD U6600 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5149), 
	.D(n5145), 
	.C(n5147), 
	.B(n5146), 
	.A(n5148));
   MUX4EHD U6601 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5150), 
	.D(\ram[79][5] ), 
	.C(\ram[77][5] ), 
	.B(\ram[78][5] ), 
	.A(\ram[76][5] ));
   MUX4EHD U6602 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5151), 
	.D(\ram[75][5] ), 
	.C(\ram[73][5] ), 
	.B(\ram[74][5] ), 
	.A(\ram[72][5] ));
   MUX4EHD U6603 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5152), 
	.D(\ram[71][5] ), 
	.C(\ram[69][5] ), 
	.B(\ram[70][5] ), 
	.A(\ram[68][5] ));
   MUX4EHD U6604 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5153), 
	.D(\ram[67][5] ), 
	.C(\ram[65][5] ), 
	.B(\ram[66][5] ), 
	.A(\ram[64][5] ));
   MUX4EHD U6605 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5154), 
	.D(n5150), 
	.C(n5152), 
	.B(n5151), 
	.A(n5153));
   MUX4EHD U6606 (.S1(n6038), 
	.S0(n7444), 
	.O(n5155), 
	.D(n5139), 
	.C(n5149), 
	.B(n5144), 
	.A(n5154));
   MUX4EHD U6607 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5156), 
	.D(\ram[63][5] ), 
	.C(\ram[61][5] ), 
	.B(\ram[62][5] ), 
	.A(\ram[60][5] ));
   MUX4EHD U6608 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5157), 
	.D(\ram[59][5] ), 
	.C(\ram[57][5] ), 
	.B(\ram[58][5] ), 
	.A(\ram[56][5] ));
   MUX4EHD U6609 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5158), 
	.D(\ram[55][5] ), 
	.C(\ram[53][5] ), 
	.B(\ram[54][5] ), 
	.A(\ram[52][5] ));
   MUX4EHD U6610 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5159), 
	.D(\ram[51][5] ), 
	.C(\ram[49][5] ), 
	.B(\ram[50][5] ), 
	.A(\ram[48][5] ));
   MUX4EHD U6611 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5160), 
	.D(n5156), 
	.C(n5158), 
	.B(n5157), 
	.A(n5159));
   MUX4EHD U6612 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5161), 
	.D(\ram[47][5] ), 
	.C(\ram[45][5] ), 
	.B(\ram[46][5] ), 
	.A(\ram[44][5] ));
   MUX4EHD U6613 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5162), 
	.D(\ram[43][5] ), 
	.C(\ram[41][5] ), 
	.B(\ram[42][5] ), 
	.A(\ram[40][5] ));
   MUX4EHD U6614 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5163), 
	.D(\ram[39][5] ), 
	.C(\ram[37][5] ), 
	.B(\ram[38][5] ), 
	.A(\ram[36][5] ));
   MUX4EHD U6615 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5164), 
	.D(\ram[35][5] ), 
	.C(\ram[33][5] ), 
	.B(\ram[34][5] ), 
	.A(\ram[32][5] ));
   MUX4EHD U6616 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5165), 
	.D(n5161), 
	.C(n5163), 
	.B(n5162), 
	.A(n5164));
   MUX4EHD U6617 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5166), 
	.D(\ram[31][5] ), 
	.C(\ram[29][5] ), 
	.B(\ram[30][5] ), 
	.A(\ram[28][5] ));
   MUX4EHD U6618 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5167), 
	.D(\ram[27][5] ), 
	.C(\ram[25][5] ), 
	.B(\ram[26][5] ), 
	.A(\ram[24][5] ));
   MUX4EHD U6619 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5168), 
	.D(\ram[23][5] ), 
	.C(\ram[21][5] ), 
	.B(\ram[22][5] ), 
	.A(\ram[20][5] ));
   MUX4EHD U6620 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5169), 
	.D(\ram[19][5] ), 
	.C(\ram[17][5] ), 
	.B(\ram[18][5] ), 
	.A(\ram[16][5] ));
   MUX4EHD U6621 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5170), 
	.D(n5166), 
	.C(n5168), 
	.B(n5167), 
	.A(n5169));
   MUX4EHD U6622 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5171), 
	.D(\ram[15][5] ), 
	.C(\ram[13][5] ), 
	.B(\ram[14][5] ), 
	.A(\ram[12][5] ));
   MUX4EHD U6623 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5172), 
	.D(\ram[11][5] ), 
	.C(\ram[9][5] ), 
	.B(\ram[10][5] ), 
	.A(\ram[8][5] ));
   MUX4EHD U6624 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5173), 
	.D(\ram[7][5] ), 
	.C(\ram[5][5] ), 
	.B(\ram[6][5] ), 
	.A(\ram[4][5] ));
   MUX4EHD U6625 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5174), 
	.D(\ram[3][5] ), 
	.C(\ram[1][5] ), 
	.B(\ram[2][5] ), 
	.A(\ram[0][5] ));
   MUX4EHD U6626 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5175), 
	.D(n5171), 
	.C(n5173), 
	.B(n5172), 
	.A(n5174));
   MUX4EHD U6627 (.S1(n6038), 
	.S0(n7444), 
	.O(n5176), 
	.D(n5160), 
	.C(n5170), 
	.B(n5165), 
	.A(n5175));
   MUX4EHD U6628 (.S1(n6469), 
	.S0(n6470), 
	.O(N4136), 
	.D(n5113), 
	.C(n5155), 
	.B(n5134), 
	.A(n5176));
   MUX4EHD U6629 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5177), 
	.D(\ram[255][6] ), 
	.C(\ram[253][6] ), 
	.B(\ram[254][6] ), 
	.A(\ram[252][6] ));
   MUX4EHD U6630 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5178), 
	.D(\ram[251][6] ), 
	.C(\ram[249][6] ), 
	.B(\ram[250][6] ), 
	.A(\ram[248][6] ));
   MUX4EHD U6631 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5179), 
	.D(\ram[247][6] ), 
	.C(\ram[245][6] ), 
	.B(\ram[246][6] ), 
	.A(\ram[244][6] ));
   MUX4EHD U6632 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5180), 
	.D(\ram[243][6] ), 
	.C(\ram[241][6] ), 
	.B(\ram[242][6] ), 
	.A(\ram[240][6] ));
   MUX4EHD U6633 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5181), 
	.D(n5177), 
	.C(n5179), 
	.B(n5178), 
	.A(n5180));
   MUX4EHD U6634 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5182), 
	.D(\ram[239][6] ), 
	.C(\ram[237][6] ), 
	.B(\ram[238][6] ), 
	.A(\ram[236][6] ));
   MUX4EHD U6635 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5183), 
	.D(\ram[235][6] ), 
	.C(\ram[233][6] ), 
	.B(\ram[234][6] ), 
	.A(\ram[232][6] ));
   MUX4EHD U6636 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5184), 
	.D(\ram[231][6] ), 
	.C(\ram[229][6] ), 
	.B(\ram[230][6] ), 
	.A(\ram[228][6] ));
   MUX4EHD U6637 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5185), 
	.D(\ram[227][6] ), 
	.C(\ram[225][6] ), 
	.B(\ram[226][6] ), 
	.A(\ram[224][6] ));
   MUX4EHD U6638 (.S1(n6136), 
	.S0(n7442), 
	.O(n5186), 
	.D(n5182), 
	.C(n5184), 
	.B(n5183), 
	.A(n5185));
   MUX4EHD U6639 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5187), 
	.D(\ram[223][6] ), 
	.C(\ram[221][6] ), 
	.B(\ram[222][6] ), 
	.A(\ram[220][6] ));
   MUX4EHD U6640 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5188), 
	.D(\ram[219][6] ), 
	.C(\ram[217][6] ), 
	.B(\ram[218][6] ), 
	.A(\ram[216][6] ));
   MUX4EHD U6641 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5189), 
	.D(\ram[215][6] ), 
	.C(\ram[213][6] ), 
	.B(\ram[214][6] ), 
	.A(\ram[212][6] ));
   MUX4EHD U6642 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5190), 
	.D(\ram[211][6] ), 
	.C(\ram[209][6] ), 
	.B(\ram[210][6] ), 
	.A(\ram[208][6] ));
   MUX4EHD U6643 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5191), 
	.D(n5187), 
	.C(n5189), 
	.B(n5188), 
	.A(n5190));
   MUX4EHD U6644 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5192), 
	.D(\ram[207][6] ), 
	.C(\ram[205][6] ), 
	.B(\ram[206][6] ), 
	.A(\ram[204][6] ));
   MUX4EHD U6645 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5193), 
	.D(\ram[203][6] ), 
	.C(\ram[201][6] ), 
	.B(\ram[202][6] ), 
	.A(\ram[200][6] ));
   MUX4EHD U6646 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5194), 
	.D(\ram[199][6] ), 
	.C(\ram[197][6] ), 
	.B(\ram[198][6] ), 
	.A(\ram[196][6] ));
   MUX4EHD U6647 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5195), 
	.D(\ram[195][6] ), 
	.C(\ram[193][6] ), 
	.B(\ram[194][6] ), 
	.A(\ram[192][6] ));
   MUX4EHD U6648 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5196), 
	.D(n5192), 
	.C(n5194), 
	.B(n5193), 
	.A(n5195));
   MUX4EHD U6649 (.S1(n6038), 
	.S0(n7444), 
	.O(n5197), 
	.D(n5181), 
	.C(n5191), 
	.B(n5186), 
	.A(n5196));
   MUX4EHD U6650 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5198), 
	.D(\ram[191][6] ), 
	.C(\ram[189][6] ), 
	.B(\ram[190][6] ), 
	.A(\ram[188][6] ));
   MUX4EHD U6651 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5199), 
	.D(\ram[187][6] ), 
	.C(\ram[185][6] ), 
	.B(\ram[186][6] ), 
	.A(\ram[184][6] ));
   MUX4EHD U6652 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5200), 
	.D(\ram[183][6] ), 
	.C(\ram[181][6] ), 
	.B(\ram[182][6] ), 
	.A(\ram[180][6] ));
   MUX4EHD U6653 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5201), 
	.D(\ram[179][6] ), 
	.C(\ram[177][6] ), 
	.B(\ram[178][6] ), 
	.A(\ram[176][6] ));
   MUX4EHD U6654 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5202), 
	.D(n5198), 
	.C(n5200), 
	.B(n5199), 
	.A(n5201));
   MUX4EHD U6655 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5203), 
	.D(\ram[175][6] ), 
	.C(\ram[173][6] ), 
	.B(\ram[174][6] ), 
	.A(\ram[172][6] ));
   MUX4EHD U6656 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5204), 
	.D(\ram[171][6] ), 
	.C(\ram[169][6] ), 
	.B(\ram[170][6] ), 
	.A(\ram[168][6] ));
   MUX4EHD U6657 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5205), 
	.D(\ram[167][6] ), 
	.C(\ram[165][6] ), 
	.B(\ram[166][6] ), 
	.A(\ram[164][6] ));
   MUX4EHD U6658 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5206), 
	.D(\ram[163][6] ), 
	.C(\ram[161][6] ), 
	.B(\ram[162][6] ), 
	.A(\ram[160][6] ));
   MUX4EHD U6659 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5207), 
	.D(n5203), 
	.C(n5205), 
	.B(n5204), 
	.A(n5206));
   MUX4EHD U6660 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5208), 
	.D(\ram[159][6] ), 
	.C(\ram[157][6] ), 
	.B(\ram[158][6] ), 
	.A(\ram[156][6] ));
   MUX4EHD U6661 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5209), 
	.D(\ram[155][6] ), 
	.C(\ram[153][6] ), 
	.B(\ram[154][6] ), 
	.A(\ram[152][6] ));
   MUX4EHD U6662 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5210), 
	.D(\ram[151][6] ), 
	.C(\ram[149][6] ), 
	.B(\ram[150][6] ), 
	.A(\ram[148][6] ));
   MUX4EHD U6663 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5211), 
	.D(\ram[147][6] ), 
	.C(\ram[145][6] ), 
	.B(\ram[146][6] ), 
	.A(\ram[144][6] ));
   MUX4EHD U6664 (.S1(n6136), 
	.S0(n7442), 
	.O(n5212), 
	.D(n5208), 
	.C(n5210), 
	.B(n5209), 
	.A(n5211));
   MUX4EHD U6665 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5213), 
	.D(\ram[143][6] ), 
	.C(\ram[141][6] ), 
	.B(\ram[142][6] ), 
	.A(\ram[140][6] ));
   MUX4EHD U6666 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5214), 
	.D(\ram[139][6] ), 
	.C(\ram[137][6] ), 
	.B(\ram[138][6] ), 
	.A(\ram[136][6] ));
   MUX4EHD U6667 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5215), 
	.D(\ram[135][6] ), 
	.C(\ram[133][6] ), 
	.B(\ram[134][6] ), 
	.A(\ram[132][6] ));
   MUX4EHD U6668 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5216), 
	.D(\ram[131][6] ), 
	.C(\ram[129][6] ), 
	.B(\ram[130][6] ), 
	.A(\ram[128][6] ));
   MUX4EHD U6669 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5217), 
	.D(n5213), 
	.C(n5215), 
	.B(n5214), 
	.A(n5216));
   MUX4EHD U6670 (.S1(n6038), 
	.S0(n7444), 
	.O(n5218), 
	.D(n5202), 
	.C(n5212), 
	.B(n5207), 
	.A(n5217));
   MUX4EHD U6671 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5219), 
	.D(\ram[127][6] ), 
	.C(\ram[125][6] ), 
	.B(\ram[126][6] ), 
	.A(\ram[124][6] ));
   MUX4EHD U6672 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5220), 
	.D(\ram[123][6] ), 
	.C(\ram[121][6] ), 
	.B(\ram[122][6] ), 
	.A(\ram[120][6] ));
   MUX4EHD U6673 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5221), 
	.D(\ram[119][6] ), 
	.C(\ram[117][6] ), 
	.B(\ram[118][6] ), 
	.A(\ram[116][6] ));
   MUX4EHD U6674 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5222), 
	.D(\ram[115][6] ), 
	.C(\ram[113][6] ), 
	.B(\ram[114][6] ), 
	.A(\ram[112][6] ));
   MUX4EHD U6675 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5223), 
	.D(n5219), 
	.C(n5221), 
	.B(n5220), 
	.A(n5222));
   MUX4EHD U6676 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5224), 
	.D(\ram[111][6] ), 
	.C(\ram[109][6] ), 
	.B(\ram[110][6] ), 
	.A(\ram[108][6] ));
   MUX4EHD U6677 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5225), 
	.D(\ram[107][6] ), 
	.C(\ram[105][6] ), 
	.B(\ram[106][6] ), 
	.A(\ram[104][6] ));
   MUX4EHD U6678 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5226), 
	.D(\ram[103][6] ), 
	.C(\ram[101][6] ), 
	.B(\ram[102][6] ), 
	.A(\ram[100][6] ));
   MUX4EHD U6679 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5227), 
	.D(\ram[99][6] ), 
	.C(\ram[97][6] ), 
	.B(\ram[98][6] ), 
	.A(\ram[96][6] ));
   MUX4EHD U6680 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5228), 
	.D(n5224), 
	.C(n5226), 
	.B(n5225), 
	.A(n5227));
   MUX4EHD U6681 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5229), 
	.D(\ram[95][6] ), 
	.C(\ram[93][6] ), 
	.B(\ram[94][6] ), 
	.A(\ram[92][6] ));
   MUX4EHD U6682 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5230), 
	.D(\ram[91][6] ), 
	.C(\ram[89][6] ), 
	.B(\ram[90][6] ), 
	.A(\ram[88][6] ));
   MUX4EHD U6683 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5231), 
	.D(\ram[87][6] ), 
	.C(\ram[85][6] ), 
	.B(\ram[86][6] ), 
	.A(\ram[84][6] ));
   MUX4EHD U6684 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5232), 
	.D(\ram[83][6] ), 
	.C(\ram[81][6] ), 
	.B(\ram[82][6] ), 
	.A(\ram[80][6] ));
   MUX4EHD U6685 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5233), 
	.D(n5229), 
	.C(n5231), 
	.B(n5230), 
	.A(n5232));
   MUX4EHD U6686 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5234), 
	.D(\ram[79][6] ), 
	.C(\ram[77][6] ), 
	.B(\ram[78][6] ), 
	.A(\ram[76][6] ));
   MUX4EHD U6687 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5235), 
	.D(\ram[75][6] ), 
	.C(\ram[73][6] ), 
	.B(\ram[74][6] ), 
	.A(\ram[72][6] ));
   MUX4EHD U6688 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5236), 
	.D(\ram[71][6] ), 
	.C(\ram[69][6] ), 
	.B(\ram[70][6] ), 
	.A(\ram[68][6] ));
   MUX4EHD U6689 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5237), 
	.D(\ram[67][6] ), 
	.C(\ram[65][6] ), 
	.B(\ram[66][6] ), 
	.A(\ram[64][6] ));
   MUX4EHD U6690 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5238), 
	.D(n5234), 
	.C(n5236), 
	.B(n5235), 
	.A(n5237));
   MUX4EHD U6691 (.S1(n6038), 
	.S0(n7444), 
	.O(n5239), 
	.D(n5223), 
	.C(n5233), 
	.B(n5228), 
	.A(n5238));
   MUX4EHD U6692 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5240), 
	.D(\ram[63][6] ), 
	.C(\ram[61][6] ), 
	.B(\ram[62][6] ), 
	.A(\ram[60][6] ));
   MUX4EHD U6693 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5241), 
	.D(\ram[59][6] ), 
	.C(\ram[57][6] ), 
	.B(\ram[58][6] ), 
	.A(\ram[56][6] ));
   MUX4EHD U6694 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5242), 
	.D(\ram[55][6] ), 
	.C(\ram[53][6] ), 
	.B(\ram[54][6] ), 
	.A(\ram[52][6] ));
   MUX4EHD U6695 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5243), 
	.D(\ram[51][6] ), 
	.C(\ram[49][6] ), 
	.B(\ram[50][6] ), 
	.A(\ram[48][6] ));
   MUX4EHD U6696 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5244), 
	.D(n5240), 
	.C(n5242), 
	.B(n5241), 
	.A(n5243));
   MUX4EHD U6697 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5245), 
	.D(\ram[47][6] ), 
	.C(\ram[45][6] ), 
	.B(\ram[46][6] ), 
	.A(\ram[44][6] ));
   MUX4EHD U6698 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5246), 
	.D(\ram[43][6] ), 
	.C(\ram[41][6] ), 
	.B(\ram[42][6] ), 
	.A(\ram[40][6] ));
   MUX4EHD U6699 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5247), 
	.D(\ram[39][6] ), 
	.C(\ram[37][6] ), 
	.B(\ram[38][6] ), 
	.A(\ram[36][6] ));
   MUX4EHD U6700 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5248), 
	.D(\ram[35][6] ), 
	.C(\ram[33][6] ), 
	.B(\ram[34][6] ), 
	.A(\ram[32][6] ));
   MUX4EHD U6701 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5249), 
	.D(n5245), 
	.C(n5247), 
	.B(n5246), 
	.A(n5248));
   MUX4EHD U6702 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5250), 
	.D(\ram[31][6] ), 
	.C(\ram[29][6] ), 
	.B(\ram[30][6] ), 
	.A(\ram[28][6] ));
   MUX4EHD U6703 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5251), 
	.D(\ram[27][6] ), 
	.C(\ram[25][6] ), 
	.B(\ram[26][6] ), 
	.A(\ram[24][6] ));
   MUX4EHD U6704 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5252), 
	.D(\ram[23][6] ), 
	.C(\ram[21][6] ), 
	.B(\ram[22][6] ), 
	.A(\ram[20][6] ));
   MUX4EHD U6705 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5253), 
	.D(\ram[19][6] ), 
	.C(\ram[17][6] ), 
	.B(\ram[18][6] ), 
	.A(\ram[16][6] ));
   MUX4EHD U6706 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5254), 
	.D(n5250), 
	.C(n5252), 
	.B(n5251), 
	.A(n5253));
   MUX4EHD U6707 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5255), 
	.D(\ram[15][6] ), 
	.C(\ram[13][6] ), 
	.B(\ram[14][6] ), 
	.A(\ram[12][6] ));
   MUX4EHD U6708 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5256), 
	.D(\ram[11][6] ), 
	.C(\ram[9][6] ), 
	.B(\ram[10][6] ), 
	.A(\ram[8][6] ));
   MUX4EHD U6709 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5257), 
	.D(\ram[7][6] ), 
	.C(\ram[5][6] ), 
	.B(\ram[6][6] ), 
	.A(\ram[4][6] ));
   MUX4EHD U6710 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5258), 
	.D(\ram[3][6] ), 
	.C(\ram[1][6] ), 
	.B(\ram[2][6] ), 
	.A(\ram[0][6] ));
   MUX4EHD U6711 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5259), 
	.D(n5255), 
	.C(n5257), 
	.B(n5256), 
	.A(n5258));
   MUX4EHD U6712 (.S1(n6038), 
	.S0(n7444), 
	.O(n5260), 
	.D(n5244), 
	.C(n5254), 
	.B(n5249), 
	.A(n5259));
   MUX4EHD U6713 (.S1(n6469), 
	.S0(n6470), 
	.O(N4135), 
	.D(n5197), 
	.C(n5239), 
	.B(n5218), 
	.A(n5260));
   MUX4EHD U6714 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5261), 
	.D(\ram[255][7] ), 
	.C(\ram[253][7] ), 
	.B(\ram[254][7] ), 
	.A(\ram[252][7] ));
   MUX4EHD U6715 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5262), 
	.D(\ram[251][7] ), 
	.C(\ram[249][7] ), 
	.B(\ram[250][7] ), 
	.A(\ram[248][7] ));
   MUX4EHD U6716 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5263), 
	.D(\ram[247][7] ), 
	.C(\ram[245][7] ), 
	.B(\ram[246][7] ), 
	.A(\ram[244][7] ));
   MUX4EHD U6717 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5264), 
	.D(\ram[243][7] ), 
	.C(\ram[241][7] ), 
	.B(\ram[242][7] ), 
	.A(\ram[240][7] ));
   MUX4EHD U6718 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5265), 
	.D(n5261), 
	.C(n5263), 
	.B(n5262), 
	.A(n5264));
   MUX4EHD U6719 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5266), 
	.D(\ram[239][7] ), 
	.C(\ram[237][7] ), 
	.B(\ram[238][7] ), 
	.A(\ram[236][7] ));
   MUX4EHD U6720 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5267), 
	.D(\ram[235][7] ), 
	.C(\ram[233][7] ), 
	.B(\ram[234][7] ), 
	.A(\ram[232][7] ));
   MUX4EHD U6721 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5268), 
	.D(\ram[231][7] ), 
	.C(\ram[229][7] ), 
	.B(\ram[230][7] ), 
	.A(\ram[228][7] ));
   MUX4EHD U6722 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5269), 
	.D(\ram[227][7] ), 
	.C(\ram[225][7] ), 
	.B(\ram[226][7] ), 
	.A(\ram[224][7] ));
   MUX4EHD U6723 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5270), 
	.D(n5266), 
	.C(n5268), 
	.B(n5267), 
	.A(n5269));
   MUX4EHD U6724 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5271), 
	.D(\ram[223][7] ), 
	.C(\ram[221][7] ), 
	.B(\ram[222][7] ), 
	.A(\ram[220][7] ));
   MUX4EHD U6725 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5272), 
	.D(\ram[219][7] ), 
	.C(\ram[217][7] ), 
	.B(\ram[218][7] ), 
	.A(\ram[216][7] ));
   MUX4EHD U6726 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5273), 
	.D(\ram[215][7] ), 
	.C(\ram[213][7] ), 
	.B(\ram[214][7] ), 
	.A(\ram[212][7] ));
   MUX4EHD U6727 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5274), 
	.D(\ram[211][7] ), 
	.C(\ram[209][7] ), 
	.B(\ram[210][7] ), 
	.A(\ram[208][7] ));
   MUX4EHD U6728 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5275), 
	.D(n5271), 
	.C(n5273), 
	.B(n5272), 
	.A(n5274));
   MUX4EHD U6729 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5276), 
	.D(\ram[207][7] ), 
	.C(\ram[205][7] ), 
	.B(\ram[206][7] ), 
	.A(\ram[204][7] ));
   MUX4EHD U6730 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5277), 
	.D(\ram[203][7] ), 
	.C(\ram[201][7] ), 
	.B(\ram[202][7] ), 
	.A(\ram[200][7] ));
   MUX4EHD U6731 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5278), 
	.D(\ram[199][7] ), 
	.C(\ram[197][7] ), 
	.B(\ram[198][7] ), 
	.A(\ram[196][7] ));
   MUX4EHD U6732 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5279), 
	.D(\ram[195][7] ), 
	.C(\ram[193][7] ), 
	.B(\ram[194][7] ), 
	.A(\ram[192][7] ));
   MUX4EHD U6733 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5280), 
	.D(n5276), 
	.C(n5278), 
	.B(n5277), 
	.A(n5279));
   MUX4EHD U6734 (.S1(n6038), 
	.S0(n7444), 
	.O(n5281), 
	.D(n5265), 
	.C(n5275), 
	.B(n5270), 
	.A(n5280));
   MUX4EHD U6735 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5282), 
	.D(\ram[191][7] ), 
	.C(\ram[189][7] ), 
	.B(\ram[190][7] ), 
	.A(\ram[188][7] ));
   MUX4EHD U6736 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5283), 
	.D(\ram[187][7] ), 
	.C(\ram[185][7] ), 
	.B(\ram[186][7] ), 
	.A(\ram[184][7] ));
   MUX4EHD U6737 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5284), 
	.D(\ram[183][7] ), 
	.C(\ram[181][7] ), 
	.B(\ram[182][7] ), 
	.A(\ram[180][7] ));
   MUX4EHD U6738 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5285), 
	.D(\ram[179][7] ), 
	.C(\ram[177][7] ), 
	.B(\ram[178][7] ), 
	.A(\ram[176][7] ));
   MUX4EHD U6739 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5286), 
	.D(n5282), 
	.C(n5284), 
	.B(n5283), 
	.A(n5285));
   MUX4EHD U6740 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5287), 
	.D(\ram[175][7] ), 
	.C(\ram[173][7] ), 
	.B(\ram[174][7] ), 
	.A(\ram[172][7] ));
   MUX4EHD U6741 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5288), 
	.D(\ram[171][7] ), 
	.C(\ram[169][7] ), 
	.B(\ram[170][7] ), 
	.A(\ram[168][7] ));
   MUX4EHD U6742 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5289), 
	.D(\ram[167][7] ), 
	.C(\ram[165][7] ), 
	.B(\ram[166][7] ), 
	.A(\ram[164][7] ));
   MUX4EHD U6743 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5290), 
	.D(\ram[163][7] ), 
	.C(\ram[161][7] ), 
	.B(\ram[162][7] ), 
	.A(\ram[160][7] ));
   MUX4EHD U6744 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5291), 
	.D(n5287), 
	.C(n5289), 
	.B(n5288), 
	.A(n5290));
   MUX4EHD U6745 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5292), 
	.D(\ram[159][7] ), 
	.C(\ram[157][7] ), 
	.B(\ram[158][7] ), 
	.A(\ram[156][7] ));
   MUX4EHD U6746 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n5293), 
	.D(\ram[155][7] ), 
	.C(\ram[153][7] ), 
	.B(\ram[154][7] ), 
	.A(\ram[152][7] ));
   MUX4EHD U6747 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5294), 
	.D(\ram[151][7] ), 
	.C(\ram[149][7] ), 
	.B(\ram[150][7] ), 
	.A(\ram[148][7] ));
   MUX4EHD U6748 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5295), 
	.D(\ram[147][7] ), 
	.C(\ram[145][7] ), 
	.B(\ram[146][7] ), 
	.A(\ram[144][7] ));
   MUX4EHD U6749 (.S1(n6136), 
	.S0(n7442), 
	.O(n5296), 
	.D(n5292), 
	.C(n5294), 
	.B(n5293), 
	.A(n5295));
   MUX4EHD U6750 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5297), 
	.D(\ram[143][7] ), 
	.C(\ram[141][7] ), 
	.B(\ram[142][7] ), 
	.A(\ram[140][7] ));
   MUX4EHD U6751 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5298), 
	.D(\ram[139][7] ), 
	.C(\ram[137][7] ), 
	.B(\ram[138][7] ), 
	.A(\ram[136][7] ));
   MUX4EHD U6752 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5299), 
	.D(\ram[135][7] ), 
	.C(\ram[133][7] ), 
	.B(\ram[134][7] ), 
	.A(\ram[132][7] ));
   MUX4EHD U6753 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5300), 
	.D(\ram[131][7] ), 
	.C(\ram[129][7] ), 
	.B(\ram[130][7] ), 
	.A(\ram[128][7] ));
   MUX4EHD U6754 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5301), 
	.D(n5297), 
	.C(n5299), 
	.B(n5298), 
	.A(n5300));
   MUX4EHD U6755 (.S1(n6038), 
	.S0(n7444), 
	.O(n5302), 
	.D(n5286), 
	.C(n5296), 
	.B(n5291), 
	.A(n5301));
   MUX4EHD U6756 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5303), 
	.D(\ram[127][7] ), 
	.C(\ram[125][7] ), 
	.B(\ram[126][7] ), 
	.A(\ram[124][7] ));
   MUX4EHD U6757 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5304), 
	.D(\ram[123][7] ), 
	.C(\ram[121][7] ), 
	.B(\ram[122][7] ), 
	.A(\ram[120][7] ));
   MUX4EHD U6758 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5305), 
	.D(\ram[119][7] ), 
	.C(\ram[117][7] ), 
	.B(\ram[118][7] ), 
	.A(\ram[116][7] ));
   MUX4EHD U6759 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5306), 
	.D(\ram[115][7] ), 
	.C(\ram[113][7] ), 
	.B(\ram[114][7] ), 
	.A(\ram[112][7] ));
   MUX4EHD U6760 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5307), 
	.D(n5303), 
	.C(n5305), 
	.B(n5304), 
	.A(n5306));
   MUX4EHD U6761 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5308), 
	.D(\ram[111][7] ), 
	.C(\ram[109][7] ), 
	.B(\ram[110][7] ), 
	.A(\ram[108][7] ));
   MUX4EHD U6762 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5309), 
	.D(\ram[107][7] ), 
	.C(\ram[105][7] ), 
	.B(\ram[106][7] ), 
	.A(\ram[104][7] ));
   MUX4EHD U6763 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5310), 
	.D(\ram[103][7] ), 
	.C(\ram[101][7] ), 
	.B(\ram[102][7] ), 
	.A(\ram[100][7] ));
   MUX4EHD U6764 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5311), 
	.D(\ram[99][7] ), 
	.C(\ram[97][7] ), 
	.B(\ram[98][7] ), 
	.A(\ram[96][7] ));
   MUX4EHD U6765 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5312), 
	.D(n5308), 
	.C(n5310), 
	.B(n5309), 
	.A(n5311));
   MUX4EHD U6766 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5313), 
	.D(\ram[95][7] ), 
	.C(\ram[93][7] ), 
	.B(\ram[94][7] ), 
	.A(\ram[92][7] ));
   MUX4EHD U6767 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5314), 
	.D(\ram[91][7] ), 
	.C(\ram[89][7] ), 
	.B(\ram[90][7] ), 
	.A(\ram[88][7] ));
   MUX4EHD U6768 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5315), 
	.D(\ram[87][7] ), 
	.C(\ram[85][7] ), 
	.B(\ram[86][7] ), 
	.A(\ram[84][7] ));
   MUX4EHD U6769 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5316), 
	.D(\ram[83][7] ), 
	.C(\ram[81][7] ), 
	.B(\ram[82][7] ), 
	.A(\ram[80][7] ));
   MUX4EHD U6770 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5317), 
	.D(n5313), 
	.C(n5315), 
	.B(n5314), 
	.A(n5316));
   MUX4EHD U6771 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5318), 
	.D(\ram[79][7] ), 
	.C(\ram[77][7] ), 
	.B(\ram[78][7] ), 
	.A(\ram[76][7] ));
   MUX4EHD U6772 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5319), 
	.D(\ram[75][7] ), 
	.C(\ram[73][7] ), 
	.B(\ram[74][7] ), 
	.A(\ram[72][7] ));
   MUX4EHD U6773 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5320), 
	.D(\ram[71][7] ), 
	.C(\ram[69][7] ), 
	.B(\ram[70][7] ), 
	.A(\ram[68][7] ));
   MUX4EHD U6774 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5321), 
	.D(\ram[67][7] ), 
	.C(\ram[65][7] ), 
	.B(\ram[66][7] ), 
	.A(\ram[64][7] ));
   MUX4EHD U6775 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5322), 
	.D(n5318), 
	.C(n5320), 
	.B(n5319), 
	.A(n5321));
   MUX4EHD U6776 (.S1(n6038), 
	.S0(n7444), 
	.O(n5323), 
	.D(n5307), 
	.C(n5317), 
	.B(n5312), 
	.A(n5322));
   MUX4EHD U6777 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5324), 
	.D(\ram[63][7] ), 
	.C(\ram[61][7] ), 
	.B(\ram[62][7] ), 
	.A(\ram[60][7] ));
   MUX4EHD U6778 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5325), 
	.D(\ram[59][7] ), 
	.C(\ram[57][7] ), 
	.B(\ram[58][7] ), 
	.A(\ram[56][7] ));
   MUX4EHD U6779 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5326), 
	.D(\ram[55][7] ), 
	.C(\ram[53][7] ), 
	.B(\ram[54][7] ), 
	.A(\ram[52][7] ));
   MUX4EHD U6780 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5327), 
	.D(\ram[51][7] ), 
	.C(\ram[49][7] ), 
	.B(\ram[50][7] ), 
	.A(\ram[48][7] ));
   MUX4EHD U6781 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5328), 
	.D(n5324), 
	.C(n5326), 
	.B(n5325), 
	.A(n5327));
   MUX4EHD U6782 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5329), 
	.D(\ram[47][7] ), 
	.C(\ram[45][7] ), 
	.B(\ram[46][7] ), 
	.A(\ram[44][7] ));
   MUX4EHD U6783 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5330), 
	.D(\ram[43][7] ), 
	.C(\ram[41][7] ), 
	.B(\ram[42][7] ), 
	.A(\ram[40][7] ));
   MUX4EHD U6784 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5331), 
	.D(\ram[39][7] ), 
	.C(\ram[37][7] ), 
	.B(\ram[38][7] ), 
	.A(\ram[36][7] ));
   MUX4EHD U6785 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5332), 
	.D(\ram[35][7] ), 
	.C(\ram[33][7] ), 
	.B(\ram[34][7] ), 
	.A(\ram[32][7] ));
   MUX4EHD U6786 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5333), 
	.D(n5329), 
	.C(n5331), 
	.B(n5330), 
	.A(n5332));
   MUX4EHD U6787 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5334), 
	.D(\ram[31][7] ), 
	.C(\ram[29][7] ), 
	.B(\ram[30][7] ), 
	.A(\ram[28][7] ));
   MUX4EHD U6788 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5335), 
	.D(\ram[27][7] ), 
	.C(\ram[25][7] ), 
	.B(\ram[26][7] ), 
	.A(\ram[24][7] ));
   MUX4EHD U6789 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5336), 
	.D(\ram[23][7] ), 
	.C(\ram[21][7] ), 
	.B(\ram[22][7] ), 
	.A(\ram[20][7] ));
   MUX4EHD U6790 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5337), 
	.D(\ram[19][7] ), 
	.C(\ram[17][7] ), 
	.B(\ram[18][7] ), 
	.A(\ram[16][7] ));
   MUX4EHD U6791 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5338), 
	.D(n5334), 
	.C(n5336), 
	.B(n5335), 
	.A(n5337));
   MUX4EHD U6792 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5339), 
	.D(\ram[15][7] ), 
	.C(\ram[13][7] ), 
	.B(\ram[14][7] ), 
	.A(\ram[12][7] ));
   MUX4EHD U6793 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5340), 
	.D(\ram[11][7] ), 
	.C(\ram[9][7] ), 
	.B(\ram[10][7] ), 
	.A(\ram[8][7] ));
   MUX4EHD U6794 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5341), 
	.D(\ram[7][7] ), 
	.C(\ram[5][7] ), 
	.B(\ram[6][7] ), 
	.A(\ram[4][7] ));
   MUX4EHD U6795 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5342), 
	.D(\ram[3][7] ), 
	.C(\ram[1][7] ), 
	.B(\ram[2][7] ), 
	.A(\ram[0][7] ));
   MUX4EHD U6796 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5343), 
	.D(n5339), 
	.C(n5341), 
	.B(n5340), 
	.A(n5342));
   MUX4EHD U6797 (.S1(n6038), 
	.S0(n7444), 
	.O(n5344), 
	.D(n5328), 
	.C(n5338), 
	.B(n5333), 
	.A(n5343));
   MUX4EHD U6798 (.S1(n6469), 
	.S0(n6470), 
	.O(N4134), 
	.D(n5281), 
	.C(n5323), 
	.B(n5302), 
	.A(n5344));
   MUX4EHD U6799 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5345), 
	.D(\ram[255][8] ), 
	.C(\ram[253][8] ), 
	.B(\ram[254][8] ), 
	.A(\ram[252][8] ));
   MUX4EHD U6800 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5346), 
	.D(\ram[251][8] ), 
	.C(\ram[249][8] ), 
	.B(\ram[250][8] ), 
	.A(\ram[248][8] ));
   MUX4EHD U6801 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5347), 
	.D(\ram[247][8] ), 
	.C(\ram[245][8] ), 
	.B(\ram[246][8] ), 
	.A(\ram[244][8] ));
   MUX4EHD U6802 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5348), 
	.D(\ram[243][8] ), 
	.C(\ram[241][8] ), 
	.B(\ram[242][8] ), 
	.A(\ram[240][8] ));
   MUX4EHD U6803 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5349), 
	.D(n5345), 
	.C(n5347), 
	.B(n5346), 
	.A(n5348));
   MUX4EHD U6804 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5350), 
	.D(\ram[239][8] ), 
	.C(\ram[237][8] ), 
	.B(\ram[238][8] ), 
	.A(\ram[236][8] ));
   MUX4EHD U6805 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5351), 
	.D(\ram[235][8] ), 
	.C(\ram[233][8] ), 
	.B(\ram[234][8] ), 
	.A(\ram[232][8] ));
   MUX4EHD U6806 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5352), 
	.D(\ram[231][8] ), 
	.C(\ram[229][8] ), 
	.B(\ram[230][8] ), 
	.A(\ram[228][8] ));
   MUX4EHD U6807 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5353), 
	.D(\ram[227][8] ), 
	.C(\ram[225][8] ), 
	.B(\ram[226][8] ), 
	.A(\ram[224][8] ));
   MUX4EHD U6808 (.S1(n6136), 
	.S0(n7442), 
	.O(n5354), 
	.D(n5350), 
	.C(n5352), 
	.B(n5351), 
	.A(n5353));
   MUX4EHD U6809 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5355), 
	.D(\ram[223][8] ), 
	.C(\ram[221][8] ), 
	.B(\ram[222][8] ), 
	.A(\ram[220][8] ));
   MUX4EHD U6810 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5356), 
	.D(\ram[219][8] ), 
	.C(\ram[217][8] ), 
	.B(\ram[218][8] ), 
	.A(\ram[216][8] ));
   MUX4EHD U6811 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5357), 
	.D(\ram[215][8] ), 
	.C(\ram[213][8] ), 
	.B(\ram[214][8] ), 
	.A(\ram[212][8] ));
   MUX4EHD U6812 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5358), 
	.D(\ram[211][8] ), 
	.C(\ram[209][8] ), 
	.B(\ram[210][8] ), 
	.A(\ram[208][8] ));
   MUX4EHD U6813 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5359), 
	.D(n5355), 
	.C(n5357), 
	.B(n5356), 
	.A(n5358));
   MUX4EHD U6814 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5360), 
	.D(\ram[207][8] ), 
	.C(\ram[205][8] ), 
	.B(\ram[206][8] ), 
	.A(\ram[204][8] ));
   MUX4EHD U6815 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5361), 
	.D(\ram[203][8] ), 
	.C(\ram[201][8] ), 
	.B(\ram[202][8] ), 
	.A(\ram[200][8] ));
   MUX4EHD U6816 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5362), 
	.D(\ram[199][8] ), 
	.C(\ram[197][8] ), 
	.B(\ram[198][8] ), 
	.A(\ram[196][8] ));
   MUX4EHD U6817 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5363), 
	.D(\ram[195][8] ), 
	.C(\ram[193][8] ), 
	.B(\ram[194][8] ), 
	.A(\ram[192][8] ));
   MUX4EHD U6818 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5364), 
	.D(n5360), 
	.C(n5362), 
	.B(n5361), 
	.A(n5363));
   MUX4EHD U6819 (.S1(n6038), 
	.S0(n7444), 
	.O(n5365), 
	.D(n5349), 
	.C(n5359), 
	.B(n5354), 
	.A(n5364));
   MUX4EHD U6820 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5366), 
	.D(\ram[191][8] ), 
	.C(\ram[189][8] ), 
	.B(\ram[190][8] ), 
	.A(\ram[188][8] ));
   MUX4EHD U6821 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5367), 
	.D(\ram[187][8] ), 
	.C(\ram[185][8] ), 
	.B(\ram[186][8] ), 
	.A(\ram[184][8] ));
   MUX4EHD U6822 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5368), 
	.D(\ram[183][8] ), 
	.C(\ram[181][8] ), 
	.B(\ram[182][8] ), 
	.A(\ram[180][8] ));
   MUX4EHD U6823 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5369), 
	.D(\ram[179][8] ), 
	.C(\ram[177][8] ), 
	.B(\ram[178][8] ), 
	.A(\ram[176][8] ));
   MUX4EHD U6824 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5370), 
	.D(n5366), 
	.C(n5368), 
	.B(n5367), 
	.A(n5369));
   MUX4EHD U6825 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5371), 
	.D(\ram[175][8] ), 
	.C(\ram[173][8] ), 
	.B(\ram[174][8] ), 
	.A(\ram[172][8] ));
   MUX4EHD U6826 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5372), 
	.D(\ram[171][8] ), 
	.C(\ram[169][8] ), 
	.B(\ram[170][8] ), 
	.A(\ram[168][8] ));
   MUX4EHD U6827 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5373), 
	.D(\ram[167][8] ), 
	.C(\ram[165][8] ), 
	.B(\ram[166][8] ), 
	.A(\ram[164][8] ));
   MUX4EHD U6828 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5374), 
	.D(\ram[163][8] ), 
	.C(\ram[161][8] ), 
	.B(\ram[162][8] ), 
	.A(\ram[160][8] ));
   MUX4EHD U6829 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5375), 
	.D(n5371), 
	.C(n5373), 
	.B(n5372), 
	.A(n5374));
   MUX4EHD U6830 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5376), 
	.D(\ram[159][8] ), 
	.C(\ram[157][8] ), 
	.B(\ram[158][8] ), 
	.A(\ram[156][8] ));
   MUX4EHD U6831 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5377), 
	.D(\ram[155][8] ), 
	.C(\ram[153][8] ), 
	.B(\ram[154][8] ), 
	.A(\ram[152][8] ));
   MUX4EHD U6832 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5378), 
	.D(\ram[151][8] ), 
	.C(\ram[149][8] ), 
	.B(\ram[150][8] ), 
	.A(\ram[148][8] ));
   MUX4EHD U6833 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5379), 
	.D(\ram[147][8] ), 
	.C(\ram[145][8] ), 
	.B(\ram[146][8] ), 
	.A(\ram[144][8] ));
   MUX4EHD U6834 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5380), 
	.D(n5376), 
	.C(n5378), 
	.B(n5377), 
	.A(n5379));
   MUX4EHD U6835 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5381), 
	.D(\ram[143][8] ), 
	.C(\ram[141][8] ), 
	.B(\ram[142][8] ), 
	.A(\ram[140][8] ));
   MUX4EHD U6836 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5382), 
	.D(\ram[139][8] ), 
	.C(\ram[137][8] ), 
	.B(\ram[138][8] ), 
	.A(\ram[136][8] ));
   MUX4EHD U6837 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5383), 
	.D(\ram[135][8] ), 
	.C(\ram[133][8] ), 
	.B(\ram[134][8] ), 
	.A(\ram[132][8] ));
   MUX4EHD U6838 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5384), 
	.D(\ram[131][8] ), 
	.C(\ram[129][8] ), 
	.B(\ram[130][8] ), 
	.A(\ram[128][8] ));
   MUX4EHD U6839 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5385), 
	.D(n5381), 
	.C(n5383), 
	.B(n5382), 
	.A(n5384));
   MUX4EHD U6840 (.S1(n6038), 
	.S0(n7444), 
	.O(n5386), 
	.D(n5370), 
	.C(n5380), 
	.B(n5375), 
	.A(n5385));
   MUX4EHD U6841 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5387), 
	.D(\ram[127][8] ), 
	.C(\ram[125][8] ), 
	.B(\ram[126][8] ), 
	.A(\ram[124][8] ));
   MUX4EHD U6842 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5388), 
	.D(\ram[123][8] ), 
	.C(\ram[121][8] ), 
	.B(\ram[122][8] ), 
	.A(\ram[120][8] ));
   MUX4EHD U6843 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5389), 
	.D(\ram[119][8] ), 
	.C(\ram[117][8] ), 
	.B(\ram[118][8] ), 
	.A(\ram[116][8] ));
   MUX4EHD U6844 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5390), 
	.D(\ram[115][8] ), 
	.C(\ram[113][8] ), 
	.B(\ram[114][8] ), 
	.A(\ram[112][8] ));
   MUX4EHD U6845 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5391), 
	.D(n5387), 
	.C(n5389), 
	.B(n5388), 
	.A(n5390));
   MUX4EHD U6846 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5392), 
	.D(\ram[111][8] ), 
	.C(\ram[109][8] ), 
	.B(\ram[110][8] ), 
	.A(\ram[108][8] ));
   MUX4EHD U6847 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5393), 
	.D(\ram[107][8] ), 
	.C(\ram[105][8] ), 
	.B(\ram[106][8] ), 
	.A(\ram[104][8] ));
   MUX4EHD U6848 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5394), 
	.D(\ram[103][8] ), 
	.C(\ram[101][8] ), 
	.B(\ram[102][8] ), 
	.A(\ram[100][8] ));
   MUX4EHD U6849 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5395), 
	.D(\ram[99][8] ), 
	.C(\ram[97][8] ), 
	.B(\ram[98][8] ), 
	.A(\ram[96][8] ));
   MUX4EHD U6850 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5396), 
	.D(n5392), 
	.C(n5394), 
	.B(n5393), 
	.A(n5395));
   MUX4EHD U6851 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5397), 
	.D(\ram[95][8] ), 
	.C(\ram[93][8] ), 
	.B(\ram[94][8] ), 
	.A(\ram[92][8] ));
   MUX4EHD U6852 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5398), 
	.D(\ram[91][8] ), 
	.C(\ram[89][8] ), 
	.B(\ram[90][8] ), 
	.A(\ram[88][8] ));
   MUX4EHD U6853 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5399), 
	.D(\ram[87][8] ), 
	.C(\ram[85][8] ), 
	.B(\ram[86][8] ), 
	.A(\ram[84][8] ));
   MUX4EHD U6854 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5400), 
	.D(\ram[83][8] ), 
	.C(\ram[81][8] ), 
	.B(\ram[82][8] ), 
	.A(\ram[80][8] ));
   MUX4EHD U6855 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5401), 
	.D(n5397), 
	.C(n5399), 
	.B(n5398), 
	.A(n5400));
   MUX4EHD U6856 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5402), 
	.D(\ram[79][8] ), 
	.C(\ram[77][8] ), 
	.B(\ram[78][8] ), 
	.A(\ram[76][8] ));
   MUX4EHD U6857 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5403), 
	.D(\ram[75][8] ), 
	.C(\ram[73][8] ), 
	.B(\ram[74][8] ), 
	.A(\ram[72][8] ));
   MUX4EHD U6858 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5404), 
	.D(\ram[71][8] ), 
	.C(\ram[69][8] ), 
	.B(\ram[70][8] ), 
	.A(\ram[68][8] ));
   MUX4EHD U6859 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5405), 
	.D(\ram[67][8] ), 
	.C(\ram[65][8] ), 
	.B(\ram[66][8] ), 
	.A(\ram[64][8] ));
   MUX4EHD U6860 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5406), 
	.D(n5402), 
	.C(n5404), 
	.B(n5403), 
	.A(n5405));
   MUX4EHD U6861 (.S1(n6038), 
	.S0(n7444), 
	.O(n5407), 
	.D(n5391), 
	.C(n5401), 
	.B(n5396), 
	.A(n5406));
   MUX4EHD U6862 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5408), 
	.D(\ram[63][8] ), 
	.C(\ram[61][8] ), 
	.B(\ram[62][8] ), 
	.A(\ram[60][8] ));
   MUX4EHD U6863 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5409), 
	.D(\ram[59][8] ), 
	.C(\ram[57][8] ), 
	.B(\ram[58][8] ), 
	.A(\ram[56][8] ));
   MUX4EHD U6864 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5410), 
	.D(\ram[55][8] ), 
	.C(\ram[53][8] ), 
	.B(\ram[54][8] ), 
	.A(\ram[52][8] ));
   MUX4EHD U6865 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5411), 
	.D(\ram[51][8] ), 
	.C(\ram[49][8] ), 
	.B(\ram[50][8] ), 
	.A(\ram[48][8] ));
   MUX4EHD U6866 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5412), 
	.D(n5408), 
	.C(n5410), 
	.B(n5409), 
	.A(n5411));
   MUX4EHD U6867 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5413), 
	.D(\ram[47][8] ), 
	.C(\ram[45][8] ), 
	.B(\ram[46][8] ), 
	.A(\ram[44][8] ));
   MUX4EHD U6868 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5414), 
	.D(\ram[43][8] ), 
	.C(\ram[41][8] ), 
	.B(\ram[42][8] ), 
	.A(\ram[40][8] ));
   MUX4EHD U6869 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5415), 
	.D(\ram[39][8] ), 
	.C(\ram[37][8] ), 
	.B(\ram[38][8] ), 
	.A(\ram[36][8] ));
   MUX4EHD U6870 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5416), 
	.D(\ram[35][8] ), 
	.C(\ram[33][8] ), 
	.B(\ram[34][8] ), 
	.A(\ram[32][8] ));
   MUX4EHD U6871 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5417), 
	.D(n5413), 
	.C(n5415), 
	.B(n5414), 
	.A(n5416));
   MUX4EHD U6872 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5418), 
	.D(\ram[31][8] ), 
	.C(\ram[29][8] ), 
	.B(\ram[30][8] ), 
	.A(\ram[28][8] ));
   MUX4EHD U6873 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5419), 
	.D(\ram[27][8] ), 
	.C(\ram[25][8] ), 
	.B(\ram[26][8] ), 
	.A(\ram[24][8] ));
   MUX4EHD U6874 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5420), 
	.D(\ram[23][8] ), 
	.C(\ram[21][8] ), 
	.B(\ram[22][8] ), 
	.A(\ram[20][8] ));
   MUX4EHD U6875 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5421), 
	.D(\ram[19][8] ), 
	.C(\ram[17][8] ), 
	.B(\ram[18][8] ), 
	.A(\ram[16][8] ));
   MUX4EHD U6876 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5422), 
	.D(n5418), 
	.C(n5420), 
	.B(n5419), 
	.A(n5421));
   MUX4EHD U6877 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5423), 
	.D(\ram[15][8] ), 
	.C(\ram[13][8] ), 
	.B(\ram[14][8] ), 
	.A(\ram[12][8] ));
   MUX4EHD U6878 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5424), 
	.D(\ram[11][8] ), 
	.C(\ram[9][8] ), 
	.B(\ram[10][8] ), 
	.A(\ram[8][8] ));
   MUX4EHD U6879 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5425), 
	.D(\ram[7][8] ), 
	.C(\ram[5][8] ), 
	.B(\ram[6][8] ), 
	.A(\ram[4][8] ));
   MUX4EHD U6880 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n5426), 
	.D(\ram[3][8] ), 
	.C(\ram[1][8] ), 
	.B(\ram[2][8] ), 
	.A(\ram[0][8] ));
   MUX4EHD U6881 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5427), 
	.D(n5423), 
	.C(n5425), 
	.B(n5424), 
	.A(n5426));
   MUX4EHD U6882 (.S1(n6038), 
	.S0(n7444), 
	.O(n5428), 
	.D(n5412), 
	.C(n5422), 
	.B(n5417), 
	.A(n5427));
   MUX4EHD U6883 (.S1(n6469), 
	.S0(n6470), 
	.O(N4133), 
	.D(n5365), 
	.C(n5407), 
	.B(n5386), 
	.A(n5428));
   MUX4EHD U6884 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5429), 
	.D(\ram[255][9] ), 
	.C(\ram[253][9] ), 
	.B(\ram[254][9] ), 
	.A(\ram[252][9] ));
   MUX4EHD U6885 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5430), 
	.D(\ram[251][9] ), 
	.C(\ram[249][9] ), 
	.B(\ram[250][9] ), 
	.A(\ram[248][9] ));
   MUX4EHD U6886 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5431), 
	.D(\ram[247][9] ), 
	.C(\ram[245][9] ), 
	.B(\ram[246][9] ), 
	.A(\ram[244][9] ));
   MUX4EHD U6887 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5432), 
	.D(\ram[243][9] ), 
	.C(\ram[241][9] ), 
	.B(\ram[242][9] ), 
	.A(\ram[240][9] ));
   MUX4EHD U6888 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5433), 
	.D(n5429), 
	.C(n5431), 
	.B(n5430), 
	.A(n5432));
   MUX4EHD U6889 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5434), 
	.D(\ram[239][9] ), 
	.C(\ram[237][9] ), 
	.B(\ram[238][9] ), 
	.A(\ram[236][9] ));
   MUX4EHD U6890 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5435), 
	.D(\ram[235][9] ), 
	.C(\ram[233][9] ), 
	.B(\ram[234][9] ), 
	.A(\ram[232][9] ));
   MUX4EHD U6891 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5436), 
	.D(\ram[231][9] ), 
	.C(\ram[229][9] ), 
	.B(\ram[230][9] ), 
	.A(\ram[228][9] ));
   MUX4EHD U6892 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5437), 
	.D(\ram[227][9] ), 
	.C(\ram[225][9] ), 
	.B(\ram[226][9] ), 
	.A(\ram[224][9] ));
   MUX4EHD U6893 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5438), 
	.D(n5434), 
	.C(n5436), 
	.B(n5435), 
	.A(n5437));
   MUX4EHD U6894 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5439), 
	.D(\ram[223][9] ), 
	.C(\ram[221][9] ), 
	.B(\ram[222][9] ), 
	.A(\ram[220][9] ));
   MUX4EHD U6895 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5440), 
	.D(\ram[219][9] ), 
	.C(\ram[217][9] ), 
	.B(\ram[218][9] ), 
	.A(\ram[216][9] ));
   MUX4EHD U6896 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5441), 
	.D(\ram[215][9] ), 
	.C(\ram[213][9] ), 
	.B(\ram[214][9] ), 
	.A(\ram[212][9] ));
   MUX4EHD U6897 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5442), 
	.D(\ram[211][9] ), 
	.C(\ram[209][9] ), 
	.B(\ram[210][9] ), 
	.A(\ram[208][9] ));
   MUX4EHD U6898 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5443), 
	.D(n5439), 
	.C(n5441), 
	.B(n5440), 
	.A(n5442));
   MUX4EHD U6899 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5444), 
	.D(\ram[207][9] ), 
	.C(\ram[205][9] ), 
	.B(\ram[206][9] ), 
	.A(\ram[204][9] ));
   MUX4EHD U6900 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5445), 
	.D(\ram[203][9] ), 
	.C(\ram[201][9] ), 
	.B(\ram[202][9] ), 
	.A(\ram[200][9] ));
   MUX4EHD U6901 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5446), 
	.D(\ram[199][9] ), 
	.C(\ram[197][9] ), 
	.B(\ram[198][9] ), 
	.A(\ram[196][9] ));
   MUX4EHD U6902 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5447), 
	.D(\ram[195][9] ), 
	.C(\ram[193][9] ), 
	.B(\ram[194][9] ), 
	.A(\ram[192][9] ));
   MUX4EHD U6903 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5448), 
	.D(n5444), 
	.C(n5446), 
	.B(n5445), 
	.A(n5447));
   MUX4EHD U6904 (.S1(n6038), 
	.S0(n7444), 
	.O(n5449), 
	.D(n5433), 
	.C(n5443), 
	.B(n5438), 
	.A(n5448));
   MUX4EHD U6905 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5450), 
	.D(\ram[191][9] ), 
	.C(\ram[189][9] ), 
	.B(\ram[190][9] ), 
	.A(\ram[188][9] ));
   MUX4EHD U6906 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5451), 
	.D(\ram[187][9] ), 
	.C(\ram[185][9] ), 
	.B(\ram[186][9] ), 
	.A(\ram[184][9] ));
   MUX4EHD U6907 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5452), 
	.D(\ram[183][9] ), 
	.C(\ram[181][9] ), 
	.B(\ram[182][9] ), 
	.A(\ram[180][9] ));
   MUX4EHD U6908 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5453), 
	.D(\ram[179][9] ), 
	.C(\ram[177][9] ), 
	.B(\ram[178][9] ), 
	.A(\ram[176][9] ));
   MUX4EHD U6909 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5454), 
	.D(n5450), 
	.C(n5452), 
	.B(n5451), 
	.A(n5453));
   MUX4EHD U6910 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5455), 
	.D(\ram[175][9] ), 
	.C(\ram[173][9] ), 
	.B(\ram[174][9] ), 
	.A(\ram[172][9] ));
   MUX4EHD U6911 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5456), 
	.D(\ram[171][9] ), 
	.C(\ram[169][9] ), 
	.B(\ram[170][9] ), 
	.A(\ram[168][9] ));
   MUX4EHD U6912 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5457), 
	.D(\ram[167][9] ), 
	.C(\ram[165][9] ), 
	.B(\ram[166][9] ), 
	.A(\ram[164][9] ));
   MUX4EHD U6913 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5458), 
	.D(\ram[163][9] ), 
	.C(\ram[161][9] ), 
	.B(\ram[162][9] ), 
	.A(\ram[160][9] ));
   MUX4EHD U6914 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5459), 
	.D(n5455), 
	.C(n5457), 
	.B(n5456), 
	.A(n5458));
   MUX4EHD U6915 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5460), 
	.D(\ram[159][9] ), 
	.C(\ram[157][9] ), 
	.B(\ram[158][9] ), 
	.A(\ram[156][9] ));
   MUX4EHD U6916 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5461), 
	.D(\ram[155][9] ), 
	.C(\ram[153][9] ), 
	.B(\ram[154][9] ), 
	.A(\ram[152][9] ));
   MUX4EHD U6917 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5462), 
	.D(\ram[151][9] ), 
	.C(\ram[149][9] ), 
	.B(\ram[150][9] ), 
	.A(\ram[148][9] ));
   MUX4EHD U6918 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5463), 
	.D(\ram[147][9] ), 
	.C(\ram[145][9] ), 
	.B(\ram[146][9] ), 
	.A(\ram[144][9] ));
   MUX4EHD U6919 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5464), 
	.D(n5460), 
	.C(n5462), 
	.B(n5461), 
	.A(n5463));
   MUX4EHD U6920 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5465), 
	.D(\ram[143][9] ), 
	.C(\ram[141][9] ), 
	.B(\ram[142][9] ), 
	.A(\ram[140][9] ));
   MUX4EHD U6921 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5466), 
	.D(\ram[139][9] ), 
	.C(\ram[137][9] ), 
	.B(\ram[138][9] ), 
	.A(\ram[136][9] ));
   MUX4EHD U6922 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5467), 
	.D(\ram[135][9] ), 
	.C(\ram[133][9] ), 
	.B(\ram[134][9] ), 
	.A(\ram[132][9] ));
   MUX4EHD U6923 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5468), 
	.D(\ram[131][9] ), 
	.C(\ram[129][9] ), 
	.B(\ram[130][9] ), 
	.A(\ram[128][9] ));
   MUX4EHD U6924 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5469), 
	.D(n5465), 
	.C(n5467), 
	.B(n5466), 
	.A(n5468));
   MUX4EHD U6925 (.S1(n6038), 
	.S0(n7444), 
	.O(n5470), 
	.D(n5454), 
	.C(n5464), 
	.B(n5459), 
	.A(n5469));
   MUX4EHD U6926 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5471), 
	.D(\ram[127][9] ), 
	.C(\ram[125][9] ), 
	.B(\ram[126][9] ), 
	.A(\ram[124][9] ));
   MUX4EHD U6927 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5472), 
	.D(\ram[123][9] ), 
	.C(\ram[121][9] ), 
	.B(\ram[122][9] ), 
	.A(\ram[120][9] ));
   MUX4EHD U6928 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5473), 
	.D(\ram[119][9] ), 
	.C(\ram[117][9] ), 
	.B(\ram[118][9] ), 
	.A(\ram[116][9] ));
   MUX4EHD U6929 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5474), 
	.D(\ram[115][9] ), 
	.C(\ram[113][9] ), 
	.B(\ram[114][9] ), 
	.A(\ram[112][9] ));
   MUX4EHD U6930 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5475), 
	.D(n5471), 
	.C(n5473), 
	.B(n5472), 
	.A(n5474));
   MUX4EHD U6931 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5476), 
	.D(\ram[111][9] ), 
	.C(\ram[109][9] ), 
	.B(\ram[110][9] ), 
	.A(\ram[108][9] ));
   MUX4EHD U6932 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5477), 
	.D(\ram[107][9] ), 
	.C(\ram[105][9] ), 
	.B(\ram[106][9] ), 
	.A(\ram[104][9] ));
   MUX4EHD U6933 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5478), 
	.D(\ram[103][9] ), 
	.C(\ram[101][9] ), 
	.B(\ram[102][9] ), 
	.A(\ram[100][9] ));
   MUX4EHD U6934 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5479), 
	.D(\ram[99][9] ), 
	.C(\ram[97][9] ), 
	.B(\ram[98][9] ), 
	.A(\ram[96][9] ));
   MUX4EHD U6935 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5480), 
	.D(n5476), 
	.C(n5478), 
	.B(n5477), 
	.A(n5479));
   MUX4EHD U6936 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5481), 
	.D(\ram[95][9] ), 
	.C(\ram[93][9] ), 
	.B(\ram[94][9] ), 
	.A(\ram[92][9] ));
   MUX4EHD U6937 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5482), 
	.D(\ram[91][9] ), 
	.C(\ram[89][9] ), 
	.B(\ram[90][9] ), 
	.A(\ram[88][9] ));
   MUX4EHD U6938 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5483), 
	.D(\ram[87][9] ), 
	.C(\ram[85][9] ), 
	.B(\ram[86][9] ), 
	.A(\ram[84][9] ));
   MUX4EHD U6939 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5484), 
	.D(\ram[83][9] ), 
	.C(\ram[81][9] ), 
	.B(\ram[82][9] ), 
	.A(\ram[80][9] ));
   MUX4EHD U6940 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5485), 
	.D(n5481), 
	.C(n5483), 
	.B(n5482), 
	.A(n5484));
   MUX4EHD U6941 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5486), 
	.D(\ram[79][9] ), 
	.C(\ram[77][9] ), 
	.B(\ram[78][9] ), 
	.A(\ram[76][9] ));
   MUX4EHD U6942 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5487), 
	.D(\ram[75][9] ), 
	.C(\ram[73][9] ), 
	.B(\ram[74][9] ), 
	.A(\ram[72][9] ));
   MUX4EHD U6943 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5488), 
	.D(\ram[71][9] ), 
	.C(\ram[69][9] ), 
	.B(\ram[70][9] ), 
	.A(\ram[68][9] ));
   MUX4EHD U6944 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5489), 
	.D(\ram[67][9] ), 
	.C(\ram[65][9] ), 
	.B(\ram[66][9] ), 
	.A(\ram[64][9] ));
   MUX4EHD U6945 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5490), 
	.D(n5486), 
	.C(n5488), 
	.B(n5487), 
	.A(n5489));
   MUX4EHD U6946 (.S1(n6038), 
	.S0(n7444), 
	.O(n5491), 
	.D(n5475), 
	.C(n5485), 
	.B(n5480), 
	.A(n5490));
   MUX4EHD U6947 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5492), 
	.D(\ram[63][9] ), 
	.C(\ram[61][9] ), 
	.B(\ram[62][9] ), 
	.A(\ram[60][9] ));
   MUX4EHD U6948 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5493), 
	.D(\ram[59][9] ), 
	.C(\ram[57][9] ), 
	.B(\ram[58][9] ), 
	.A(\ram[56][9] ));
   MUX4EHD U6949 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5494), 
	.D(\ram[55][9] ), 
	.C(\ram[53][9] ), 
	.B(\ram[54][9] ), 
	.A(\ram[52][9] ));
   MUX4EHD U6950 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5495), 
	.D(\ram[51][9] ), 
	.C(\ram[49][9] ), 
	.B(\ram[50][9] ), 
	.A(\ram[48][9] ));
   MUX4EHD U6951 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5496), 
	.D(n5492), 
	.C(n5494), 
	.B(n5493), 
	.A(n5495));
   MUX4EHD U6952 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5497), 
	.D(\ram[47][9] ), 
	.C(\ram[45][9] ), 
	.B(\ram[46][9] ), 
	.A(\ram[44][9] ));
   MUX4EHD U6953 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5498), 
	.D(\ram[43][9] ), 
	.C(\ram[41][9] ), 
	.B(\ram[42][9] ), 
	.A(\ram[40][9] ));
   MUX4EHD U6954 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5499), 
	.D(\ram[39][9] ), 
	.C(\ram[37][9] ), 
	.B(\ram[38][9] ), 
	.A(\ram[36][9] ));
   MUX4EHD U6955 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5500), 
	.D(\ram[35][9] ), 
	.C(\ram[33][9] ), 
	.B(\ram[34][9] ), 
	.A(\ram[32][9] ));
   MUX4EHD U6956 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5501), 
	.D(n5497), 
	.C(n5499), 
	.B(n5498), 
	.A(n5500));
   MUX4EHD U6957 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5502), 
	.D(\ram[31][9] ), 
	.C(\ram[29][9] ), 
	.B(\ram[30][9] ), 
	.A(\ram[28][9] ));
   MUX4EHD U6958 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5503), 
	.D(\ram[27][9] ), 
	.C(\ram[25][9] ), 
	.B(\ram[26][9] ), 
	.A(\ram[24][9] ));
   MUX4EHD U6959 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5504), 
	.D(\ram[23][9] ), 
	.C(\ram[21][9] ), 
	.B(\ram[22][9] ), 
	.A(\ram[20][9] ));
   MUX4EHD U6960 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5505), 
	.D(\ram[19][9] ), 
	.C(\ram[17][9] ), 
	.B(\ram[18][9] ), 
	.A(\ram[16][9] ));
   MUX4EHD U6961 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5506), 
	.D(n5502), 
	.C(n5504), 
	.B(n5503), 
	.A(n5505));
   MUX4EHD U6962 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5507), 
	.D(\ram[15][9] ), 
	.C(\ram[13][9] ), 
	.B(\ram[14][9] ), 
	.A(\ram[12][9] ));
   MUX4EHD U6963 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5508), 
	.D(\ram[11][9] ), 
	.C(\ram[9][9] ), 
	.B(\ram[10][9] ), 
	.A(\ram[8][9] ));
   MUX4EHD U6964 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5509), 
	.D(\ram[7][9] ), 
	.C(\ram[5][9] ), 
	.B(\ram[6][9] ), 
	.A(\ram[4][9] ));
   MUX4EHD U6965 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5510), 
	.D(\ram[3][9] ), 
	.C(\ram[1][9] ), 
	.B(\ram[2][9] ), 
	.A(\ram[0][9] ));
   MUX4EHD U6966 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5511), 
	.D(n5507), 
	.C(n5509), 
	.B(n5508), 
	.A(n5510));
   MUX4EHD U6967 (.S1(n6038), 
	.S0(n7444), 
	.O(n5512), 
	.D(n5496), 
	.C(n5506), 
	.B(n5501), 
	.A(n5511));
   MUX4EHD U6968 (.S1(n6469), 
	.S0(n6470), 
	.O(N4132), 
	.D(n5449), 
	.C(n5491), 
	.B(n5470), 
	.A(n5512));
   MUX4EHD U6969 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5513), 
	.D(\ram[255][10] ), 
	.C(\ram[253][10] ), 
	.B(\ram[254][10] ), 
	.A(\ram[252][10] ));
   MUX4EHD U6970 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5514), 
	.D(\ram[251][10] ), 
	.C(\ram[249][10] ), 
	.B(\ram[250][10] ), 
	.A(\ram[248][10] ));
   MUX4EHD U6971 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5515), 
	.D(\ram[247][10] ), 
	.C(\ram[245][10] ), 
	.B(\ram[246][10] ), 
	.A(\ram[244][10] ));
   MUX4EHD U6972 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5516), 
	.D(\ram[243][10] ), 
	.C(\ram[241][10] ), 
	.B(\ram[242][10] ), 
	.A(\ram[240][10] ));
   MUX4EHD U6973 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5517), 
	.D(n5513), 
	.C(n5515), 
	.B(n5514), 
	.A(n5516));
   MUX4EHD U6974 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5518), 
	.D(\ram[239][10] ), 
	.C(\ram[237][10] ), 
	.B(\ram[238][10] ), 
	.A(\ram[236][10] ));
   MUX4EHD U6975 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5519), 
	.D(\ram[235][10] ), 
	.C(\ram[233][10] ), 
	.B(\ram[234][10] ), 
	.A(\ram[232][10] ));
   MUX4EHD U6976 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5520), 
	.D(\ram[231][10] ), 
	.C(\ram[229][10] ), 
	.B(\ram[230][10] ), 
	.A(\ram[228][10] ));
   MUX4EHD U6977 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5521), 
	.D(\ram[227][10] ), 
	.C(\ram[225][10] ), 
	.B(\ram[226][10] ), 
	.A(\ram[224][10] ));
   MUX4EHD U6978 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5522), 
	.D(n5518), 
	.C(n5520), 
	.B(n5519), 
	.A(n5521));
   MUX4EHD U6979 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5523), 
	.D(\ram[223][10] ), 
	.C(\ram[221][10] ), 
	.B(\ram[222][10] ), 
	.A(\ram[220][10] ));
   MUX4EHD U6980 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5524), 
	.D(\ram[219][10] ), 
	.C(\ram[217][10] ), 
	.B(\ram[218][10] ), 
	.A(\ram[216][10] ));
   MUX4EHD U6981 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5525), 
	.D(\ram[215][10] ), 
	.C(\ram[213][10] ), 
	.B(\ram[214][10] ), 
	.A(\ram[212][10] ));
   MUX4EHD U6982 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5526), 
	.D(\ram[211][10] ), 
	.C(\ram[209][10] ), 
	.B(\ram[210][10] ), 
	.A(\ram[208][10] ));
   MUX4EHD U6983 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5527), 
	.D(n5523), 
	.C(n5525), 
	.B(n5524), 
	.A(n5526));
   MUX4EHD U6984 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5528), 
	.D(\ram[207][10] ), 
	.C(\ram[205][10] ), 
	.B(\ram[206][10] ), 
	.A(\ram[204][10] ));
   MUX4EHD U6985 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5529), 
	.D(\ram[203][10] ), 
	.C(\ram[201][10] ), 
	.B(\ram[202][10] ), 
	.A(\ram[200][10] ));
   MUX4EHD U6986 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5530), 
	.D(\ram[199][10] ), 
	.C(\ram[197][10] ), 
	.B(\ram[198][10] ), 
	.A(\ram[196][10] ));
   MUX4EHD U6987 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5531), 
	.D(\ram[195][10] ), 
	.C(\ram[193][10] ), 
	.B(\ram[194][10] ), 
	.A(\ram[192][10] ));
   MUX4EHD U6988 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5532), 
	.D(n5528), 
	.C(n5530), 
	.B(n5529), 
	.A(n5531));
   MUX4EHD U6989 (.S1(n6038), 
	.S0(n7444), 
	.O(n5533), 
	.D(n5517), 
	.C(n5527), 
	.B(n5522), 
	.A(n5532));
   MUX4EHD U6990 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5534), 
	.D(\ram[191][10] ), 
	.C(\ram[189][10] ), 
	.B(\ram[190][10] ), 
	.A(\ram[188][10] ));
   MUX4EHD U6991 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5535), 
	.D(\ram[187][10] ), 
	.C(\ram[185][10] ), 
	.B(\ram[186][10] ), 
	.A(\ram[184][10] ));
   MUX4EHD U6992 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5536), 
	.D(\ram[183][10] ), 
	.C(\ram[181][10] ), 
	.B(\ram[182][10] ), 
	.A(\ram[180][10] ));
   MUX4EHD U6993 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5537), 
	.D(\ram[179][10] ), 
	.C(\ram[177][10] ), 
	.B(\ram[178][10] ), 
	.A(\ram[176][10] ));
   MUX4EHD U6994 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5538), 
	.D(n5534), 
	.C(n5536), 
	.B(n5535), 
	.A(n5537));
   MUX4EHD U6995 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5539), 
	.D(\ram[175][10] ), 
	.C(\ram[173][10] ), 
	.B(\ram[174][10] ), 
	.A(\ram[172][10] ));
   MUX4EHD U6996 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5540), 
	.D(\ram[171][10] ), 
	.C(\ram[169][10] ), 
	.B(\ram[170][10] ), 
	.A(\ram[168][10] ));
   MUX4EHD U6997 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5541), 
	.D(\ram[167][10] ), 
	.C(\ram[165][10] ), 
	.B(\ram[166][10] ), 
	.A(\ram[164][10] ));
   MUX4EHD U6998 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5542), 
	.D(\ram[163][10] ), 
	.C(\ram[161][10] ), 
	.B(\ram[162][10] ), 
	.A(\ram[160][10] ));
   MUX4EHD U6999 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5543), 
	.D(n5539), 
	.C(n5541), 
	.B(n5540), 
	.A(n5542));
   MUX4EHD U7000 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5544), 
	.D(\ram[159][10] ), 
	.C(\ram[157][10] ), 
	.B(\ram[158][10] ), 
	.A(\ram[156][10] ));
   MUX4EHD U7001 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5545), 
	.D(\ram[155][10] ), 
	.C(\ram[153][10] ), 
	.B(\ram[154][10] ), 
	.A(\ram[152][10] ));
   MUX4EHD U7002 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5546), 
	.D(\ram[151][10] ), 
	.C(\ram[149][10] ), 
	.B(\ram[150][10] ), 
	.A(\ram[148][10] ));
   MUX4EHD U7003 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5547), 
	.D(\ram[147][10] ), 
	.C(\ram[145][10] ), 
	.B(\ram[146][10] ), 
	.A(\ram[144][10] ));
   MUX4EHD U7004 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5548), 
	.D(n5544), 
	.C(n5546), 
	.B(n5545), 
	.A(n5547));
   MUX4EHD U7005 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5549), 
	.D(\ram[143][10] ), 
	.C(\ram[141][10] ), 
	.B(\ram[142][10] ), 
	.A(\ram[140][10] ));
   MUX4EHD U7006 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5550), 
	.D(\ram[139][10] ), 
	.C(\ram[137][10] ), 
	.B(\ram[138][10] ), 
	.A(\ram[136][10] ));
   MUX4EHD U7007 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5551), 
	.D(\ram[135][10] ), 
	.C(\ram[133][10] ), 
	.B(\ram[134][10] ), 
	.A(\ram[132][10] ));
   MUX4EHD U7008 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5552), 
	.D(\ram[131][10] ), 
	.C(\ram[129][10] ), 
	.B(\ram[130][10] ), 
	.A(\ram[128][10] ));
   MUX4EHD U7009 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5553), 
	.D(n5549), 
	.C(n5551), 
	.B(n5550), 
	.A(n5552));
   MUX4EHD U7010 (.S1(n6038), 
	.S0(n7444), 
	.O(n5554), 
	.D(n5538), 
	.C(n5548), 
	.B(n5543), 
	.A(n5553));
   MUX4EHD U7011 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5555), 
	.D(\ram[127][10] ), 
	.C(\ram[125][10] ), 
	.B(\ram[126][10] ), 
	.A(\ram[124][10] ));
   MUX4EHD U7012 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5556), 
	.D(\ram[123][10] ), 
	.C(\ram[121][10] ), 
	.B(\ram[122][10] ), 
	.A(\ram[120][10] ));
   MUX4EHD U7013 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5557), 
	.D(\ram[119][10] ), 
	.C(\ram[117][10] ), 
	.B(\ram[118][10] ), 
	.A(\ram[116][10] ));
   MUX4EHD U7014 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5558), 
	.D(\ram[115][10] ), 
	.C(\ram[113][10] ), 
	.B(\ram[114][10] ), 
	.A(\ram[112][10] ));
   MUX4EHD U7015 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5559), 
	.D(n5555), 
	.C(n5557), 
	.B(n5556), 
	.A(n5558));
   MUX4EHD U7016 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5560), 
	.D(\ram[111][10] ), 
	.C(\ram[109][10] ), 
	.B(\ram[110][10] ), 
	.A(\ram[108][10] ));
   MUX4EHD U7017 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5561), 
	.D(\ram[107][10] ), 
	.C(\ram[105][10] ), 
	.B(\ram[106][10] ), 
	.A(\ram[104][10] ));
   MUX4EHD U7018 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5562), 
	.D(\ram[103][10] ), 
	.C(\ram[101][10] ), 
	.B(\ram[102][10] ), 
	.A(\ram[100][10] ));
   MUX4EHD U7019 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5563), 
	.D(\ram[99][10] ), 
	.C(\ram[97][10] ), 
	.B(\ram[98][10] ), 
	.A(\ram[96][10] ));
   MUX4EHD U7020 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5564), 
	.D(n5560), 
	.C(n5562), 
	.B(n5561), 
	.A(n5563));
   MUX4EHD U7021 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5565), 
	.D(\ram[95][10] ), 
	.C(\ram[93][10] ), 
	.B(\ram[94][10] ), 
	.A(\ram[92][10] ));
   MUX4EHD U7022 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5566), 
	.D(\ram[91][10] ), 
	.C(\ram[89][10] ), 
	.B(\ram[90][10] ), 
	.A(\ram[88][10] ));
   MUX4EHD U7023 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5567), 
	.D(\ram[87][10] ), 
	.C(\ram[85][10] ), 
	.B(\ram[86][10] ), 
	.A(\ram[84][10] ));
   MUX4EHD U7024 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5568), 
	.D(\ram[83][10] ), 
	.C(\ram[81][10] ), 
	.B(\ram[82][10] ), 
	.A(\ram[80][10] ));
   MUX4EHD U7025 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5569), 
	.D(n5565), 
	.C(n5567), 
	.B(n5566), 
	.A(n5568));
   MUX4EHD U7026 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5570), 
	.D(\ram[79][10] ), 
	.C(\ram[77][10] ), 
	.B(\ram[78][10] ), 
	.A(\ram[76][10] ));
   MUX4EHD U7027 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5571), 
	.D(\ram[75][10] ), 
	.C(\ram[73][10] ), 
	.B(\ram[74][10] ), 
	.A(\ram[72][10] ));
   MUX4EHD U7028 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5572), 
	.D(\ram[71][10] ), 
	.C(\ram[69][10] ), 
	.B(\ram[70][10] ), 
	.A(\ram[68][10] ));
   MUX4EHD U7029 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5573), 
	.D(\ram[67][10] ), 
	.C(\ram[65][10] ), 
	.B(\ram[66][10] ), 
	.A(\ram[64][10] ));
   MUX4EHD U7030 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5574), 
	.D(n5570), 
	.C(n5572), 
	.B(n5571), 
	.A(n5573));
   MUX4EHD U7031 (.S1(n6038), 
	.S0(n7444), 
	.O(n5575), 
	.D(n5559), 
	.C(n5569), 
	.B(n5564), 
	.A(n5574));
   MUX4EHD U7032 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5576), 
	.D(\ram[63][10] ), 
	.C(\ram[61][10] ), 
	.B(\ram[62][10] ), 
	.A(\ram[60][10] ));
   MUX4EHD U7033 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5577), 
	.D(\ram[59][10] ), 
	.C(\ram[57][10] ), 
	.B(\ram[58][10] ), 
	.A(\ram[56][10] ));
   MUX4EHD U7034 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5578), 
	.D(\ram[55][10] ), 
	.C(\ram[53][10] ), 
	.B(\ram[54][10] ), 
	.A(\ram[52][10] ));
   MUX4EHD U7035 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5579), 
	.D(\ram[51][10] ), 
	.C(\ram[49][10] ), 
	.B(\ram[50][10] ), 
	.A(\ram[48][10] ));
   MUX4EHD U7036 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5580), 
	.D(n5576), 
	.C(n5578), 
	.B(n5577), 
	.A(n5579));
   MUX4EHD U7037 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5581), 
	.D(\ram[47][10] ), 
	.C(\ram[45][10] ), 
	.B(\ram[46][10] ), 
	.A(\ram[44][10] ));
   MUX4EHD U7038 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5582), 
	.D(\ram[43][10] ), 
	.C(\ram[41][10] ), 
	.B(\ram[42][10] ), 
	.A(\ram[40][10] ));
   MUX4EHD U7039 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5583), 
	.D(\ram[39][10] ), 
	.C(\ram[37][10] ), 
	.B(\ram[38][10] ), 
	.A(\ram[36][10] ));
   MUX4EHD U7040 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5584), 
	.D(\ram[35][10] ), 
	.C(\ram[33][10] ), 
	.B(\ram[34][10] ), 
	.A(\ram[32][10] ));
   MUX4EHD U7041 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5585), 
	.D(n5581), 
	.C(n5583), 
	.B(n5582), 
	.A(n5584));
   MUX4EHD U7042 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5586), 
	.D(\ram[31][10] ), 
	.C(\ram[29][10] ), 
	.B(\ram[30][10] ), 
	.A(\ram[28][10] ));
   MUX4EHD U7043 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5587), 
	.D(\ram[27][10] ), 
	.C(\ram[25][10] ), 
	.B(\ram[26][10] ), 
	.A(\ram[24][10] ));
   MUX4EHD U7044 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5588), 
	.D(\ram[23][10] ), 
	.C(\ram[21][10] ), 
	.B(\ram[22][10] ), 
	.A(\ram[20][10] ));
   MUX4EHD U7045 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5589), 
	.D(\ram[19][10] ), 
	.C(\ram[17][10] ), 
	.B(\ram[18][10] ), 
	.A(\ram[16][10] ));
   MUX4EHD U7046 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5590), 
	.D(n5586), 
	.C(n5588), 
	.B(n5587), 
	.A(n5589));
   MUX4EHD U7047 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5591), 
	.D(\ram[15][10] ), 
	.C(\ram[13][10] ), 
	.B(\ram[14][10] ), 
	.A(\ram[12][10] ));
   MUX4EHD U7048 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5592), 
	.D(\ram[11][10] ), 
	.C(\ram[9][10] ), 
	.B(\ram[10][10] ), 
	.A(\ram[8][10] ));
   MUX4EHD U7049 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5593), 
	.D(\ram[7][10] ), 
	.C(\ram[5][10] ), 
	.B(\ram[6][10] ), 
	.A(\ram[4][10] ));
   MUX4EHD U7050 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5594), 
	.D(\ram[3][10] ), 
	.C(\ram[1][10] ), 
	.B(\ram[2][10] ), 
	.A(\ram[0][10] ));
   MUX4EHD U7051 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5595), 
	.D(n5591), 
	.C(n5593), 
	.B(n5592), 
	.A(n5594));
   MUX4EHD U7052 (.S1(n6038), 
	.S0(n7444), 
	.O(n5596), 
	.D(n5580), 
	.C(n5590), 
	.B(n5585), 
	.A(n5595));
   MUX4EHD U7053 (.S1(n6469), 
	.S0(n6470), 
	.O(N4131), 
	.D(n5533), 
	.C(n5575), 
	.B(n5554), 
	.A(n5596));
   MUX4EHD U7054 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5597), 
	.D(\ram[255][11] ), 
	.C(\ram[253][11] ), 
	.B(\ram[254][11] ), 
	.A(\ram[252][11] ));
   MUX4EHD U7055 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5598), 
	.D(\ram[251][11] ), 
	.C(\ram[249][11] ), 
	.B(\ram[250][11] ), 
	.A(\ram[248][11] ));
   MUX4EHD U7056 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5599), 
	.D(\ram[247][11] ), 
	.C(\ram[245][11] ), 
	.B(\ram[246][11] ), 
	.A(\ram[244][11] ));
   MUX4EHD U7057 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5600), 
	.D(\ram[243][11] ), 
	.C(\ram[241][11] ), 
	.B(\ram[242][11] ), 
	.A(\ram[240][11] ));
   MUX4EHD U7058 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5601), 
	.D(n5597), 
	.C(n5599), 
	.B(n5598), 
	.A(n5600));
   MUX4EHD U7059 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5602), 
	.D(\ram[239][11] ), 
	.C(\ram[237][11] ), 
	.B(\ram[238][11] ), 
	.A(\ram[236][11] ));
   MUX4EHD U7060 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5603), 
	.D(\ram[235][11] ), 
	.C(\ram[233][11] ), 
	.B(\ram[234][11] ), 
	.A(\ram[232][11] ));
   MUX4EHD U7061 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5604), 
	.D(\ram[231][11] ), 
	.C(\ram[229][11] ), 
	.B(\ram[230][11] ), 
	.A(\ram[228][11] ));
   MUX4EHD U7062 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5605), 
	.D(\ram[227][11] ), 
	.C(\ram[225][11] ), 
	.B(\ram[226][11] ), 
	.A(\ram[224][11] ));
   MUX4EHD U7063 (.S1(n6136), 
	.S0(n7442), 
	.O(n5606), 
	.D(n5602), 
	.C(n5604), 
	.B(n5603), 
	.A(n5605));
   MUX4EHD U7064 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5607), 
	.D(\ram[223][11] ), 
	.C(\ram[221][11] ), 
	.B(\ram[222][11] ), 
	.A(\ram[220][11] ));
   MUX4EHD U7065 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5608), 
	.D(\ram[219][11] ), 
	.C(\ram[217][11] ), 
	.B(\ram[218][11] ), 
	.A(\ram[216][11] ));
   MUX4EHD U7066 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5609), 
	.D(\ram[215][11] ), 
	.C(\ram[213][11] ), 
	.B(\ram[214][11] ), 
	.A(\ram[212][11] ));
   MUX4EHD U7067 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5610), 
	.D(\ram[211][11] ), 
	.C(\ram[209][11] ), 
	.B(\ram[210][11] ), 
	.A(\ram[208][11] ));
   MUX4EHD U7068 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5611), 
	.D(n5607), 
	.C(n5609), 
	.B(n5608), 
	.A(n5610));
   MUX4EHD U7069 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5612), 
	.D(\ram[207][11] ), 
	.C(\ram[205][11] ), 
	.B(\ram[206][11] ), 
	.A(\ram[204][11] ));
   MUX4EHD U7070 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5613), 
	.D(\ram[203][11] ), 
	.C(\ram[201][11] ), 
	.B(\ram[202][11] ), 
	.A(\ram[200][11] ));
   MUX4EHD U7071 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5614), 
	.D(\ram[199][11] ), 
	.C(\ram[197][11] ), 
	.B(\ram[198][11] ), 
	.A(\ram[196][11] ));
   MUX4EHD U7072 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5615), 
	.D(\ram[195][11] ), 
	.C(\ram[193][11] ), 
	.B(\ram[194][11] ), 
	.A(\ram[192][11] ));
   MUX4EHD U7073 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5616), 
	.D(n5612), 
	.C(n5614), 
	.B(n5613), 
	.A(n5615));
   MUX4EHD U7074 (.S1(n6038), 
	.S0(n7444), 
	.O(n5617), 
	.D(n5601), 
	.C(n5611), 
	.B(n5606), 
	.A(n5616));
   MUX4EHD U7075 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5618), 
	.D(\ram[191][11] ), 
	.C(\ram[189][11] ), 
	.B(\ram[190][11] ), 
	.A(\ram[188][11] ));
   MUX4EHD U7076 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5619), 
	.D(\ram[187][11] ), 
	.C(\ram[185][11] ), 
	.B(\ram[186][11] ), 
	.A(\ram[184][11] ));
   MUX4EHD U7077 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5620), 
	.D(\ram[183][11] ), 
	.C(\ram[181][11] ), 
	.B(\ram[182][11] ), 
	.A(\ram[180][11] ));
   MUX4EHD U7078 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5621), 
	.D(\ram[179][11] ), 
	.C(\ram[177][11] ), 
	.B(\ram[178][11] ), 
	.A(\ram[176][11] ));
   MUX4EHD U7079 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5622), 
	.D(n5618), 
	.C(n5620), 
	.B(n5619), 
	.A(n5621));
   MUX4EHD U7080 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5623), 
	.D(\ram[175][11] ), 
	.C(\ram[173][11] ), 
	.B(\ram[174][11] ), 
	.A(\ram[172][11] ));
   MUX4EHD U7081 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5624), 
	.D(\ram[171][11] ), 
	.C(\ram[169][11] ), 
	.B(\ram[170][11] ), 
	.A(\ram[168][11] ));
   MUX4EHD U7082 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5625), 
	.D(\ram[167][11] ), 
	.C(\ram[165][11] ), 
	.B(\ram[166][11] ), 
	.A(\ram[164][11] ));
   MUX4EHD U7083 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5626), 
	.D(\ram[163][11] ), 
	.C(\ram[161][11] ), 
	.B(\ram[162][11] ), 
	.A(\ram[160][11] ));
   MUX4EHD U7084 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5627), 
	.D(n5623), 
	.C(n5625), 
	.B(n5624), 
	.A(n5626));
   MUX4EHD U7085 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5628), 
	.D(\ram[159][11] ), 
	.C(\ram[157][11] ), 
	.B(\ram[158][11] ), 
	.A(\ram[156][11] ));
   MUX4EHD U7086 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5629), 
	.D(\ram[155][11] ), 
	.C(\ram[153][11] ), 
	.B(\ram[154][11] ), 
	.A(\ram[152][11] ));
   MUX4EHD U7087 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5630), 
	.D(\ram[151][11] ), 
	.C(\ram[149][11] ), 
	.B(\ram[150][11] ), 
	.A(\ram[148][11] ));
   MUX4EHD U7088 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5631), 
	.D(\ram[147][11] ), 
	.C(\ram[145][11] ), 
	.B(\ram[146][11] ), 
	.A(\ram[144][11] ));
   MUX4EHD U7089 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5632), 
	.D(n5628), 
	.C(n5630), 
	.B(n5629), 
	.A(n5631));
   MUX4EHD U7090 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5633), 
	.D(\ram[143][11] ), 
	.C(\ram[141][11] ), 
	.B(\ram[142][11] ), 
	.A(\ram[140][11] ));
   MUX4EHD U7091 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5634), 
	.D(\ram[139][11] ), 
	.C(\ram[137][11] ), 
	.B(\ram[138][11] ), 
	.A(\ram[136][11] ));
   MUX4EHD U7092 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5635), 
	.D(\ram[135][11] ), 
	.C(\ram[133][11] ), 
	.B(\ram[134][11] ), 
	.A(\ram[132][11] ));
   MUX4EHD U7093 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5636), 
	.D(\ram[131][11] ), 
	.C(\ram[129][11] ), 
	.B(\ram[130][11] ), 
	.A(\ram[128][11] ));
   MUX4EHD U7094 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5637), 
	.D(n5633), 
	.C(n5635), 
	.B(n5634), 
	.A(n5636));
   MUX4EHD U7095 (.S1(n6038), 
	.S0(n7444), 
	.O(n5638), 
	.D(n5622), 
	.C(n5632), 
	.B(n5627), 
	.A(n5637));
   MUX4EHD U7096 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5639), 
	.D(\ram[127][11] ), 
	.C(\ram[125][11] ), 
	.B(\ram[126][11] ), 
	.A(\ram[124][11] ));
   MUX4EHD U7097 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5640), 
	.D(\ram[123][11] ), 
	.C(\ram[121][11] ), 
	.B(\ram[122][11] ), 
	.A(\ram[120][11] ));
   MUX4EHD U7098 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5641), 
	.D(\ram[119][11] ), 
	.C(\ram[117][11] ), 
	.B(\ram[118][11] ), 
	.A(\ram[116][11] ));
   MUX4EHD U7099 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5642), 
	.D(\ram[115][11] ), 
	.C(\ram[113][11] ), 
	.B(\ram[114][11] ), 
	.A(\ram[112][11] ));
   MUX4EHD U7100 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5643), 
	.D(n5639), 
	.C(n5641), 
	.B(n5640), 
	.A(n5642));
   MUX4EHD U7101 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5644), 
	.D(\ram[111][11] ), 
	.C(\ram[109][11] ), 
	.B(\ram[110][11] ), 
	.A(\ram[108][11] ));
   MUX4EHD U7102 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5645), 
	.D(\ram[107][11] ), 
	.C(\ram[105][11] ), 
	.B(\ram[106][11] ), 
	.A(\ram[104][11] ));
   MUX4EHD U7103 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5646), 
	.D(\ram[103][11] ), 
	.C(\ram[101][11] ), 
	.B(\ram[102][11] ), 
	.A(\ram[100][11] ));
   MUX4EHD U7104 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5647), 
	.D(\ram[99][11] ), 
	.C(\ram[97][11] ), 
	.B(\ram[98][11] ), 
	.A(\ram[96][11] ));
   MUX4EHD U7105 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5648), 
	.D(n5644), 
	.C(n5646), 
	.B(n5645), 
	.A(n5647));
   MUX4EHD U7106 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5649), 
	.D(\ram[95][11] ), 
	.C(\ram[93][11] ), 
	.B(\ram[94][11] ), 
	.A(\ram[92][11] ));
   MUX4EHD U7107 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5650), 
	.D(\ram[91][11] ), 
	.C(\ram[89][11] ), 
	.B(\ram[90][11] ), 
	.A(\ram[88][11] ));
   MUX4EHD U7108 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5651), 
	.D(\ram[87][11] ), 
	.C(\ram[85][11] ), 
	.B(\ram[86][11] ), 
	.A(\ram[84][11] ));
   MUX4EHD U7109 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5652), 
	.D(\ram[83][11] ), 
	.C(\ram[81][11] ), 
	.B(\ram[82][11] ), 
	.A(\ram[80][11] ));
   MUX4EHD U7110 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5653), 
	.D(n5649), 
	.C(n5651), 
	.B(n5650), 
	.A(n5652));
   MUX4EHD U7111 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5654), 
	.D(\ram[79][11] ), 
	.C(\ram[77][11] ), 
	.B(\ram[78][11] ), 
	.A(\ram[76][11] ));
   MUX4EHD U7112 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5655), 
	.D(\ram[75][11] ), 
	.C(\ram[73][11] ), 
	.B(\ram[74][11] ), 
	.A(\ram[72][11] ));
   MUX4EHD U7113 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5656), 
	.D(\ram[71][11] ), 
	.C(\ram[69][11] ), 
	.B(\ram[70][11] ), 
	.A(\ram[68][11] ));
   MUX4EHD U7114 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5657), 
	.D(\ram[67][11] ), 
	.C(\ram[65][11] ), 
	.B(\ram[66][11] ), 
	.A(\ram[64][11] ));
   MUX4EHD U7115 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5658), 
	.D(n5654), 
	.C(n5656), 
	.B(n5655), 
	.A(n5657));
   MUX4EHD U7116 (.S1(n6038), 
	.S0(n7444), 
	.O(n5659), 
	.D(n5643), 
	.C(n5653), 
	.B(n5648), 
	.A(n5658));
   MUX4EHD U7117 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5660), 
	.D(\ram[63][11] ), 
	.C(\ram[61][11] ), 
	.B(\ram[62][11] ), 
	.A(\ram[60][11] ));
   MUX4EHD U7118 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5661), 
	.D(\ram[59][11] ), 
	.C(\ram[57][11] ), 
	.B(\ram[58][11] ), 
	.A(\ram[56][11] ));
   MUX4EHD U7119 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5662), 
	.D(\ram[55][11] ), 
	.C(\ram[53][11] ), 
	.B(\ram[54][11] ), 
	.A(\ram[52][11] ));
   MUX4EHD U7120 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5663), 
	.D(\ram[51][11] ), 
	.C(\ram[49][11] ), 
	.B(\ram[50][11] ), 
	.A(\ram[48][11] ));
   MUX4EHD U7121 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5664), 
	.D(n5660), 
	.C(n5662), 
	.B(n5661), 
	.A(n5663));
   MUX4EHD U7122 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5665), 
	.D(\ram[47][11] ), 
	.C(\ram[45][11] ), 
	.B(\ram[46][11] ), 
	.A(\ram[44][11] ));
   MUX4EHD U7123 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5666), 
	.D(\ram[43][11] ), 
	.C(\ram[41][11] ), 
	.B(\ram[42][11] ), 
	.A(\ram[40][11] ));
   MUX4EHD U7124 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5667), 
	.D(\ram[39][11] ), 
	.C(\ram[37][11] ), 
	.B(\ram[38][11] ), 
	.A(\ram[36][11] ));
   MUX4EHD U7125 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5668), 
	.D(\ram[35][11] ), 
	.C(\ram[33][11] ), 
	.B(\ram[34][11] ), 
	.A(\ram[32][11] ));
   MUX4EHD U7126 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5669), 
	.D(n5665), 
	.C(n5667), 
	.B(n5666), 
	.A(n5668));
   MUX4EHD U7127 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5670), 
	.D(\ram[31][11] ), 
	.C(\ram[29][11] ), 
	.B(\ram[30][11] ), 
	.A(\ram[28][11] ));
   MUX4EHD U7128 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5671), 
	.D(\ram[27][11] ), 
	.C(\ram[25][11] ), 
	.B(\ram[26][11] ), 
	.A(\ram[24][11] ));
   MUX4EHD U7129 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5672), 
	.D(\ram[23][11] ), 
	.C(\ram[21][11] ), 
	.B(\ram[22][11] ), 
	.A(\ram[20][11] ));
   MUX4EHD U7130 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5673), 
	.D(\ram[19][11] ), 
	.C(\ram[17][11] ), 
	.B(\ram[18][11] ), 
	.A(\ram[16][11] ));
   MUX4EHD U7131 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5674), 
	.D(n5670), 
	.C(n5672), 
	.B(n5671), 
	.A(n5673));
   MUX4EHD U7132 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5675), 
	.D(\ram[15][11] ), 
	.C(\ram[13][11] ), 
	.B(\ram[14][11] ), 
	.A(\ram[12][11] ));
   MUX4EHD U7133 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5676), 
	.D(\ram[11][11] ), 
	.C(\ram[9][11] ), 
	.B(\ram[10][11] ), 
	.A(\ram[8][11] ));
   MUX4EHD U7134 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5677), 
	.D(\ram[7][11] ), 
	.C(\ram[5][11] ), 
	.B(\ram[6][11] ), 
	.A(\ram[4][11] ));
   MUX4EHD U7135 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5678), 
	.D(\ram[3][11] ), 
	.C(\ram[1][11] ), 
	.B(\ram[2][11] ), 
	.A(\ram[0][11] ));
   MUX4EHD U7136 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5679), 
	.D(n5675), 
	.C(n5677), 
	.B(n5676), 
	.A(n5678));
   MUX4EHD U7137 (.S1(n6038), 
	.S0(n7444), 
	.O(n5680), 
	.D(n5664), 
	.C(n5674), 
	.B(n5669), 
	.A(n5679));
   MUX4EHD U7138 (.S1(n6469), 
	.S0(n6470), 
	.O(N4130), 
	.D(n5617), 
	.C(n5659), 
	.B(n5638), 
	.A(n5680));
   MUX4EHD U7139 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5681), 
	.D(\ram[255][12] ), 
	.C(\ram[253][12] ), 
	.B(\ram[254][12] ), 
	.A(\ram[252][12] ));
   MUX4EHD U7140 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5682), 
	.D(\ram[251][12] ), 
	.C(\ram[249][12] ), 
	.B(\ram[250][12] ), 
	.A(\ram[248][12] ));
   MUX4EHD U7141 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5683), 
	.D(\ram[247][12] ), 
	.C(\ram[245][12] ), 
	.B(\ram[246][12] ), 
	.A(\ram[244][12] ));
   MUX4EHD U7142 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5684), 
	.D(\ram[243][12] ), 
	.C(\ram[241][12] ), 
	.B(\ram[242][12] ), 
	.A(\ram[240][12] ));
   MUX4EHD U7143 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5685), 
	.D(n5681), 
	.C(n5683), 
	.B(n5682), 
	.A(n5684));
   MUX4EHD U7144 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5686), 
	.D(\ram[239][12] ), 
	.C(\ram[237][12] ), 
	.B(\ram[238][12] ), 
	.A(\ram[236][12] ));
   MUX4EHD U7145 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5687), 
	.D(\ram[235][12] ), 
	.C(\ram[233][12] ), 
	.B(\ram[234][12] ), 
	.A(\ram[232][12] ));
   MUX4EHD U7146 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5688), 
	.D(\ram[231][12] ), 
	.C(\ram[229][12] ), 
	.B(\ram[230][12] ), 
	.A(\ram[228][12] ));
   MUX4EHD U7147 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5689), 
	.D(\ram[227][12] ), 
	.C(\ram[225][12] ), 
	.B(\ram[226][12] ), 
	.A(\ram[224][12] ));
   MUX4EHD U7148 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5690), 
	.D(n5686), 
	.C(n5688), 
	.B(n5687), 
	.A(n5689));
   MUX4EHD U7149 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5691), 
	.D(\ram[223][12] ), 
	.C(\ram[221][12] ), 
	.B(\ram[222][12] ), 
	.A(\ram[220][12] ));
   MUX4EHD U7150 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5692), 
	.D(\ram[219][12] ), 
	.C(\ram[217][12] ), 
	.B(\ram[218][12] ), 
	.A(\ram[216][12] ));
   MUX4EHD U7151 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5693), 
	.D(\ram[215][12] ), 
	.C(\ram[213][12] ), 
	.B(\ram[214][12] ), 
	.A(\ram[212][12] ));
   MUX4EHD U7152 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5694), 
	.D(\ram[211][12] ), 
	.C(\ram[209][12] ), 
	.B(\ram[210][12] ), 
	.A(\ram[208][12] ));
   MUX4EHD U7153 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5695), 
	.D(n5691), 
	.C(n5693), 
	.B(n5692), 
	.A(n5694));
   MUX4EHD U7154 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5696), 
	.D(\ram[207][12] ), 
	.C(\ram[205][12] ), 
	.B(\ram[206][12] ), 
	.A(\ram[204][12] ));
   MUX4EHD U7155 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5697), 
	.D(\ram[203][12] ), 
	.C(\ram[201][12] ), 
	.B(\ram[202][12] ), 
	.A(\ram[200][12] ));
   MUX4EHD U7156 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5698), 
	.D(\ram[199][12] ), 
	.C(\ram[197][12] ), 
	.B(\ram[198][12] ), 
	.A(\ram[196][12] ));
   MUX4EHD U7157 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5699), 
	.D(\ram[195][12] ), 
	.C(\ram[193][12] ), 
	.B(\ram[194][12] ), 
	.A(\ram[192][12] ));
   MUX4EHD U7158 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5700), 
	.D(n5696), 
	.C(n5698), 
	.B(n5697), 
	.A(n5699));
   MUX4EHD U7159 (.S1(n6038), 
	.S0(n7444), 
	.O(n5701), 
	.D(n5685), 
	.C(n5695), 
	.B(n5690), 
	.A(n5700));
   MUX4EHD U7160 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5702), 
	.D(\ram[191][12] ), 
	.C(\ram[189][12] ), 
	.B(\ram[190][12] ), 
	.A(\ram[188][12] ));
   MUX4EHD U7161 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5703), 
	.D(\ram[187][12] ), 
	.C(\ram[185][12] ), 
	.B(\ram[186][12] ), 
	.A(\ram[184][12] ));
   MUX4EHD U7162 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5704), 
	.D(\ram[183][12] ), 
	.C(\ram[181][12] ), 
	.B(\ram[182][12] ), 
	.A(\ram[180][12] ));
   MUX4EHD U7163 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5705), 
	.D(\ram[179][12] ), 
	.C(\ram[177][12] ), 
	.B(\ram[178][12] ), 
	.A(\ram[176][12] ));
   MUX4EHD U7164 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5706), 
	.D(n5702), 
	.C(n5704), 
	.B(n5703), 
	.A(n5705));
   MUX4EHD U7165 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5707), 
	.D(\ram[175][12] ), 
	.C(\ram[173][12] ), 
	.B(\ram[174][12] ), 
	.A(\ram[172][12] ));
   MUX4EHD U7166 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5708), 
	.D(\ram[171][12] ), 
	.C(\ram[169][12] ), 
	.B(\ram[170][12] ), 
	.A(\ram[168][12] ));
   MUX4EHD U7167 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5709), 
	.D(\ram[167][12] ), 
	.C(\ram[165][12] ), 
	.B(\ram[166][12] ), 
	.A(\ram[164][12] ));
   MUX4EHD U7168 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5710), 
	.D(\ram[163][12] ), 
	.C(\ram[161][12] ), 
	.B(\ram[162][12] ), 
	.A(\ram[160][12] ));
   MUX4EHD U7169 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5711), 
	.D(n5707), 
	.C(n5709), 
	.B(n5708), 
	.A(n5710));
   MUX4EHD U7170 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5712), 
	.D(\ram[159][12] ), 
	.C(\ram[157][12] ), 
	.B(\ram[158][12] ), 
	.A(\ram[156][12] ));
   MUX4EHD U7171 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5713), 
	.D(\ram[155][12] ), 
	.C(\ram[153][12] ), 
	.B(\ram[154][12] ), 
	.A(\ram[152][12] ));
   MUX4EHD U7172 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5714), 
	.D(\ram[151][12] ), 
	.C(\ram[149][12] ), 
	.B(\ram[150][12] ), 
	.A(\ram[148][12] ));
   MUX4EHD U7173 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5715), 
	.D(\ram[147][12] ), 
	.C(\ram[145][12] ), 
	.B(\ram[146][12] ), 
	.A(\ram[144][12] ));
   MUX4EHD U7174 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5716), 
	.D(n5712), 
	.C(n5714), 
	.B(n5713), 
	.A(n5715));
   MUX4EHD U7175 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5717), 
	.D(\ram[143][12] ), 
	.C(\ram[141][12] ), 
	.B(\ram[142][12] ), 
	.A(\ram[140][12] ));
   MUX4EHD U7176 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5718), 
	.D(\ram[139][12] ), 
	.C(\ram[137][12] ), 
	.B(\ram[138][12] ), 
	.A(\ram[136][12] ));
   MUX4EHD U7177 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5719), 
	.D(\ram[135][12] ), 
	.C(\ram[133][12] ), 
	.B(\ram[134][12] ), 
	.A(\ram[132][12] ));
   MUX4EHD U7178 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5720), 
	.D(\ram[131][12] ), 
	.C(\ram[129][12] ), 
	.B(\ram[130][12] ), 
	.A(\ram[128][12] ));
   MUX4EHD U7179 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5721), 
	.D(n5717), 
	.C(n5719), 
	.B(n5718), 
	.A(n5720));
   MUX4EHD U7180 (.S1(n6038), 
	.S0(n7444), 
	.O(n5722), 
	.D(n5706), 
	.C(n5716), 
	.B(n5711), 
	.A(n5721));
   MUX4EHD U7181 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5723), 
	.D(\ram[127][12] ), 
	.C(\ram[125][12] ), 
	.B(\ram[126][12] ), 
	.A(\ram[124][12] ));
   MUX4EHD U7182 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5724), 
	.D(\ram[123][12] ), 
	.C(\ram[121][12] ), 
	.B(\ram[122][12] ), 
	.A(\ram[120][12] ));
   MUX4EHD U7183 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5725), 
	.D(\ram[119][12] ), 
	.C(\ram[117][12] ), 
	.B(\ram[118][12] ), 
	.A(\ram[116][12] ));
   MUX4EHD U7184 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5726), 
	.D(\ram[115][12] ), 
	.C(\ram[113][12] ), 
	.B(\ram[114][12] ), 
	.A(\ram[112][12] ));
   MUX4EHD U7185 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5727), 
	.D(n5723), 
	.C(n5725), 
	.B(n5724), 
	.A(n5726));
   MUX4EHD U7186 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5728), 
	.D(\ram[111][12] ), 
	.C(\ram[109][12] ), 
	.B(\ram[110][12] ), 
	.A(\ram[108][12] ));
   MUX4EHD U7187 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5729), 
	.D(\ram[107][12] ), 
	.C(\ram[105][12] ), 
	.B(\ram[106][12] ), 
	.A(\ram[104][12] ));
   MUX4EHD U7188 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5730), 
	.D(\ram[103][12] ), 
	.C(\ram[101][12] ), 
	.B(\ram[102][12] ), 
	.A(\ram[100][12] ));
   MUX4EHD U7189 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5731), 
	.D(\ram[99][12] ), 
	.C(\ram[97][12] ), 
	.B(\ram[98][12] ), 
	.A(\ram[96][12] ));
   MUX4EHD U7190 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5732), 
	.D(n5728), 
	.C(n5730), 
	.B(n5729), 
	.A(n5731));
   MUX4EHD U7191 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5733), 
	.D(\ram[95][12] ), 
	.C(\ram[93][12] ), 
	.B(\ram[94][12] ), 
	.A(\ram[92][12] ));
   MUX4EHD U7192 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5734), 
	.D(\ram[91][12] ), 
	.C(\ram[89][12] ), 
	.B(\ram[90][12] ), 
	.A(\ram[88][12] ));
   MUX4EHD U7193 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5735), 
	.D(\ram[87][12] ), 
	.C(\ram[85][12] ), 
	.B(\ram[86][12] ), 
	.A(\ram[84][12] ));
   MUX4EHD U7194 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5736), 
	.D(\ram[83][12] ), 
	.C(\ram[81][12] ), 
	.B(\ram[82][12] ), 
	.A(\ram[80][12] ));
   MUX4EHD U7195 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5737), 
	.D(n5733), 
	.C(n5735), 
	.B(n5734), 
	.A(n5736));
   MUX4EHD U7196 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5738), 
	.D(\ram[79][12] ), 
	.C(\ram[77][12] ), 
	.B(\ram[78][12] ), 
	.A(\ram[76][12] ));
   MUX4EHD U7197 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5739), 
	.D(\ram[75][12] ), 
	.C(\ram[73][12] ), 
	.B(\ram[74][12] ), 
	.A(\ram[72][12] ));
   MUX4EHD U7198 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5740), 
	.D(\ram[71][12] ), 
	.C(\ram[69][12] ), 
	.B(\ram[70][12] ), 
	.A(\ram[68][12] ));
   MUX4EHD U7199 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5741), 
	.D(\ram[67][12] ), 
	.C(\ram[65][12] ), 
	.B(\ram[66][12] ), 
	.A(\ram[64][12] ));
   MUX4EHD U7200 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5742), 
	.D(n5738), 
	.C(n5740), 
	.B(n5739), 
	.A(n5741));
   MUX4EHD U7201 (.S1(n6038), 
	.S0(n7444), 
	.O(n5743), 
	.D(n5727), 
	.C(n5737), 
	.B(n5732), 
	.A(n5742));
   MUX4EHD U7202 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5744), 
	.D(\ram[63][12] ), 
	.C(\ram[61][12] ), 
	.B(\ram[62][12] ), 
	.A(\ram[60][12] ));
   MUX4EHD U7203 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5745), 
	.D(\ram[59][12] ), 
	.C(\ram[57][12] ), 
	.B(\ram[58][12] ), 
	.A(\ram[56][12] ));
   MUX4EHD U7204 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5746), 
	.D(\ram[55][12] ), 
	.C(\ram[53][12] ), 
	.B(\ram[54][12] ), 
	.A(\ram[52][12] ));
   MUX4EHD U7205 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5747), 
	.D(\ram[51][12] ), 
	.C(\ram[49][12] ), 
	.B(\ram[50][12] ), 
	.A(\ram[48][12] ));
   MUX4EHD U7206 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5748), 
	.D(n5744), 
	.C(n5746), 
	.B(n5745), 
	.A(n5747));
   MUX4EHD U7207 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5749), 
	.D(\ram[47][12] ), 
	.C(\ram[45][12] ), 
	.B(\ram[46][12] ), 
	.A(\ram[44][12] ));
   MUX4EHD U7208 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5750), 
	.D(\ram[43][12] ), 
	.C(\ram[41][12] ), 
	.B(\ram[42][12] ), 
	.A(\ram[40][12] ));
   MUX4EHD U7209 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5751), 
	.D(\ram[39][12] ), 
	.C(\ram[37][12] ), 
	.B(\ram[38][12] ), 
	.A(\ram[36][12] ));
   MUX4EHD U7210 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5752), 
	.D(\ram[35][12] ), 
	.C(\ram[33][12] ), 
	.B(\ram[34][12] ), 
	.A(\ram[32][12] ));
   MUX4EHD U7211 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5753), 
	.D(n5749), 
	.C(n5751), 
	.B(n5750), 
	.A(n5752));
   MUX4EHD U7212 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5754), 
	.D(\ram[31][12] ), 
	.C(\ram[29][12] ), 
	.B(\ram[30][12] ), 
	.A(\ram[28][12] ));
   MUX4EHD U7213 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5755), 
	.D(\ram[27][12] ), 
	.C(\ram[25][12] ), 
	.B(\ram[26][12] ), 
	.A(\ram[24][12] ));
   MUX4EHD U7214 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5756), 
	.D(\ram[23][12] ), 
	.C(\ram[21][12] ), 
	.B(\ram[22][12] ), 
	.A(\ram[20][12] ));
   MUX4EHD U7215 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5757), 
	.D(\ram[19][12] ), 
	.C(\ram[17][12] ), 
	.B(\ram[18][12] ), 
	.A(\ram[16][12] ));
   MUX4EHD U7216 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5758), 
	.D(n5754), 
	.C(n5756), 
	.B(n5755), 
	.A(n5757));
   MUX4EHD U7217 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5759), 
	.D(\ram[15][12] ), 
	.C(\ram[13][12] ), 
	.B(\ram[14][12] ), 
	.A(\ram[12][12] ));
   MUX4EHD U7218 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5760), 
	.D(\ram[11][12] ), 
	.C(\ram[9][12] ), 
	.B(\ram[10][12] ), 
	.A(\ram[8][12] ));
   MUX4EHD U7219 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5761), 
	.D(\ram[7][12] ), 
	.C(\ram[5][12] ), 
	.B(\ram[6][12] ), 
	.A(\ram[4][12] ));
   MUX4EHD U7220 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5762), 
	.D(\ram[3][12] ), 
	.C(\ram[1][12] ), 
	.B(\ram[2][12] ), 
	.A(\ram[0][12] ));
   MUX4EHD U7221 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5763), 
	.D(n5759), 
	.C(n5761), 
	.B(n5760), 
	.A(n5762));
   MUX4EHD U7222 (.S1(n6038), 
	.S0(n7444), 
	.O(n5764), 
	.D(n5748), 
	.C(n5758), 
	.B(n5753), 
	.A(n5763));
   MUX4EHD U7223 (.S1(n6469), 
	.S0(n6470), 
	.O(N4129), 
	.D(n5701), 
	.C(n5743), 
	.B(n5722), 
	.A(n5764));
   MUX4EHD U7224 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5765), 
	.D(\ram[255][13] ), 
	.C(\ram[253][13] ), 
	.B(\ram[254][13] ), 
	.A(\ram[252][13] ));
   MUX4EHD U7225 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5766), 
	.D(\ram[251][13] ), 
	.C(\ram[249][13] ), 
	.B(\ram[250][13] ), 
	.A(\ram[248][13] ));
   MUX4EHD U7226 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5767), 
	.D(\ram[247][13] ), 
	.C(\ram[245][13] ), 
	.B(\ram[246][13] ), 
	.A(\ram[244][13] ));
   MUX4EHD U7227 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5768), 
	.D(\ram[243][13] ), 
	.C(\ram[241][13] ), 
	.B(\ram[242][13] ), 
	.A(\ram[240][13] ));
   MUX4EHD U7228 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5769), 
	.D(n5765), 
	.C(n5767), 
	.B(n5766), 
	.A(n5768));
   MUX4EHD U7229 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5770), 
	.D(\ram[239][13] ), 
	.C(\ram[237][13] ), 
	.B(\ram[238][13] ), 
	.A(\ram[236][13] ));
   MUX4EHD U7230 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5771), 
	.D(\ram[235][13] ), 
	.C(\ram[233][13] ), 
	.B(\ram[234][13] ), 
	.A(\ram[232][13] ));
   MUX4EHD U7231 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5772), 
	.D(\ram[231][13] ), 
	.C(\ram[229][13] ), 
	.B(\ram[230][13] ), 
	.A(\ram[228][13] ));
   MUX4EHD U7232 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5773), 
	.D(\ram[227][13] ), 
	.C(\ram[225][13] ), 
	.B(\ram[226][13] ), 
	.A(\ram[224][13] ));
   MUX4EHD U7233 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5774), 
	.D(n5770), 
	.C(n5772), 
	.B(n5771), 
	.A(n5773));
   MUX4EHD U7234 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5775), 
	.D(\ram[223][13] ), 
	.C(\ram[221][13] ), 
	.B(\ram[222][13] ), 
	.A(\ram[220][13] ));
   MUX4EHD U7235 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5776), 
	.D(\ram[219][13] ), 
	.C(\ram[217][13] ), 
	.B(\ram[218][13] ), 
	.A(\ram[216][13] ));
   MUX4EHD U7236 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5777), 
	.D(\ram[215][13] ), 
	.C(\ram[213][13] ), 
	.B(\ram[214][13] ), 
	.A(\ram[212][13] ));
   MUX4EHD U7237 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5778), 
	.D(\ram[211][13] ), 
	.C(\ram[209][13] ), 
	.B(\ram[210][13] ), 
	.A(\ram[208][13] ));
   MUX4EHD U7238 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5779), 
	.D(n5775), 
	.C(n5777), 
	.B(n5776), 
	.A(n5778));
   MUX4EHD U7239 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5780), 
	.D(\ram[207][13] ), 
	.C(\ram[205][13] ), 
	.B(\ram[206][13] ), 
	.A(\ram[204][13] ));
   MUX4EHD U7240 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5781), 
	.D(\ram[203][13] ), 
	.C(\ram[201][13] ), 
	.B(\ram[202][13] ), 
	.A(\ram[200][13] ));
   MUX4EHD U7241 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5782), 
	.D(\ram[199][13] ), 
	.C(\ram[197][13] ), 
	.B(\ram[198][13] ), 
	.A(\ram[196][13] ));
   MUX4EHD U7242 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5783), 
	.D(\ram[195][13] ), 
	.C(\ram[193][13] ), 
	.B(\ram[194][13] ), 
	.A(\ram[192][13] ));
   MUX4EHD U7243 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5784), 
	.D(n5780), 
	.C(n5782), 
	.B(n5781), 
	.A(n5783));
   MUX4EHD U7244 (.S1(n6038), 
	.S0(n7444), 
	.O(n5785), 
	.D(n5769), 
	.C(n5779), 
	.B(n5774), 
	.A(n5784));
   MUX4EHD U7245 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5786), 
	.D(\ram[191][13] ), 
	.C(\ram[189][13] ), 
	.B(\ram[190][13] ), 
	.A(\ram[188][13] ));
   MUX4EHD U7246 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5787), 
	.D(\ram[187][13] ), 
	.C(\ram[185][13] ), 
	.B(\ram[186][13] ), 
	.A(\ram[184][13] ));
   MUX4EHD U7247 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5788), 
	.D(\ram[183][13] ), 
	.C(\ram[181][13] ), 
	.B(\ram[182][13] ), 
	.A(\ram[180][13] ));
   MUX4EHD U7248 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5789), 
	.D(\ram[179][13] ), 
	.C(\ram[177][13] ), 
	.B(\ram[178][13] ), 
	.A(\ram[176][13] ));
   MUX4EHD U7249 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5790), 
	.D(n5786), 
	.C(n5788), 
	.B(n5787), 
	.A(n5789));
   MUX4EHD U7250 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5791), 
	.D(\ram[175][13] ), 
	.C(\ram[173][13] ), 
	.B(\ram[174][13] ), 
	.A(\ram[172][13] ));
   MUX4EHD U7251 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5792), 
	.D(\ram[171][13] ), 
	.C(\ram[169][13] ), 
	.B(\ram[170][13] ), 
	.A(\ram[168][13] ));
   MUX4EHD U7252 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5793), 
	.D(\ram[167][13] ), 
	.C(\ram[165][13] ), 
	.B(\ram[166][13] ), 
	.A(\ram[164][13] ));
   MUX4EHD U7253 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5794), 
	.D(\ram[163][13] ), 
	.C(\ram[161][13] ), 
	.B(\ram[162][13] ), 
	.A(\ram[160][13] ));
   MUX4EHD U7254 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5795), 
	.D(n5791), 
	.C(n5793), 
	.B(n5792), 
	.A(n5794));
   MUX4EHD U7255 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5796), 
	.D(\ram[159][13] ), 
	.C(\ram[157][13] ), 
	.B(\ram[158][13] ), 
	.A(\ram[156][13] ));
   MUX4EHD U7256 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5797), 
	.D(\ram[155][13] ), 
	.C(\ram[153][13] ), 
	.B(\ram[154][13] ), 
	.A(\ram[152][13] ));
   MUX4EHD U7257 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5798), 
	.D(\ram[151][13] ), 
	.C(\ram[149][13] ), 
	.B(\ram[150][13] ), 
	.A(\ram[148][13] ));
   MUX4EHD U7258 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5799), 
	.D(\ram[147][13] ), 
	.C(\ram[145][13] ), 
	.B(\ram[146][13] ), 
	.A(\ram[144][13] ));
   MUX4EHD U7259 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5800), 
	.D(n5796), 
	.C(n5798), 
	.B(n5797), 
	.A(n5799));
   MUX4EHD U7260 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5801), 
	.D(\ram[143][13] ), 
	.C(\ram[141][13] ), 
	.B(\ram[142][13] ), 
	.A(\ram[140][13] ));
   MUX4EHD U7261 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5802), 
	.D(\ram[139][13] ), 
	.C(\ram[137][13] ), 
	.B(\ram[138][13] ), 
	.A(\ram[136][13] ));
   MUX4EHD U7262 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5803), 
	.D(\ram[135][13] ), 
	.C(\ram[133][13] ), 
	.B(\ram[134][13] ), 
	.A(\ram[132][13] ));
   MUX4EHD U7263 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5804), 
	.D(\ram[131][13] ), 
	.C(\ram[129][13] ), 
	.B(\ram[130][13] ), 
	.A(\ram[128][13] ));
   MUX4EHD U7264 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5805), 
	.D(n5801), 
	.C(n5803), 
	.B(n5802), 
	.A(n5804));
   MUX4EHD U7265 (.S1(n6038), 
	.S0(n7444), 
	.O(n5806), 
	.D(n5790), 
	.C(n5800), 
	.B(n5795), 
	.A(n5805));
   MUX4EHD U7266 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5807), 
	.D(\ram[127][13] ), 
	.C(\ram[125][13] ), 
	.B(\ram[126][13] ), 
	.A(\ram[124][13] ));
   MUX4EHD U7267 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5808), 
	.D(\ram[123][13] ), 
	.C(\ram[121][13] ), 
	.B(\ram[122][13] ), 
	.A(\ram[120][13] ));
   MUX4EHD U7268 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5809), 
	.D(\ram[119][13] ), 
	.C(\ram[117][13] ), 
	.B(\ram[118][13] ), 
	.A(\ram[116][13] ));
   MUX4EHD U7269 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5810), 
	.D(\ram[115][13] ), 
	.C(\ram[113][13] ), 
	.B(\ram[114][13] ), 
	.A(\ram[112][13] ));
   MUX4EHD U7270 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5811), 
	.D(n5807), 
	.C(n5809), 
	.B(n5808), 
	.A(n5810));
   MUX4EHD U7271 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5812), 
	.D(\ram[111][13] ), 
	.C(\ram[109][13] ), 
	.B(\ram[110][13] ), 
	.A(\ram[108][13] ));
   MUX4EHD U7272 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5813), 
	.D(\ram[107][13] ), 
	.C(\ram[105][13] ), 
	.B(\ram[106][13] ), 
	.A(\ram[104][13] ));
   MUX4EHD U7273 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5814), 
	.D(\ram[103][13] ), 
	.C(\ram[101][13] ), 
	.B(\ram[102][13] ), 
	.A(\ram[100][13] ));
   MUX4EHD U7274 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5815), 
	.D(\ram[99][13] ), 
	.C(\ram[97][13] ), 
	.B(\ram[98][13] ), 
	.A(\ram[96][13] ));
   MUX4EHD U7275 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5816), 
	.D(n5812), 
	.C(n5814), 
	.B(n5813), 
	.A(n5815));
   MUX4EHD U7276 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5817), 
	.D(\ram[95][13] ), 
	.C(\ram[93][13] ), 
	.B(\ram[94][13] ), 
	.A(\ram[92][13] ));
   MUX4EHD U7277 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5818), 
	.D(\ram[91][13] ), 
	.C(\ram[89][13] ), 
	.B(\ram[90][13] ), 
	.A(\ram[88][13] ));
   MUX4EHD U7278 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5819), 
	.D(\ram[87][13] ), 
	.C(\ram[85][13] ), 
	.B(\ram[86][13] ), 
	.A(\ram[84][13] ));
   MUX4EHD U7279 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5820), 
	.D(\ram[83][13] ), 
	.C(\ram[81][13] ), 
	.B(\ram[82][13] ), 
	.A(\ram[80][13] ));
   MUX4EHD U7280 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5821), 
	.D(n5817), 
	.C(n5819), 
	.B(n5818), 
	.A(n5820));
   MUX4EHD U7281 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5822), 
	.D(\ram[79][13] ), 
	.C(\ram[77][13] ), 
	.B(\ram[78][13] ), 
	.A(\ram[76][13] ));
   MUX4EHD U7282 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5823), 
	.D(\ram[75][13] ), 
	.C(\ram[73][13] ), 
	.B(\ram[74][13] ), 
	.A(\ram[72][13] ));
   MUX4EHD U7283 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5824), 
	.D(\ram[71][13] ), 
	.C(\ram[69][13] ), 
	.B(\ram[70][13] ), 
	.A(\ram[68][13] ));
   MUX4EHD U7284 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5825), 
	.D(\ram[67][13] ), 
	.C(\ram[65][13] ), 
	.B(\ram[66][13] ), 
	.A(\ram[64][13] ));
   MUX4EHD U7285 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5826), 
	.D(n5822), 
	.C(n5824), 
	.B(n5823), 
	.A(n5825));
   MUX4EHD U7286 (.S1(n6038), 
	.S0(n7444), 
	.O(n5827), 
	.D(n5811), 
	.C(n5821), 
	.B(n5816), 
	.A(n5826));
   MUX4EHD U7287 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5828), 
	.D(\ram[63][13] ), 
	.C(\ram[61][13] ), 
	.B(\ram[62][13] ), 
	.A(\ram[60][13] ));
   MUX4EHD U7288 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5829), 
	.D(\ram[59][13] ), 
	.C(\ram[57][13] ), 
	.B(\ram[58][13] ), 
	.A(\ram[56][13] ));
   MUX4EHD U7289 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5830), 
	.D(\ram[55][13] ), 
	.C(\ram[53][13] ), 
	.B(\ram[54][13] ), 
	.A(\ram[52][13] ));
   MUX4EHD U7290 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5831), 
	.D(\ram[51][13] ), 
	.C(\ram[49][13] ), 
	.B(\ram[50][13] ), 
	.A(\ram[48][13] ));
   MUX4EHD U7291 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5832), 
	.D(n5828), 
	.C(n5830), 
	.B(n5829), 
	.A(n5831));
   MUX4EHD U7292 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5833), 
	.D(\ram[47][13] ), 
	.C(\ram[45][13] ), 
	.B(\ram[46][13] ), 
	.A(\ram[44][13] ));
   MUX4EHD U7293 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5834), 
	.D(\ram[43][13] ), 
	.C(\ram[41][13] ), 
	.B(\ram[42][13] ), 
	.A(\ram[40][13] ));
   MUX4EHD U7294 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5835), 
	.D(\ram[39][13] ), 
	.C(\ram[37][13] ), 
	.B(\ram[38][13] ), 
	.A(\ram[36][13] ));
   MUX4EHD U7295 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5836), 
	.D(\ram[35][13] ), 
	.C(\ram[33][13] ), 
	.B(\ram[34][13] ), 
	.A(\ram[32][13] ));
   MUX4EHD U7296 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5837), 
	.D(n5833), 
	.C(n5835), 
	.B(n5834), 
	.A(n5836));
   MUX4EHD U7297 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5838), 
	.D(\ram[31][13] ), 
	.C(\ram[29][13] ), 
	.B(\ram[30][13] ), 
	.A(\ram[28][13] ));
   MUX4EHD U7298 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5839), 
	.D(\ram[27][13] ), 
	.C(\ram[25][13] ), 
	.B(\ram[26][13] ), 
	.A(\ram[24][13] ));
   MUX4EHD U7299 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5840), 
	.D(\ram[23][13] ), 
	.C(\ram[21][13] ), 
	.B(\ram[22][13] ), 
	.A(\ram[20][13] ));
   MUX4EHD U7300 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5841), 
	.D(\ram[19][13] ), 
	.C(\ram[17][13] ), 
	.B(\ram[18][13] ), 
	.A(\ram[16][13] ));
   MUX4EHD U7301 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5842), 
	.D(n5838), 
	.C(n5840), 
	.B(n5839), 
	.A(n5841));
   MUX4EHD U7302 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5843), 
	.D(\ram[15][13] ), 
	.C(\ram[13][13] ), 
	.B(\ram[14][13] ), 
	.A(\ram[12][13] ));
   MUX4EHD U7303 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5844), 
	.D(\ram[11][13] ), 
	.C(\ram[9][13] ), 
	.B(\ram[10][13] ), 
	.A(\ram[8][13] ));
   MUX4EHD U7304 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5845), 
	.D(\ram[7][13] ), 
	.C(\ram[5][13] ), 
	.B(\ram[6][13] ), 
	.A(\ram[4][13] ));
   MUX4EHD U7305 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5846), 
	.D(\ram[3][13] ), 
	.C(\ram[1][13] ), 
	.B(\ram[2][13] ), 
	.A(\ram[0][13] ));
   MUX4EHD U7306 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5847), 
	.D(n5843), 
	.C(n5845), 
	.B(n5844), 
	.A(n5846));
   MUX4EHD U7307 (.S1(n6038), 
	.S0(n7444), 
	.O(n5848), 
	.D(n5832), 
	.C(n5842), 
	.B(n5837), 
	.A(n5847));
   MUX4EHD U7308 (.S1(n6469), 
	.S0(n6470), 
	.O(N4128), 
	.D(n5785), 
	.C(n5827), 
	.B(n5806), 
	.A(n5848));
   MUX4EHD U7309 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5849), 
	.D(\ram[255][14] ), 
	.C(\ram[253][14] ), 
	.B(\ram[254][14] ), 
	.A(\ram[252][14] ));
   MUX4EHD U7310 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5850), 
	.D(\ram[251][14] ), 
	.C(\ram[249][14] ), 
	.B(\ram[250][14] ), 
	.A(\ram[248][14] ));
   MUX4EHD U7311 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5851), 
	.D(\ram[247][14] ), 
	.C(\ram[245][14] ), 
	.B(\ram[246][14] ), 
	.A(\ram[244][14] ));
   MUX4EHD U7312 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5852), 
	.D(\ram[243][14] ), 
	.C(\ram[241][14] ), 
	.B(\ram[242][14] ), 
	.A(\ram[240][14] ));
   MUX4EHD U7313 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5853), 
	.D(n5849), 
	.C(n5851), 
	.B(n5850), 
	.A(n5852));
   MUX4EHD U7314 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5854), 
	.D(\ram[239][14] ), 
	.C(\ram[237][14] ), 
	.B(\ram[238][14] ), 
	.A(\ram[236][14] ));
   MUX4EHD U7315 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5855), 
	.D(\ram[235][14] ), 
	.C(\ram[233][14] ), 
	.B(\ram[234][14] ), 
	.A(\ram[232][14] ));
   MUX4EHD U7316 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5856), 
	.D(\ram[231][14] ), 
	.C(\ram[229][14] ), 
	.B(\ram[230][14] ), 
	.A(\ram[228][14] ));
   MUX4EHD U7317 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5857), 
	.D(\ram[227][14] ), 
	.C(\ram[225][14] ), 
	.B(\ram[226][14] ), 
	.A(\ram[224][14] ));
   MUX4EHD U7318 (.S1(n6136), 
	.S0(n7442), 
	.O(n5858), 
	.D(n5854), 
	.C(n5856), 
	.B(n5855), 
	.A(n5857));
   MUX4EHD U7319 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5859), 
	.D(\ram[223][14] ), 
	.C(\ram[221][14] ), 
	.B(\ram[222][14] ), 
	.A(\ram[220][14] ));
   MUX4EHD U7320 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5860), 
	.D(\ram[219][14] ), 
	.C(\ram[217][14] ), 
	.B(\ram[218][14] ), 
	.A(\ram[216][14] ));
   MUX4EHD U7321 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5861), 
	.D(\ram[215][14] ), 
	.C(\ram[213][14] ), 
	.B(\ram[214][14] ), 
	.A(\ram[212][14] ));
   MUX4EHD U7322 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5862), 
	.D(\ram[211][14] ), 
	.C(\ram[209][14] ), 
	.B(\ram[210][14] ), 
	.A(\ram[208][14] ));
   MUX4EHD U7323 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5863), 
	.D(n5859), 
	.C(n5861), 
	.B(n5860), 
	.A(n5862));
   MUX4EHD U7324 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5864), 
	.D(\ram[207][14] ), 
	.C(\ram[205][14] ), 
	.B(\ram[206][14] ), 
	.A(\ram[204][14] ));
   MUX4EHD U7325 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5865), 
	.D(\ram[203][14] ), 
	.C(\ram[201][14] ), 
	.B(\ram[202][14] ), 
	.A(\ram[200][14] ));
   MUX4EHD U7326 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5866), 
	.D(\ram[199][14] ), 
	.C(\ram[197][14] ), 
	.B(\ram[198][14] ), 
	.A(\ram[196][14] ));
   MUX4EHD U7327 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5867), 
	.D(\ram[195][14] ), 
	.C(\ram[193][14] ), 
	.B(\ram[194][14] ), 
	.A(\ram[192][14] ));
   MUX4EHD U7328 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5868), 
	.D(n5864), 
	.C(n5866), 
	.B(n5865), 
	.A(n5867));
   MUX4EHD U7329 (.S1(n6038), 
	.S0(n7444), 
	.O(n5869), 
	.D(n5853), 
	.C(n5863), 
	.B(n5858), 
	.A(n5868));
   MUX4EHD U7330 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5870), 
	.D(\ram[191][14] ), 
	.C(\ram[189][14] ), 
	.B(\ram[190][14] ), 
	.A(\ram[188][14] ));
   MUX4EHD U7331 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5871), 
	.D(\ram[187][14] ), 
	.C(\ram[185][14] ), 
	.B(\ram[186][14] ), 
	.A(\ram[184][14] ));
   MUX4EHD U7332 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5872), 
	.D(\ram[183][14] ), 
	.C(\ram[181][14] ), 
	.B(\ram[182][14] ), 
	.A(\ram[180][14] ));
   MUX4EHD U7333 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5873), 
	.D(\ram[179][14] ), 
	.C(\ram[177][14] ), 
	.B(\ram[178][14] ), 
	.A(\ram[176][14] ));
   MUX4EHD U7334 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5874), 
	.D(n5870), 
	.C(n5872), 
	.B(n5871), 
	.A(n5873));
   MUX4EHD U7335 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5875), 
	.D(\ram[175][14] ), 
	.C(\ram[173][14] ), 
	.B(\ram[174][14] ), 
	.A(\ram[172][14] ));
   MUX4EHD U7336 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5876), 
	.D(\ram[171][14] ), 
	.C(\ram[169][14] ), 
	.B(\ram[170][14] ), 
	.A(\ram[168][14] ));
   MUX4EHD U7337 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5877), 
	.D(\ram[167][14] ), 
	.C(\ram[165][14] ), 
	.B(\ram[166][14] ), 
	.A(\ram[164][14] ));
   MUX4EHD U7338 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5878), 
	.D(\ram[163][14] ), 
	.C(\ram[161][14] ), 
	.B(\ram[162][14] ), 
	.A(\ram[160][14] ));
   MUX4EHD U7339 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5879), 
	.D(n5875), 
	.C(n5877), 
	.B(n5876), 
	.A(n5878));
   MUX4EHD U7340 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5880), 
	.D(\ram[159][14] ), 
	.C(\ram[157][14] ), 
	.B(\ram[158][14] ), 
	.A(\ram[156][14] ));
   MUX4EHD U7341 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5881), 
	.D(\ram[155][14] ), 
	.C(\ram[153][14] ), 
	.B(\ram[154][14] ), 
	.A(\ram[152][14] ));
   MUX4EHD U7342 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5882), 
	.D(\ram[151][14] ), 
	.C(\ram[149][14] ), 
	.B(\ram[150][14] ), 
	.A(\ram[148][14] ));
   MUX4EHD U7343 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5883), 
	.D(\ram[147][14] ), 
	.C(\ram[145][14] ), 
	.B(\ram[146][14] ), 
	.A(\ram[144][14] ));
   MUX4EHD U7344 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5884), 
	.D(n5880), 
	.C(n5882), 
	.B(n5881), 
	.A(n5883));
   MUX4EHD U7345 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5885), 
	.D(\ram[143][14] ), 
	.C(\ram[141][14] ), 
	.B(\ram[142][14] ), 
	.A(\ram[140][14] ));
   MUX4EHD U7346 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5886), 
	.D(\ram[139][14] ), 
	.C(\ram[137][14] ), 
	.B(\ram[138][14] ), 
	.A(\ram[136][14] ));
   MUX4EHD U7347 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5887), 
	.D(\ram[135][14] ), 
	.C(\ram[133][14] ), 
	.B(\ram[134][14] ), 
	.A(\ram[132][14] ));
   MUX4EHD U7348 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5888), 
	.D(\ram[131][14] ), 
	.C(\ram[129][14] ), 
	.B(\ram[130][14] ), 
	.A(\ram[128][14] ));
   MUX4EHD U7349 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5889), 
	.D(n5885), 
	.C(n5887), 
	.B(n5886), 
	.A(n5888));
   MUX4EHD U7350 (.S1(n6038), 
	.S0(n7444), 
	.O(n5890), 
	.D(n5874), 
	.C(n5884), 
	.B(n5879), 
	.A(n5889));
   MUX4EHD U7351 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5891), 
	.D(\ram[127][14] ), 
	.C(\ram[125][14] ), 
	.B(\ram[126][14] ), 
	.A(\ram[124][14] ));
   MUX4EHD U7352 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5892), 
	.D(\ram[123][14] ), 
	.C(\ram[121][14] ), 
	.B(\ram[122][14] ), 
	.A(\ram[120][14] ));
   MUX4EHD U7353 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5893), 
	.D(\ram[119][14] ), 
	.C(\ram[117][14] ), 
	.B(\ram[118][14] ), 
	.A(\ram[116][14] ));
   MUX4EHD U7354 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5894), 
	.D(\ram[115][14] ), 
	.C(\ram[113][14] ), 
	.B(\ram[114][14] ), 
	.A(\ram[112][14] ));
   MUX4EHD U7355 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5895), 
	.D(n5891), 
	.C(n5893), 
	.B(n5892), 
	.A(n5894));
   MUX4EHD U7356 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5896), 
	.D(\ram[111][14] ), 
	.C(\ram[109][14] ), 
	.B(\ram[110][14] ), 
	.A(\ram[108][14] ));
   MUX4EHD U7357 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5897), 
	.D(\ram[107][14] ), 
	.C(\ram[105][14] ), 
	.B(\ram[106][14] ), 
	.A(\ram[104][14] ));
   MUX4EHD U7358 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5898), 
	.D(\ram[103][14] ), 
	.C(\ram[101][14] ), 
	.B(\ram[102][14] ), 
	.A(\ram[100][14] ));
   MUX4EHD U7359 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5899), 
	.D(\ram[99][14] ), 
	.C(\ram[97][14] ), 
	.B(\ram[98][14] ), 
	.A(\ram[96][14] ));
   MUX4EHD U7360 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5900), 
	.D(n5896), 
	.C(n5898), 
	.B(n5897), 
	.A(n5899));
   MUX4EHD U7361 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5901), 
	.D(\ram[95][14] ), 
	.C(\ram[93][14] ), 
	.B(\ram[94][14] ), 
	.A(\ram[92][14] ));
   MUX4EHD U7362 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5902), 
	.D(\ram[91][14] ), 
	.C(\ram[89][14] ), 
	.B(\ram[90][14] ), 
	.A(\ram[88][14] ));
   MUX4EHD U7363 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5903), 
	.D(\ram[87][14] ), 
	.C(\ram[85][14] ), 
	.B(\ram[86][14] ), 
	.A(\ram[84][14] ));
   MUX4EHD U7364 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5904), 
	.D(\ram[83][14] ), 
	.C(\ram[81][14] ), 
	.B(\ram[82][14] ), 
	.A(\ram[80][14] ));
   MUX4EHD U7365 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5905), 
	.D(n5901), 
	.C(n5903), 
	.B(n5902), 
	.A(n5904));
   MUX4EHD U7366 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5906), 
	.D(\ram[79][14] ), 
	.C(\ram[77][14] ), 
	.B(\ram[78][14] ), 
	.A(\ram[76][14] ));
   MUX4EHD U7367 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5907), 
	.D(\ram[75][14] ), 
	.C(\ram[73][14] ), 
	.B(\ram[74][14] ), 
	.A(\ram[72][14] ));
   MUX4EHD U7368 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5908), 
	.D(\ram[71][14] ), 
	.C(\ram[69][14] ), 
	.B(\ram[70][14] ), 
	.A(\ram[68][14] ));
   MUX4EHD U7369 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5909), 
	.D(\ram[67][14] ), 
	.C(\ram[65][14] ), 
	.B(\ram[66][14] ), 
	.A(\ram[64][14] ));
   MUX4EHD U7370 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5910), 
	.D(n5906), 
	.C(n5908), 
	.B(n5907), 
	.A(n5909));
   MUX4EHD U7371 (.S1(n6038), 
	.S0(n7444), 
	.O(n5911), 
	.D(n5895), 
	.C(n5905), 
	.B(n5900), 
	.A(n5910));
   MUX4EHD U7372 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5912), 
	.D(\ram[63][14] ), 
	.C(\ram[61][14] ), 
	.B(\ram[62][14] ), 
	.A(\ram[60][14] ));
   MUX4EHD U7373 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5913), 
	.D(\ram[59][14] ), 
	.C(\ram[57][14] ), 
	.B(\ram[58][14] ), 
	.A(\ram[56][14] ));
   MUX4EHD U7374 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5914), 
	.D(\ram[55][14] ), 
	.C(\ram[53][14] ), 
	.B(\ram[54][14] ), 
	.A(\ram[52][14] ));
   MUX4EHD U7375 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5915), 
	.D(\ram[51][14] ), 
	.C(\ram[49][14] ), 
	.B(\ram[50][14] ), 
	.A(\ram[48][14] ));
   MUX4EHD U7376 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5916), 
	.D(n5912), 
	.C(n5914), 
	.B(n5913), 
	.A(n5915));
   MUX4EHD U7377 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5917), 
	.D(\ram[47][14] ), 
	.C(\ram[45][14] ), 
	.B(\ram[46][14] ), 
	.A(\ram[44][14] ));
   MUX4EHD U7378 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5918), 
	.D(\ram[43][14] ), 
	.C(\ram[41][14] ), 
	.B(\ram[42][14] ), 
	.A(\ram[40][14] ));
   MUX4EHD U7379 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5919), 
	.D(\ram[39][14] ), 
	.C(\ram[37][14] ), 
	.B(\ram[38][14] ), 
	.A(\ram[36][14] ));
   MUX4EHD U7380 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5920), 
	.D(\ram[35][14] ), 
	.C(\ram[33][14] ), 
	.B(\ram[34][14] ), 
	.A(\ram[32][14] ));
   MUX4EHD U7381 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5921), 
	.D(n5917), 
	.C(n5919), 
	.B(n5918), 
	.A(n5920));
   MUX4EHD U7382 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5922), 
	.D(\ram[31][14] ), 
	.C(\ram[29][14] ), 
	.B(\ram[30][14] ), 
	.A(\ram[28][14] ));
   MUX4EHD U7383 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5923), 
	.D(\ram[27][14] ), 
	.C(\ram[25][14] ), 
	.B(\ram[26][14] ), 
	.A(\ram[24][14] ));
   MUX4EHD U7384 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5924), 
	.D(\ram[23][14] ), 
	.C(\ram[21][14] ), 
	.B(\ram[22][14] ), 
	.A(\ram[20][14] ));
   MUX4EHD U7385 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5925), 
	.D(\ram[19][14] ), 
	.C(\ram[17][14] ), 
	.B(\ram[18][14] ), 
	.A(\ram[16][14] ));
   MUX4EHD U7386 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5926), 
	.D(n5922), 
	.C(n5924), 
	.B(n5923), 
	.A(n5925));
   MUX4EHD U7387 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5927), 
	.D(\ram[15][14] ), 
	.C(\ram[13][14] ), 
	.B(\ram[14][14] ), 
	.A(\ram[12][14] ));
   MUX4EHD U7388 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5928), 
	.D(\ram[11][14] ), 
	.C(\ram[9][14] ), 
	.B(\ram[10][14] ), 
	.A(\ram[8][14] ));
   MUX4EHD U7389 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5929), 
	.D(\ram[7][14] ), 
	.C(\ram[5][14] ), 
	.B(\ram[6][14] ), 
	.A(\ram[4][14] ));
   MUX4EHD U7390 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n5930), 
	.D(\ram[3][14] ), 
	.C(\ram[1][14] ), 
	.B(\ram[2][14] ), 
	.A(\ram[0][14] ));
   MUX4EHD U7391 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5931), 
	.D(n5927), 
	.C(n5929), 
	.B(n5928), 
	.A(n5930));
   MUX4EHD U7392 (.S1(n6038), 
	.S0(n7444), 
	.O(n5932), 
	.D(n5916), 
	.C(n5926), 
	.B(n5921), 
	.A(n5931));
   MUX4EHD U7393 (.S1(n6469), 
	.S0(n6470), 
	.O(N4127), 
	.D(n5869), 
	.C(n5911), 
	.B(n5890), 
	.A(n5932));
   MUX4EHD U7394 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5933), 
	.D(\ram[255][15] ), 
	.C(\ram[253][15] ), 
	.B(\ram[254][15] ), 
	.A(\ram[252][15] ));
   MUX4EHD U7395 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5934), 
	.D(\ram[251][15] ), 
	.C(\ram[249][15] ), 
	.B(\ram[250][15] ), 
	.A(\ram[248][15] ));
   MUX4EHD U7396 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5935), 
	.D(\ram[247][15] ), 
	.C(\ram[245][15] ), 
	.B(\ram[246][15] ), 
	.A(\ram[244][15] ));
   MUX4EHD U7397 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5936), 
	.D(\ram[243][15] ), 
	.C(\ram[241][15] ), 
	.B(\ram[242][15] ), 
	.A(\ram[240][15] ));
   MUX4EHD U7398 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5937), 
	.D(n5933), 
	.C(n5935), 
	.B(n5934), 
	.A(n5936));
   MUX4EHD U7399 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5938), 
	.D(\ram[239][15] ), 
	.C(\ram[237][15] ), 
	.B(\ram[238][15] ), 
	.A(\ram[236][15] ));
   MUX4EHD U7400 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5939), 
	.D(\ram[235][15] ), 
	.C(\ram[233][15] ), 
	.B(\ram[234][15] ), 
	.A(\ram[232][15] ));
   MUX4EHD U7401 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5940), 
	.D(\ram[231][15] ), 
	.C(\ram[229][15] ), 
	.B(\ram[230][15] ), 
	.A(\ram[228][15] ));
   MUX4EHD U7402 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5941), 
	.D(\ram[227][15] ), 
	.C(\ram[225][15] ), 
	.B(\ram[226][15] ), 
	.A(\ram[224][15] ));
   MUX4EHD U7403 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5942), 
	.D(n5938), 
	.C(n5940), 
	.B(n5939), 
	.A(n5941));
   MUX4EHD U7404 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5943), 
	.D(\ram[223][15] ), 
	.C(\ram[221][15] ), 
	.B(\ram[222][15] ), 
	.A(\ram[220][15] ));
   MUX4EHD U7405 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5944), 
	.D(\ram[219][15] ), 
	.C(\ram[217][15] ), 
	.B(\ram[218][15] ), 
	.A(\ram[216][15] ));
   MUX4EHD U7406 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5945), 
	.D(\ram[215][15] ), 
	.C(\ram[213][15] ), 
	.B(\ram[214][15] ), 
	.A(\ram[212][15] ));
   MUX4EHD U7407 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5946), 
	.D(\ram[211][15] ), 
	.C(\ram[209][15] ), 
	.B(\ram[210][15] ), 
	.A(\ram[208][15] ));
   MUX4EHD U7408 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5947), 
	.D(n5943), 
	.C(n5945), 
	.B(n5944), 
	.A(n5946));
   MUX4EHD U7409 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5948), 
	.D(\ram[207][15] ), 
	.C(\ram[205][15] ), 
	.B(\ram[206][15] ), 
	.A(\ram[204][15] ));
   MUX4EHD U7410 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5949), 
	.D(\ram[203][15] ), 
	.C(\ram[201][15] ), 
	.B(\ram[202][15] ), 
	.A(\ram[200][15] ));
   MUX4EHD U7411 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5950), 
	.D(\ram[199][15] ), 
	.C(\ram[197][15] ), 
	.B(\ram[198][15] ), 
	.A(\ram[196][15] ));
   MUX4EHD U7412 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5951), 
	.D(\ram[195][15] ), 
	.C(\ram[193][15] ), 
	.B(\ram[194][15] ), 
	.A(\ram[192][15] ));
   MUX4EHD U7413 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5952), 
	.D(n5948), 
	.C(n5950), 
	.B(n5949), 
	.A(n5951));
   MUX4EHD U7414 (.S1(n6038), 
	.S0(n7444), 
	.O(n5953), 
	.D(n5937), 
	.C(n5947), 
	.B(n5942), 
	.A(n5952));
   MUX4EHD U7415 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5954), 
	.D(\ram[191][15] ), 
	.C(\ram[189][15] ), 
	.B(\ram[190][15] ), 
	.A(\ram[188][15] ));
   MUX4EHD U7416 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5955), 
	.D(\ram[187][15] ), 
	.C(\ram[185][15] ), 
	.B(\ram[186][15] ), 
	.A(\ram[184][15] ));
   MUX4EHD U7417 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5956), 
	.D(\ram[183][15] ), 
	.C(\ram[181][15] ), 
	.B(\ram[182][15] ), 
	.A(\ram[180][15] ));
   MUX4EHD U7418 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5957), 
	.D(\ram[179][15] ), 
	.C(\ram[177][15] ), 
	.B(\ram[178][15] ), 
	.A(\ram[176][15] ));
   MUX4EHD U7419 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5958), 
	.D(n5954), 
	.C(n5956), 
	.B(n5955), 
	.A(n5957));
   MUX4EHD U7420 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5959), 
	.D(\ram[175][15] ), 
	.C(\ram[173][15] ), 
	.B(\ram[174][15] ), 
	.A(\ram[172][15] ));
   MUX4EHD U7421 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5960), 
	.D(\ram[171][15] ), 
	.C(\ram[169][15] ), 
	.B(\ram[170][15] ), 
	.A(\ram[168][15] ));
   MUX4EHD U7422 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5961), 
	.D(\ram[167][15] ), 
	.C(\ram[165][15] ), 
	.B(\ram[166][15] ), 
	.A(\ram[164][15] ));
   MUX4EHD U7423 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5962), 
	.D(\ram[163][15] ), 
	.C(\ram[161][15] ), 
	.B(\ram[162][15] ), 
	.A(\ram[160][15] ));
   MUX4EHD U7424 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5963), 
	.D(n5959), 
	.C(n5961), 
	.B(n5960), 
	.A(n5962));
   MUX4EHD U7425 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5964), 
	.D(\ram[159][15] ), 
	.C(\ram[157][15] ), 
	.B(\ram[158][15] ), 
	.A(\ram[156][15] ));
   MUX4EHD U7426 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5965), 
	.D(\ram[155][15] ), 
	.C(\ram[153][15] ), 
	.B(\ram[154][15] ), 
	.A(\ram[152][15] ));
   MUX4EHD U7427 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5966), 
	.D(\ram[151][15] ), 
	.C(\ram[149][15] ), 
	.B(\ram[150][15] ), 
	.A(\ram[148][15] ));
   MUX4EHD U7428 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5967), 
	.D(\ram[147][15] ), 
	.C(\ram[145][15] ), 
	.B(\ram[146][15] ), 
	.A(\ram[144][15] ));
   MUX4EHD U7429 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5968), 
	.D(n5964), 
	.C(n5966), 
	.B(n5965), 
	.A(n5967));
   MUX4EHD U7430 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5969), 
	.D(\ram[143][15] ), 
	.C(\ram[141][15] ), 
	.B(\ram[142][15] ), 
	.A(\ram[140][15] ));
   MUX4EHD U7431 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5970), 
	.D(\ram[139][15] ), 
	.C(\ram[137][15] ), 
	.B(\ram[138][15] ), 
	.A(\ram[136][15] ));
   MUX4EHD U7432 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5971), 
	.D(\ram[135][15] ), 
	.C(\ram[133][15] ), 
	.B(\ram[134][15] ), 
	.A(\ram[132][15] ));
   MUX4EHD U7433 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5972), 
	.D(\ram[131][15] ), 
	.C(\ram[129][15] ), 
	.B(\ram[130][15] ), 
	.A(\ram[128][15] ));
   MUX4EHD U7434 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5973), 
	.D(n5969), 
	.C(n5971), 
	.B(n5970), 
	.A(n5972));
   MUX4EHD U7435 (.S1(n6038), 
	.S0(n7444), 
	.O(n5974), 
	.D(n5958), 
	.C(n5968), 
	.B(n5963), 
	.A(n5973));
   MUX4EHD U7436 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5975), 
	.D(\ram[127][15] ), 
	.C(\ram[125][15] ), 
	.B(\ram[126][15] ), 
	.A(\ram[124][15] ));
   MUX4EHD U7437 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5976), 
	.D(\ram[123][15] ), 
	.C(\ram[121][15] ), 
	.B(\ram[122][15] ), 
	.A(\ram[120][15] ));
   MUX4EHD U7438 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5977), 
	.D(\ram[119][15] ), 
	.C(\ram[117][15] ), 
	.B(\ram[118][15] ), 
	.A(\ram[116][15] ));
   MUX4EHD U7439 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5978), 
	.D(\ram[115][15] ), 
	.C(\ram[113][15] ), 
	.B(\ram[114][15] ), 
	.A(\ram[112][15] ));
   MUX4EHD U7440 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5979), 
	.D(n5975), 
	.C(n5977), 
	.B(n5976), 
	.A(n5978));
   MUX4EHD U7441 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5980), 
	.D(\ram[111][15] ), 
	.C(\ram[109][15] ), 
	.B(\ram[110][15] ), 
	.A(\ram[108][15] ));
   MUX4EHD U7442 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5981), 
	.D(\ram[107][15] ), 
	.C(\ram[105][15] ), 
	.B(\ram[106][15] ), 
	.A(\ram[104][15] ));
   MUX4EHD U7443 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5982), 
	.D(\ram[103][15] ), 
	.C(\ram[101][15] ), 
	.B(\ram[102][15] ), 
	.A(\ram[100][15] ));
   MUX4EHD U7444 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5983), 
	.D(\ram[99][15] ), 
	.C(\ram[97][15] ), 
	.B(\ram[98][15] ), 
	.A(\ram[96][15] ));
   MUX4EHD U7445 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5984), 
	.D(n5980), 
	.C(n5982), 
	.B(n5981), 
	.A(n5983));
   MUX4EHD U7446 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5985), 
	.D(\ram[95][15] ), 
	.C(\ram[93][15] ), 
	.B(\ram[94][15] ), 
	.A(\ram[92][15] ));
   MUX4EHD U7447 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5986), 
	.D(\ram[91][15] ), 
	.C(\ram[89][15] ), 
	.B(\ram[90][15] ), 
	.A(\ram[88][15] ));
   MUX4EHD U7448 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5987), 
	.D(\ram[87][15] ), 
	.C(\ram[85][15] ), 
	.B(\ram[86][15] ), 
	.A(\ram[84][15] ));
   MUX4EHD U7449 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5988), 
	.D(\ram[83][15] ), 
	.C(\ram[81][15] ), 
	.B(\ram[82][15] ), 
	.A(\ram[80][15] ));
   MUX4EHD U7450 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5989), 
	.D(n5985), 
	.C(n5987), 
	.B(n5986), 
	.A(n5988));
   MUX4EHD U7451 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5990), 
	.D(\ram[79][15] ), 
	.C(\ram[77][15] ), 
	.B(\ram[78][15] ), 
	.A(\ram[76][15] ));
   MUX4EHD U7452 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5991), 
	.D(\ram[75][15] ), 
	.C(\ram[73][15] ), 
	.B(\ram[74][15] ), 
	.A(\ram[72][15] ));
   MUX4EHD U7453 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5992), 
	.D(\ram[71][15] ), 
	.C(\ram[69][15] ), 
	.B(\ram[70][15] ), 
	.A(\ram[68][15] ));
   MUX4EHD U7454 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5993), 
	.D(\ram[67][15] ), 
	.C(\ram[65][15] ), 
	.B(\ram[66][15] ), 
	.A(\ram[64][15] ));
   MUX4EHD U7455 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5994), 
	.D(n5990), 
	.C(n5992), 
	.B(n5991), 
	.A(n5993));
   MUX4EHD U7456 (.S1(n6038), 
	.S0(n7444), 
	.O(n5995), 
	.D(n5979), 
	.C(n5989), 
	.B(n5984), 
	.A(n5994));
   MUX4EHD U7457 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5996), 
	.D(\ram[63][15] ), 
	.C(\ram[61][15] ), 
	.B(\ram[62][15] ), 
	.A(\ram[60][15] ));
   MUX4EHD U7458 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5997), 
	.D(\ram[59][15] ), 
	.C(\ram[57][15] ), 
	.B(\ram[58][15] ), 
	.A(\ram[56][15] ));
   MUX4EHD U7459 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5998), 
	.D(\ram[55][15] ), 
	.C(\ram[53][15] ), 
	.B(\ram[54][15] ), 
	.A(\ram[52][15] ));
   MUX4EHD U7460 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5999), 
	.D(\ram[51][15] ), 
	.C(\ram[49][15] ), 
	.B(\ram[50][15] ), 
	.A(\ram[48][15] ));
   MUX4EHD U7461 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n6000), 
	.D(n5996), 
	.C(n5998), 
	.B(n5997), 
	.A(n5999));
   MUX4EHD U7462 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6001), 
	.D(\ram[47][15] ), 
	.C(\ram[45][15] ), 
	.B(\ram[46][15] ), 
	.A(\ram[44][15] ));
   MUX4EHD U7463 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6002), 
	.D(\ram[43][15] ), 
	.C(\ram[41][15] ), 
	.B(\ram[42][15] ), 
	.A(\ram[40][15] ));
   MUX4EHD U7464 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6003), 
	.D(\ram[39][15] ), 
	.C(\ram[37][15] ), 
	.B(\ram[38][15] ), 
	.A(\ram[36][15] ));
   MUX4EHD U7465 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6004), 
	.D(\ram[35][15] ), 
	.C(\ram[33][15] ), 
	.B(\ram[34][15] ), 
	.A(\ram[32][15] ));
   MUX4EHD U7466 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n6005), 
	.D(n6001), 
	.C(n6003), 
	.B(n6002), 
	.A(n6004));
   MUX4EHD U7467 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n6006), 
	.D(\ram[31][15] ), 
	.C(\ram[29][15] ), 
	.B(\ram[30][15] ), 
	.A(\ram[28][15] ));
   MUX4EHD U7468 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n6007), 
	.D(\ram[27][15] ), 
	.C(\ram[25][15] ), 
	.B(\ram[26][15] ), 
	.A(\ram[24][15] ));
   MUX4EHD U7469 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n6008), 
	.D(\ram[23][15] ), 
	.C(\ram[21][15] ), 
	.B(\ram[22][15] ), 
	.A(\ram[20][15] ));
   MUX4EHD U7470 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n6009), 
	.D(\ram[19][15] ), 
	.C(\ram[17][15] ), 
	.B(\ram[18][15] ), 
	.A(\ram[16][15] ));
   MUX4EHD U7471 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n6010), 
	.D(n6006), 
	.C(n6008), 
	.B(n6007), 
	.A(n6009));
   MUX4EHD U7472 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n6011), 
	.D(\ram[15][15] ), 
	.C(\ram[13][15] ), 
	.B(\ram[14][15] ), 
	.A(\ram[12][15] ));
   MUX4EHD U7473 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n6012), 
	.D(\ram[11][15] ), 
	.C(\ram[9][15] ), 
	.B(\ram[10][15] ), 
	.A(\ram[8][15] ));
   MUX4EHD U7474 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n6013), 
	.D(\ram[7][15] ), 
	.C(\ram[5][15] ), 
	.B(\ram[6][15] ), 
	.A(\ram[4][15] ));
   MUX4EHD U7475 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n6014), 
	.D(\ram[3][15] ), 
	.C(\ram[1][15] ), 
	.B(\ram[2][15] ), 
	.A(\ram[0][15] ));
   MUX4EHD U7476 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n6015), 
	.D(n6011), 
	.C(n6013), 
	.B(n6012), 
	.A(n6014));
   MUX4EHD U7477 (.S1(n6038), 
	.S0(n7444), 
	.O(n6016), 
	.D(n6000), 
	.C(n6010), 
	.B(n6005), 
	.A(n6015));
   MUX4EHD U7478 (.S1(n6469), 
	.S0(n6470), 
	.O(N4126), 
	.D(n5953), 
	.C(n5995), 
	.B(n5974), 
	.A(n6016));
endmodule

module alu (
	a, 
	b, 
	alu_control, 
	result, 
	zero);
   input [15:0] a;
   input [15:0] b;
   input [2:0] alu_control;
   output [15:0] result;
   output zero;

   // Internal wires
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N46;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N90;
   wire n10;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;

   OR3B1EHD U19 (.O(n31), 
	.I2(result[14]), 
	.I1(result[13]), 
	.B1(n44));
   NR6EHD U69 (.O(zero), 
	.I6(result[0]), 
	.I5(result[10]), 
	.I4(result[11]), 
	.I3(result[12]), 
	.I2(n31), 
	.I1(n74));
   NR8EHD U70 (.O(n49), 
	.I8(result[9]), 
	.I7(result[8]), 
	.I6(result[7]), 
	.I5(result[6]), 
	.I4(result[5]), 
	.I3(result[4]), 
	.I2(result[3]), 
	.I1(result[2]));
   alu_DW01_sub_0 sub_14 (.A({ a[15],
		a[14],
		a[13],
		a[12],
		a[11],
		a[10],
		a[9],
		a[8],
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }), 
	.B({ b[15],
		b[14],
		b[13],
		b[12],
		b[11],
		b[10],
		b[9],
		b[8],
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }), 
	.CI(n10), 
	.DIFF({ N57,
		N56,
		N55,
		N54,
		N53,
		N52,
		N51,
		N50,
		N49,
		N48,
		N47,
		N46,
		N45,
		N44,
		N43,
		N42 }));
   alu_DW01_add_0 r53 (.A({ a[15],
		a[14],
		a[13],
		a[12],
		a[11],
		a[10],
		a[9],
		a[8],
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }), 
	.B({ b[15],
		b[14],
		b[13],
		b[12],
		b[11],
		b[10],
		b[9],
		b[8],
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }), 
	.CI(n10), 
	.SUM({ N41,
		N40,
		N39,
		N38,
		N37,
		N36,
		N35,
		N34,
		N33,
		N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26 }));
   XNR2EHD U2 (.O(n35), 
	.I2(n37), 
	.I1(n80));
   INVDHD U3 (.O(n79), 
	.I(n32));
   NR2CHD U4 (.O(n44), 
	.I2(result[15]), 
	.I1(result[1]));
   AO2222EHD U5 (.O(result[9]), 
	.D2(n50), 
	.D1(b[9]), 
	.C2(n35), 
	.C1(N35), 
	.B2(a[9]), 
	.B1(n79), 
	.A2(n40), 
	.A1(N51));
   OAI12CHD U6 (.O(n50), 
	.B2(n64), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U7 (.O(result[15]), 
	.D2(n45), 
	.D1(b[15]), 
	.C2(n35), 
	.C1(N41), 
	.B2(n79), 
	.B1(a[15]), 
	.A2(n40), 
	.A1(N57));
   OAI12CHD U8 (.O(n45), 
	.B2(n73), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U9 (.O(result[13]), 
	.D2(n48), 
	.D1(b[13]), 
	.C2(n35), 
	.C1(N39), 
	.B2(n79), 
	.B1(a[13]), 
	.A2(n40), 
	.A1(N55));
   OAI12CHD U10 (.O(n48), 
	.B2(n70), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U11 (.O(result[11]), 
	.D2(n42), 
	.D1(b[11]), 
	.C2(n35), 
	.C1(N37), 
	.B2(n79), 
	.B1(a[11]), 
	.A2(n40), 
	.A1(N53));
   OAI12CHD U12 (.O(n42), 
	.B2(n67), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U13 (.O(result[14]), 
	.D2(n47), 
	.D1(b[14]), 
	.C2(n35), 
	.C1(N40), 
	.B2(n79), 
	.B1(a[14]), 
	.A2(n40), 
	.A1(N56));
   OAI12CHD U14 (.O(n47), 
	.B2(n75), 
	.B1(n39), 
	.A1(n32));
   INVDHD U15 (.O(n75), 
	.I(a[14]));
   AO2222CHD U16 (.O(result[12]), 
	.D2(n43), 
	.D1(b[12]), 
	.C2(n35), 
	.C1(N38), 
	.B2(n79), 
	.B1(a[12]), 
	.A2(n40), 
	.A1(N54));
   OAI12CHD U17 (.O(n43), 
	.B2(n69), 
	.B1(n39), 
	.A1(n32));
   INVDHD U18 (.O(n29), 
	.I(b[4]));
   INVDHD U20 (.O(n30), 
	.I(a[4]));
   INVDHD U21 (.O(n59), 
	.I(b[6]));
   INVDHD U22 (.O(n60), 
	.I(a[6]));
   INVDHD U23 (.O(n62), 
	.I(b[8]));
   INVDHD U24 (.O(n63), 
	.I(a[8]));
   INVDHD U25 (.O(n65), 
	.I(b[10]));
   INVDHD U26 (.O(n66), 
	.I(a[10]));
   INVDHD U27 (.O(n68), 
	.I(b[12]));
   INVDHD U28 (.O(n69), 
	.I(a[12]));
   INVDHD U29 (.O(n27), 
	.I(b[2]));
   INVDHD U30 (.O(n26), 
	.I(b[1]));
   INVDHD U31 (.O(n71), 
	.I(b[14]));
   AN2EHD U32 (.O(n36), 
	.I2(alu_control[2]), 
	.I1(N90));
   INVDHD U33 (.O(n72), 
	.I(b[15]));
   OAI112BHD U34 (.O(result[0]), 
	.C2(n78), 
	.C1(n32), 
	.B1(n34), 
	.A1(n33));
   ND2DHD U35 (.O(n33), 
	.I2(n40), 
	.I1(N42));
   AOI222BHD U36 (.O(n34), 
	.C2(n38), 
	.C1(b[0]), 
	.B2(n37), 
	.B1(n36), 
	.A2(n35), 
	.A1(N26));
   OAI12CHD U37 (.O(n38), 
	.B2(n78), 
	.B1(n39), 
	.A1(n32));
   AO2222EHD U38 (.O(result[8]), 
	.D2(n51), 
	.D1(b[8]), 
	.C2(n35), 
	.C1(N34), 
	.B2(n79), 
	.B1(a[8]), 
	.A2(n40), 
	.A1(N50));
   OAI12CHD U39 (.O(n51), 
	.B2(n63), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U40 (.O(result[10]), 
	.D2(n41), 
	.D1(b[10]), 
	.C2(n35), 
	.C1(N36), 
	.B2(n79), 
	.B1(a[10]), 
	.A2(n40), 
	.A1(N52));
   OAI12CHD U41 (.O(n41), 
	.B2(n66), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U42 (.O(result[7]), 
	.D2(n52), 
	.D1(b[7]), 
	.C2(n35), 
	.C1(N33), 
	.B2(n79), 
	.B1(a[7]), 
	.A2(n40), 
	.A1(N49));
   OAI12CHD U43 (.O(n52), 
	.B2(n61), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U44 (.O(result[6]), 
	.D2(n53), 
	.D1(b[6]), 
	.C2(n35), 
	.C1(N32), 
	.B2(n79), 
	.B1(a[6]), 
	.A2(n40), 
	.A1(N48));
   OAI12CHD U45 (.O(n53), 
	.B2(n60), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U46 (.O(result[1]), 
	.D2(n46), 
	.D1(b[1]), 
	.C2(n35), 
	.C1(N27), 
	.B2(n79), 
	.B1(a[1]), 
	.A2(n40), 
	.A1(N43));
   OAI12CHD U47 (.O(n46), 
	.B2(n77), 
	.B1(n39), 
	.A1(n32));
   INVDHD U48 (.O(n77), 
	.I(a[1]));
   ND3CHD U49 (.O(n32), 
	.I3(alu_control[0]), 
	.I2(n80), 
	.I1(alu_control[1]));
   AO2222CHD U50 (.O(result[5]), 
	.D2(n54), 
	.D1(b[5]), 
	.C2(n35), 
	.C1(N31), 
	.B2(n79), 
	.B1(a[5]), 
	.A2(n40), 
	.A1(N47));
   OAI12CHD U51 (.O(n54), 
	.B2(n58), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U52 (.O(result[3]), 
	.D2(n56), 
	.D1(b[3]), 
	.C2(n35), 
	.C1(N29), 
	.B2(n79), 
	.B1(a[3]), 
	.A2(n40), 
	.A1(N45));
   OAI12CHD U53 (.O(n56), 
	.B2(n28), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U54 (.O(result[4]), 
	.D2(n55), 
	.D1(b[4]), 
	.C2(n35), 
	.C1(N30), 
	.B2(n79), 
	.B1(a[4]), 
	.A2(n40), 
	.A1(N46));
   OAI12CHD U55 (.O(n55), 
	.B2(n30), 
	.B1(n39), 
	.A1(n32));
   ND2DHD U56 (.O(n39), 
	.I2(n80), 
	.I1(alu_control[1]));
   NR2CHD U57 (.O(n37), 
	.I2(alu_control[0]), 
	.I1(alu_control[1]));
   INVDHD U58 (.O(n80), 
	.I(alu_control[2]));
   AN3B2BHD U60 (.O(n40), 
	.I1(alu_control[0]), 
	.B2(alu_control[2]), 
	.B1(alu_control[1]));
   AO2222CHD U61 (.O(result[2]), 
	.D2(n57), 
	.D1(b[2]), 
	.C2(n35), 
	.C1(N28), 
	.B2(n79), 
	.B1(a[2]), 
	.A2(n40), 
	.A1(N44));
   OAI12CHD U62 (.O(n57), 
	.B2(n76), 
	.B1(n39), 
	.A1(n32));
   INVDHD U63 (.O(n76), 
	.I(a[2]));
   INVDHD U64 (.O(n74), 
	.I(n49));
   INVDHD U65 (.O(n28), 
	.I(a[3]));
   INVDHD U66 (.O(n58), 
	.I(a[5]));
   INVDHD U67 (.O(n64), 
	.I(a[9]));
   INVDHD U68 (.O(n61), 
	.I(a[7]));
   INVDHD U71 (.O(n67), 
	.I(a[11]));
   INVDHD U72 (.O(n70), 
	.I(a[13]));
   INVDHD U73 (.O(n78), 
	.I(a[0]));
   INVDHD U74 (.O(n73), 
	.I(a[15]));
   TIE0DHD U75 (.O(n10));
   AN2CHD U76 (.O(n22), 
	.I2(b[13]), 
	.I1(n70));
   AN2CHD U77 (.O(n19), 
	.I2(b[11]), 
	.I1(n67));
   AN2CHD U78 (.O(n16), 
	.I2(b[9]), 
	.I1(n64));
   AN2CHD U79 (.O(n13), 
	.I2(b[7]), 
	.I1(n61));
   AN2CHD U80 (.O(n9), 
	.I2(b[5]), 
	.I1(n58));
   AN2CHD U81 (.O(n6), 
	.I2(b[3]), 
	.I1(n28));
   OR2B1CHD U82 (.O(n3), 
	.I1(a[0]), 
	.B1(b[0]));
   OR2CHD U83 (.O(n2), 
	.I2(n3), 
	.I1(a[1]));
   AO222CHD U84 (.O(n4), 
	.C2(a[2]), 
	.C1(n27), 
	.B2(n2), 
	.B1(n26), 
	.A2(a[1]), 
	.A1(n3));
   OAI12CHD U85 (.O(n5), 
	.B2(n27), 
	.B1(a[2]), 
	.A1(n4));
   OAI222BHD U86 (.O(n7), 
	.C2(n30), 
	.C1(b[4]), 
	.B2(n5), 
	.B1(n6), 
	.A2(n28), 
	.A1(b[3]));
   OAI12CHD U87 (.O(n8), 
	.B2(n29), 
	.B1(a[4]), 
	.A1(n7));
   OAI222BHD U88 (.O(n11), 
	.C2(n60), 
	.C1(b[6]), 
	.B2(n8), 
	.B1(n9), 
	.A2(n58), 
	.A1(b[5]));
   OAI12CHD U89 (.O(n12), 
	.B2(n59), 
	.B1(a[6]), 
	.A1(n11));
   OAI222BHD U90 (.O(n14), 
	.C2(n63), 
	.C1(b[8]), 
	.B2(n12), 
	.B1(n13), 
	.A2(n61), 
	.A1(b[7]));
   OAI12CHD U91 (.O(n15), 
	.B2(n62), 
	.B1(a[8]), 
	.A1(n14));
   OAI222BHD U92 (.O(n17), 
	.C2(n64), 
	.C1(b[9]), 
	.B2(n15), 
	.B1(n16), 
	.A2(n66), 
	.A1(b[10]));
   OAI12CHD U93 (.O(n18), 
	.B2(n65), 
	.B1(a[10]), 
	.A1(n17));
   OAI222BHD U94 (.O(n20), 
	.C2(n69), 
	.C1(b[12]), 
	.B2(n18), 
	.B1(n19), 
	.A2(n67), 
	.A1(b[11]));
   OAI12CHD U95 (.O(n21), 
	.B2(n68), 
	.B1(a[12]), 
	.A1(n20));
   OAI222BHD U96 (.O(n23), 
	.C2(n75), 
	.C1(b[14]), 
	.B2(n21), 
	.B1(n22), 
	.A2(n70), 
	.A1(b[13]));
   OAI12CHD U97 (.O(n24), 
	.B2(n71), 
	.B1(a[14]), 
	.A1(n23));
   OAI12CHD U98 (.O(n25), 
	.B2(n73), 
	.B1(b[15]), 
	.A1(n24));
   OAI12CHD U99 (.O(N90), 
	.B2(n72), 
	.B1(a[15]), 
	.A1(n25));
endmodule

module ALUControl (
	ALU_Control, 
	ALUOp, 
	Function);
   output [2:0] ALU_Control;
   input [1:0] ALUOp;
   input [3:0] Function;

   // Internal wires
   wire N9;
   wire N15;
   wire N20;
   wire n3;
   wire n4;
   wire n5;
   wire n1;
   wire n2;

   assign ALU_Control[2] = N9 ;
   assign ALU_Control[1] = N15 ;
   assign ALU_Control[0] = N20 ;

   OAI22CHD U8 (.O(N20), 
	.B2(n2), 
	.B1(n5), 
	.A2(n1), 
	.A1(ALUOp[1]));
   INVDHD U1 (.O(n1), 
	.I(ALUOp[0]));
   AN3B2BHD U2 (.O(N15), 
	.I1(Function[1]), 
	.B2(n5), 
	.B1(ALUOp[0]));
   NR2CHD U3 (.O(N9), 
	.I2(n3), 
	.I1(ALUOp[0]));
   AOI13BHD U4 (.O(n3), 
	.B3(n4), 
	.B2(n2), 
	.B1(Function[2]), 
	.A1(ALUOp[1]));
   NR2CHD U5 (.O(n4), 
	.I2(Function[1]), 
	.I1(Function[3]));
   OR3EHD U6 (.O(n5), 
	.I3(ALUOp[1]), 
	.I2(Function[3]), 
	.I1(Function[2]));
   INVDHD U7 (.O(n2), 
	.I(Function[0]));
endmodule

module JR_Control (
	alu_op, 
	funct, 
	JRControl);
   input [1:0] alu_op;
   input [3:0] funct;
   output JRControl;

   // Internal wires
   wire n1;

   NR6EHD U2 (.O(JRControl), 
	.I6(alu_op[0]), 
	.I5(alu_op[1]), 
	.I4(n1), 
	.I3(funct[1]), 
	.I2(funct[2]), 
	.I1(funct[0]));
   INVDHD U1 (.O(n1), 
	.I(funct[3]));
endmodule

module register_file (
	clk, 
	rst, 
	reg_write_en, 
	reg_write_dest, 
	reg_write_data, 
	reg_read_addr_1, 
	reg_read_data_1, 
	reg_read_addr_2, 
	reg_read_data_2, 
	clk_m__L3_N123, 
	clk_m__L3_N124, 
	clk_m__L3_N126, 
	clk_m__L3_N154, 
	clk_m__L3_N49, 
	clk_m__L3_N50, 
	clk_m__L3_N51, 
	clk_m__L3_N53, 
	clk_m__L3_N54, 
	clk_m__L3_N80);
   input clk;
   input rst;
   input reg_write_en;
   input [2:0] reg_write_dest;
   input [15:0] reg_write_data;
   input [2:0] reg_read_addr_1;
   output [15:0] reg_read_data_1;
   input [2:0] reg_read_addr_2;
   output [15:0] reg_read_data_2;
   input clk_m__L3_N123;
   input clk_m__L3_N124;
   input clk_m__L3_N126;
   input clk_m__L3_N154;
   input clk_m__L3_N49;
   input clk_m__L3_N50;
   input clk_m__L3_N51;
   input clk_m__L3_N53;
   input clk_m__L3_N54;
   input clk_m__L3_N80;

   // Internal wires
   wire FE_OFN95_n240;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire \reg_array[7][15] ;
   wire \reg_array[7][14] ;
   wire \reg_array[7][13] ;
   wire \reg_array[7][12] ;
   wire \reg_array[7][11] ;
   wire \reg_array[7][10] ;
   wire \reg_array[7][9] ;
   wire \reg_array[7][8] ;
   wire \reg_array[7][7] ;
   wire \reg_array[7][6] ;
   wire \reg_array[7][5] ;
   wire \reg_array[7][4] ;
   wire \reg_array[7][3] ;
   wire \reg_array[7][2] ;
   wire \reg_array[7][1] ;
   wire \reg_array[7][0] ;
   wire \reg_array[6][15] ;
   wire \reg_array[6][14] ;
   wire \reg_array[6][13] ;
   wire \reg_array[6][12] ;
   wire \reg_array[6][11] ;
   wire \reg_array[6][10] ;
   wire \reg_array[6][9] ;
   wire \reg_array[6][8] ;
   wire \reg_array[6][7] ;
   wire \reg_array[6][6] ;
   wire \reg_array[6][5] ;
   wire \reg_array[6][4] ;
   wire \reg_array[6][3] ;
   wire \reg_array[6][2] ;
   wire \reg_array[6][1] ;
   wire \reg_array[6][0] ;
   wire \reg_array[5][15] ;
   wire \reg_array[5][14] ;
   wire \reg_array[5][13] ;
   wire \reg_array[5][12] ;
   wire \reg_array[5][11] ;
   wire \reg_array[5][10] ;
   wire \reg_array[5][9] ;
   wire \reg_array[5][8] ;
   wire \reg_array[5][7] ;
   wire \reg_array[5][6] ;
   wire \reg_array[5][5] ;
   wire \reg_array[5][4] ;
   wire \reg_array[5][3] ;
   wire \reg_array[5][2] ;
   wire \reg_array[5][1] ;
   wire \reg_array[5][0] ;
   wire \reg_array[4][15] ;
   wire \reg_array[4][14] ;
   wire \reg_array[4][13] ;
   wire \reg_array[4][12] ;
   wire \reg_array[4][11] ;
   wire \reg_array[4][10] ;
   wire \reg_array[4][9] ;
   wire \reg_array[4][8] ;
   wire \reg_array[4][7] ;
   wire \reg_array[4][6] ;
   wire \reg_array[4][5] ;
   wire \reg_array[4][4] ;
   wire \reg_array[4][3] ;
   wire \reg_array[4][2] ;
   wire \reg_array[4][1] ;
   wire \reg_array[4][0] ;
   wire \reg_array[3][15] ;
   wire \reg_array[3][14] ;
   wire \reg_array[3][13] ;
   wire \reg_array[3][12] ;
   wire \reg_array[3][11] ;
   wire \reg_array[3][10] ;
   wire \reg_array[3][9] ;
   wire \reg_array[3][8] ;
   wire \reg_array[3][7] ;
   wire \reg_array[3][6] ;
   wire \reg_array[3][5] ;
   wire \reg_array[3][4] ;
   wire \reg_array[3][3] ;
   wire \reg_array[3][2] ;
   wire \reg_array[3][1] ;
   wire \reg_array[3][0] ;
   wire \reg_array[2][15] ;
   wire \reg_array[2][14] ;
   wire \reg_array[2][13] ;
   wire \reg_array[2][12] ;
   wire \reg_array[2][11] ;
   wire \reg_array[2][10] ;
   wire \reg_array[2][9] ;
   wire \reg_array[2][8] ;
   wire \reg_array[2][7] ;
   wire \reg_array[2][6] ;
   wire \reg_array[2][5] ;
   wire \reg_array[2][4] ;
   wire \reg_array[2][3] ;
   wire \reg_array[2][2] ;
   wire \reg_array[2][1] ;
   wire \reg_array[2][0] ;
   wire \reg_array[1][15] ;
   wire \reg_array[1][14] ;
   wire \reg_array[1][13] ;
   wire \reg_array[1][12] ;
   wire \reg_array[1][11] ;
   wire \reg_array[1][10] ;
   wire \reg_array[1][9] ;
   wire \reg_array[1][8] ;
   wire \reg_array[1][7] ;
   wire \reg_array[1][6] ;
   wire \reg_array[1][5] ;
   wire \reg_array[1][4] ;
   wire \reg_array[1][3] ;
   wire \reg_array[1][2] ;
   wire \reg_array[1][1] ;
   wire \reg_array[1][0] ;
   wire \reg_array[0][15] ;
   wire \reg_array[0][14] ;
   wire \reg_array[0][13] ;
   wire \reg_array[0][12] ;
   wire \reg_array[0][11] ;
   wire \reg_array[0][10] ;
   wire \reg_array[0][9] ;
   wire \reg_array[0][8] ;
   wire \reg_array[0][7] ;
   wire \reg_array[0][6] ;
   wire \reg_array[0][5] ;
   wire \reg_array[0][4] ;
   wire \reg_array[0][3] ;
   wire \reg_array[0][2] ;
   wire \reg_array[0][1] ;
   wire \reg_array[0][0] ;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n238;
   wire n239;
   wire n240;

   assign N18 = reg_read_addr_1[0] ;
   assign N19 = reg_read_addr_1[1] ;
   assign N20 = reg_read_addr_1[2] ;
   assign N21 = reg_read_addr_2[0] ;
   assign N22 = reg_read_addr_2[1] ;
   assign N23 = reg_read_addr_2[2] ;

   BUFGHD FE_OFC95_n240 (.O(FE_OFN95_n240), 
	.I(n240));
   DFERBCHD \reg_array_reg[5][15]  (.RB(n240), 
	.Q(\reg_array[5][15] ), 
	.EB(n144), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[1][15]  (.RB(n240), 
	.Q(\reg_array[1][15] ), 
	.EB(n137), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[1][14]  (.RB(n240), 
	.Q(\reg_array[1][14] ), 
	.EB(n137), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[6][15]  (.RB(n240), 
	.Q(\reg_array[6][15] ), 
	.EB(n146), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[6][14]  (.RB(n240), 
	.Q(\reg_array[6][14] ), 
	.EB(n146), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[2][15]  (.RB(n240), 
	.Q(\reg_array[2][15] ), 
	.EB(n138), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[2][14]  (.RB(n240), 
	.Q(\reg_array[2][14] ), 
	.EB(n138), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[4][15]  (.RB(n240), 
	.Q(\reg_array[4][15] ), 
	.EB(n142), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[4][14]  (.RB(n240), 
	.Q(\reg_array[4][14] ), 
	.EB(n142), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[0][15]  (.RB(n240), 
	.Q(\reg_array[0][15] ), 
	.EB(n135), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[0][14]  (.RB(n240), 
	.Q(\reg_array[0][14] ), 
	.EB(n135), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[7][15]  (.RB(n240), 
	.Q(\reg_array[7][15] ), 
	.EB(n148), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[7][14]  (.RB(n240), 
	.Q(\reg_array[7][14] ), 
	.EB(n148), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[3][15]  (.RB(n240), 
	.Q(\reg_array[3][15] ), 
	.EB(n140), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[3][14]  (.RB(n240), 
	.Q(\reg_array[3][14] ), 
	.EB(n140), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[5][14]  (.RB(n240), 
	.Q(\reg_array[5][14] ), 
	.EB(n144), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[5][13]  (.RB(n240), 
	.Q(\reg_array[5][13] ), 
	.EB(n144), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[5][12]  (.RB(n240), 
	.Q(\reg_array[5][12] ), 
	.EB(n144), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[5][11]  (.RB(n240), 
	.Q(\reg_array[5][11] ), 
	.EB(n144), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[5][10]  (.RB(n240), 
	.Q(\reg_array[5][10] ), 
	.EB(n144), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[5][9]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][9] ), 
	.EB(n144), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[1][13]  (.RB(n240), 
	.Q(\reg_array[1][13] ), 
	.EB(n137), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[1][12]  (.RB(n240), 
	.Q(\reg_array[1][12] ), 
	.EB(n137), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[1][11]  (.RB(n240), 
	.Q(\reg_array[1][11] ), 
	.EB(n137), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[1][10]  (.RB(n240), 
	.Q(\reg_array[1][10] ), 
	.EB(n137), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[1][9]  (.RB(n240), 
	.Q(\reg_array[1][9] ), 
	.EB(n137), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[6][13]  (.RB(n240), 
	.Q(\reg_array[6][13] ), 
	.EB(n146), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[6][12]  (.RB(n240), 
	.Q(\reg_array[6][12] ), 
	.EB(n146), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[6][11]  (.RB(n240), 
	.Q(\reg_array[6][11] ), 
	.EB(n146), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[6][10]  (.RB(n240), 
	.Q(\reg_array[6][10] ), 
	.EB(n146), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[6][9]  (.RB(n240), 
	.Q(\reg_array[6][9] ), 
	.EB(n146), 
	.D(reg_write_data[9]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[2][13]  (.RB(n240), 
	.Q(\reg_array[2][13] ), 
	.EB(n138), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[2][12]  (.RB(n240), 
	.Q(\reg_array[2][12] ), 
	.EB(n138), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[2][11]  (.RB(n240), 
	.Q(\reg_array[2][11] ), 
	.EB(n138), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[2][10]  (.RB(n240), 
	.Q(\reg_array[2][10] ), 
	.EB(n138), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[2][9]  (.RB(n240), 
	.Q(\reg_array[2][9] ), 
	.EB(n138), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[4][13]  (.RB(n240), 
	.Q(\reg_array[4][13] ), 
	.EB(n142), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[4][12]  (.RB(n240), 
	.Q(\reg_array[4][12] ), 
	.EB(n142), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[4][11]  (.RB(n240), 
	.Q(\reg_array[4][11] ), 
	.EB(n142), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[4][10]  (.RB(n240), 
	.Q(\reg_array[4][10] ), 
	.EB(n142), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[4][9]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][9] ), 
	.EB(n142), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[0][13]  (.RB(n240), 
	.Q(\reg_array[0][13] ), 
	.EB(n135), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[0][12]  (.RB(n240), 
	.Q(\reg_array[0][12] ), 
	.EB(n135), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[0][11]  (.RB(n240), 
	.Q(\reg_array[0][11] ), 
	.EB(n135), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[0][10]  (.RB(n240), 
	.Q(\reg_array[0][10] ), 
	.EB(n135), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[0][9]  (.RB(n240), 
	.Q(\reg_array[0][9] ), 
	.EB(n135), 
	.D(reg_write_data[9]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[7][13]  (.RB(n240), 
	.Q(\reg_array[7][13] ), 
	.EB(n148), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[7][12]  (.RB(n240), 
	.Q(\reg_array[7][12] ), 
	.EB(n148), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[7][11]  (.RB(n240), 
	.Q(\reg_array[7][11] ), 
	.EB(n148), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[7][10]  (.RB(n240), 
	.Q(\reg_array[7][10] ), 
	.EB(n148), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[7][9]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][9] ), 
	.EB(n148), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[7][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][8] ), 
	.EB(n148), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[3][13]  (.RB(n240), 
	.Q(\reg_array[3][13] ), 
	.EB(n140), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[3][12]  (.RB(n240), 
	.Q(\reg_array[3][12] ), 
	.EB(n140), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[3][11]  (.RB(n240), 
	.Q(\reg_array[3][11] ), 
	.EB(n140), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[3][10]  (.RB(n240), 
	.Q(\reg_array[3][10] ), 
	.EB(n140), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[3][9]  (.RB(n240), 
	.Q(\reg_array[3][9] ), 
	.EB(n140), 
	.D(reg_write_data[9]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[3][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][8] ), 
	.EB(n140), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[5][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][8] ), 
	.EB(n144), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[5][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][7] ), 
	.EB(n144), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[5][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][6] ), 
	.EB(n144), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[5][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][5] ), 
	.EB(n144), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[5][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][4] ), 
	.EB(n144), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[5][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][3] ), 
	.EB(n144), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[1][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][8] ), 
	.EB(n137), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[1][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][7] ), 
	.EB(n137), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[1][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][6] ), 
	.EB(n137), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[1][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][5] ), 
	.EB(n137), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[1][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][4] ), 
	.EB(n137), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[1][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][3] ), 
	.EB(n137), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[6][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][8] ), 
	.EB(n146), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[6][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][7] ), 
	.EB(n146), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[6][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][6] ), 
	.EB(n146), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[6][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][5] ), 
	.EB(n146), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[6][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][4] ), 
	.EB(n146), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[6][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][3] ), 
	.EB(n146), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[2][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][8] ), 
	.EB(n138), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[2][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][7] ), 
	.EB(n138), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[2][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][6] ), 
	.EB(n138), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[2][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][5] ), 
	.EB(n138), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[2][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][4] ), 
	.EB(n138), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[2][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][3] ), 
	.EB(n138), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[4][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][8] ), 
	.EB(n142), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[4][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][7] ), 
	.EB(n142), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[4][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][6] ), 
	.EB(n142), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[4][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][5] ), 
	.EB(n142), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[4][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][4] ), 
	.EB(n142), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[4][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][3] ), 
	.EB(n142), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][8] ), 
	.EB(n135), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[0][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][7] ), 
	.EB(n135), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[0][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][6] ), 
	.EB(n135), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[0][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][5] ), 
	.EB(n135), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[0][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][4] ), 
	.EB(n135), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][3] ), 
	.EB(n135), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[7][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][7] ), 
	.EB(n148), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[7][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][6] ), 
	.EB(n148), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[7][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][5] ), 
	.EB(n148), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[7][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][4] ), 
	.EB(n148), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[7][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][3] ), 
	.EB(n148), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[3][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][7] ), 
	.EB(n140), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][6] ), 
	.EB(n140), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][5] ), 
	.EB(n140), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][4] ), 
	.EB(n140), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][3] ), 
	.EB(n140), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N54));
   DFERBCHD \reg_array_reg[5][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][2] ), 
	.EB(n144), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[5][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][1] ), 
	.EB(n144), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[5][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][0] ), 
	.EB(n144), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[1][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][2] ), 
	.EB(n137), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[1][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][1] ), 
	.EB(n137), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[1][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][0] ), 
	.EB(n137), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[6][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][2] ), 
	.EB(n146), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[6][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][1] ), 
	.EB(n146), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[6][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][0] ), 
	.EB(n146), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[2][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][2] ), 
	.EB(n138), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[2][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][1] ), 
	.EB(n138), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[2][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][0] ), 
	.EB(n138), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[4][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][2] ), 
	.EB(n142), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N80));
   DFERBCHD \reg_array_reg[4][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][1] ), 
	.EB(n142), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[4][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][0] ), 
	.EB(n142), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[0][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][2] ), 
	.EB(n135), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][1] ), 
	.EB(n135), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][0] ), 
	.EB(n135), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[7][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][2] ), 
	.EB(n148), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[7][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][1] ), 
	.EB(n148), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N80));
   DFERBCHD \reg_array_reg[7][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][0] ), 
	.EB(n148), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[3][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][2] ), 
	.EB(n140), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[3][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][1] ), 
	.EB(n140), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[3][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][0] ), 
	.EB(n140), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   NR2CHD U2 (.O(n136), 
	.I2(reg_write_dest[1]), 
	.I1(reg_write_dest[2]));
   INVDHD U3 (.O(n239), 
	.I(reg_write_dest[0]));
   ND3CHD U17 (.O(n140), 
	.I3(n141), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[1]));
   NR2CHD U18 (.O(n141), 
	.I2(n238), 
	.I1(reg_write_dest[2]));
   ND3CHD U20 (.O(n144), 
	.I3(n145), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[2]));
   NR2CHD U21 (.O(n145), 
	.I2(n238), 
	.I1(reg_write_dest[1]));
   ND3CHD U23 (.O(n146), 
	.I3(n147), 
	.I2(reg_write_dest[1]), 
	.I1(reg_write_dest[2]));
   NR2CHD U24 (.O(n147), 
	.I2(n238), 
	.I1(reg_write_dest[0]));
   ND3CHD U26 (.O(n148), 
	.I3(n149), 
	.I2(reg_write_dest[1]), 
	.I1(reg_write_dest[2]));
   NR2CHD U27 (.O(n149), 
	.I2(n239), 
	.I1(n238));
   INVDHD U34 (.O(n238), 
	.I(reg_write_en));
   ND3CHD U36 (.O(n137), 
	.I3(n136), 
	.I2(reg_write_en), 
	.I1(reg_write_dest[0]));
   ND3CHD U38 (.O(n138), 
	.I3(n139), 
	.I2(reg_write_en), 
	.I1(reg_write_dest[1]));
   NR2CHD U39 (.O(n139), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[2]));
   ND3CHD U41 (.O(n142), 
	.I3(n143), 
	.I2(reg_write_en), 
	.I1(reg_write_dest[2]));
   NR2CHD U42 (.O(n143), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[1]));
   ND3CHD U44 (.O(n135), 
	.I3(n136), 
	.I2(n239), 
	.I1(reg_write_en));
   AN2EHD U47 (.O(reg_read_data_1[1]), 
	.I2(n134), 
	.I1(N167));
   MUX2EHD U48 (.S(N20), 
	.O(N167), 
	.B(n131), 
	.A(n132));
   AN2EHD U49 (.O(reg_read_data_2[1]), 
	.I2(n133), 
	.I1(N183));
   MUX2EHD U50 (.S(N23), 
	.O(N183), 
	.B(n180), 
	.A(n181));
   AN2EHD U51 (.O(reg_read_data_2[2]), 
	.I2(n133), 
	.I1(N182));
   MUX2EHD U52 (.S(N23), 
	.O(N182), 
	.B(n182), 
	.A(n183));
   AN2EHD U53 (.O(reg_read_data_2[0]), 
	.I2(n133), 
	.I1(N184));
   MUX2EHD U54 (.S(N23), 
	.O(N184), 
	.B(n178), 
	.A(n179));
   AN2EHD U55 (.O(reg_read_data_1[0]), 
	.I2(n134), 
	.I1(N168));
   MUX2EHD U56 (.S(N20), 
	.O(N168), 
	.B(n129), 
	.A(n130));
   AN2EHD U57 (.O(reg_read_data_2[7]), 
	.I2(n133), 
	.I1(N177));
   MUX2EHD U58 (.S(N23), 
	.O(N177), 
	.B(n192), 
	.A(n193));
   AN2EHD U59 (.O(reg_read_data_2[8]), 
	.I2(n133), 
	.I1(N176));
   MUX2EHD U60 (.S(N23), 
	.O(N176), 
	.B(n194), 
	.A(n195));
   AN2EHD U61 (.O(reg_read_data_2[3]), 
	.I2(n133), 
	.I1(N181));
   MUX2EHD U62 (.S(N23), 
	.O(N181), 
	.B(n184), 
	.A(n185));
   AN2EHD U63 (.O(reg_read_data_2[4]), 
	.I2(n133), 
	.I1(N180));
   MUX2EHD U64 (.S(N23), 
	.O(N180), 
	.B(n186), 
	.A(n187));
   AN2EHD U65 (.O(reg_read_data_2[5]), 
	.I2(n133), 
	.I1(N179));
   MUX2EHD U66 (.S(N23), 
	.O(N179), 
	.B(n188), 
	.A(n189));
   AN2EHD U67 (.O(reg_read_data_2[6]), 
	.I2(n133), 
	.I1(N178));
   MUX2EHD U68 (.S(N23), 
	.O(N178), 
	.B(n190), 
	.A(n191));
   AN2EHD U69 (.O(reg_read_data_1[2]), 
	.I2(n134), 
	.I1(N166));
   MUX2EHD U70 (.S(N20), 
	.O(N166), 
	.B(n150), 
	.A(n151));
   AN2EHD U71 (.O(reg_read_data_1[3]), 
	.I2(n134), 
	.I1(N165));
   MUX2EHD U72 (.S(N20), 
	.O(N165), 
	.B(n152), 
	.A(n153));
   AN2EHD U73 (.O(reg_read_data_1[4]), 
	.I2(n134), 
	.I1(N164));
   MUX2EHD U74 (.S(N20), 
	.O(N164), 
	.B(n154), 
	.A(n155));
   AN2EHD U75 (.O(reg_read_data_1[5]), 
	.I2(n134), 
	.I1(N163));
   MUX2EHD U76 (.S(N20), 
	.O(N163), 
	.B(n156), 
	.A(n157));
   AN2EHD U77 (.O(reg_read_data_1[6]), 
	.I2(n134), 
	.I1(N162));
   MUX2EHD U78 (.S(N20), 
	.O(N162), 
	.B(n158), 
	.A(n159));
   AN2EHD U79 (.O(reg_read_data_1[7]), 
	.I2(n134), 
	.I1(N161));
   MUX2EHD U80 (.S(N20), 
	.O(N161), 
	.B(n160), 
	.A(n161));
   AN2EHD U81 (.O(reg_read_data_1[9]), 
	.I2(n134), 
	.I1(N159));
   MUX2EHD U82 (.S(N20), 
	.O(N159), 
	.B(n164), 
	.A(n165));
   AN2EHD U83 (.O(reg_read_data_1[13]), 
	.I2(n134), 
	.I1(N155));
   MUX2EHD U84 (.S(N20), 
	.O(N155), 
	.B(n172), 
	.A(n173));
   AN2EHD U85 (.O(reg_read_data_2[9]), 
	.I2(n133), 
	.I1(N175));
   MUX2EHD U86 (.S(N23), 
	.O(N175), 
	.B(n196), 
	.A(n197));
   AN2EHD U87 (.O(reg_read_data_2[10]), 
	.I2(n133), 
	.I1(N174));
   MUX2EHD U88 (.S(N23), 
	.O(N174), 
	.B(n198), 
	.A(n199));
   AN2EHD U89 (.O(reg_read_data_2[11]), 
	.I2(n133), 
	.I1(N173));
   MUX2EHD U90 (.S(N23), 
	.O(N173), 
	.B(n200), 
	.A(n201));
   AN2EHD U91 (.O(reg_read_data_2[12]), 
	.I2(n133), 
	.I1(N172));
   MUX2EHD U92 (.S(N23), 
	.O(N172), 
	.B(n202), 
	.A(n203));
   AN2EHD U93 (.O(reg_read_data_2[13]), 
	.I2(n133), 
	.I1(N171));
   MUX2EHD U94 (.S(N23), 
	.O(N171), 
	.B(n204), 
	.A(n205));
   AN2EHD U95 (.O(reg_read_data_2[14]), 
	.I2(n133), 
	.I1(N170));
   MUX2EHD U96 (.S(N23), 
	.O(N170), 
	.B(n206), 
	.A(n207));
   AN2EHD U97 (.O(reg_read_data_1[12]), 
	.I2(n134), 
	.I1(N156));
   MUX2EHD U98 (.S(N20), 
	.O(N156), 
	.B(n170), 
	.A(n171));
   AN2EHD U99 (.O(reg_read_data_1[8]), 
	.I2(n134), 
	.I1(N160));
   MUX2EHD U100 (.S(N20), 
	.O(N160), 
	.B(n162), 
	.A(n163));
   AN2EHD U101 (.O(reg_read_data_1[10]), 
	.I2(n134), 
	.I1(N158));
   MUX2EHD U102 (.S(N20), 
	.O(N158), 
	.B(n166), 
	.A(n167));
   AN2EHD U103 (.O(reg_read_data_1[11]), 
	.I2(n134), 
	.I1(N157));
   MUX2EHD U104 (.S(N20), 
	.O(N157), 
	.B(n168), 
	.A(n169));
   AN2EHD U105 (.O(reg_read_data_1[15]), 
	.I2(n134), 
	.I1(N153));
   MUX2EHD U106 (.S(N20), 
	.O(N153), 
	.B(n176), 
	.A(n177));
   AN2EHD U107 (.O(reg_read_data_2[15]), 
	.I2(n133), 
	.I1(N169));
   MUX2EHD U108 (.S(N23), 
	.O(N169), 
	.B(n208), 
	.A(n209));
   AN2EHD U109 (.O(reg_read_data_1[14]), 
	.I2(n134), 
	.I1(N154));
   MUX2EHD U110 (.S(N20), 
	.O(N154), 
	.B(n174), 
	.A(n175));
   INVDHD U111 (.O(n240), 
	.I(rst));
   OR3EHD U112 (.O(n133), 
	.I3(N21), 
	.I2(N23), 
	.I1(N22));
   OR3EHD U113 (.O(n134), 
	.I3(N18), 
	.I2(N20), 
	.I1(N19));
   MUX4EHD U114 (.S1(N18), 
	.S0(N19), 
	.O(n129), 
	.D(\reg_array[7][0] ), 
	.C(\reg_array[5][0] ), 
	.B(\reg_array[6][0] ), 
	.A(\reg_array[4][0] ));
   MUX4EHD U115 (.S1(N18), 
	.S0(N19), 
	.O(n130), 
	.D(\reg_array[3][0] ), 
	.C(\reg_array[1][0] ), 
	.B(\reg_array[2][0] ), 
	.A(\reg_array[0][0] ));
   MUX4EHD U116 (.S1(N18), 
	.S0(N19), 
	.O(n131), 
	.D(\reg_array[7][1] ), 
	.C(\reg_array[5][1] ), 
	.B(\reg_array[6][1] ), 
	.A(\reg_array[4][1] ));
   MUX4EHD U117 (.S1(N18), 
	.S0(N19), 
	.O(n132), 
	.D(\reg_array[3][1] ), 
	.C(\reg_array[1][1] ), 
	.B(\reg_array[2][1] ), 
	.A(\reg_array[0][1] ));
   MUX4EHD U118 (.S1(N18), 
	.S0(N19), 
	.O(n150), 
	.D(\reg_array[7][2] ), 
	.C(\reg_array[5][2] ), 
	.B(\reg_array[6][2] ), 
	.A(\reg_array[4][2] ));
   MUX4EHD U119 (.S1(N18), 
	.S0(N19), 
	.O(n151), 
	.D(\reg_array[3][2] ), 
	.C(\reg_array[1][2] ), 
	.B(\reg_array[2][2] ), 
	.A(\reg_array[0][2] ));
   MUX4EHD U120 (.S1(N18), 
	.S0(N19), 
	.O(n152), 
	.D(\reg_array[7][3] ), 
	.C(\reg_array[5][3] ), 
	.B(\reg_array[6][3] ), 
	.A(\reg_array[4][3] ));
   MUX4EHD U121 (.S1(N18), 
	.S0(N19), 
	.O(n153), 
	.D(\reg_array[3][3] ), 
	.C(\reg_array[1][3] ), 
	.B(\reg_array[2][3] ), 
	.A(\reg_array[0][3] ));
   MUX4EHD U122 (.S1(N18), 
	.S0(N19), 
	.O(n154), 
	.D(\reg_array[7][4] ), 
	.C(\reg_array[5][4] ), 
	.B(\reg_array[6][4] ), 
	.A(\reg_array[4][4] ));
   MUX4EHD U123 (.S1(N18), 
	.S0(N19), 
	.O(n155), 
	.D(\reg_array[3][4] ), 
	.C(\reg_array[1][4] ), 
	.B(\reg_array[2][4] ), 
	.A(\reg_array[0][4] ));
   MUX4EHD U124 (.S1(N18), 
	.S0(N19), 
	.O(n156), 
	.D(\reg_array[7][5] ), 
	.C(\reg_array[5][5] ), 
	.B(\reg_array[6][5] ), 
	.A(\reg_array[4][5] ));
   MUX4EHD U125 (.S1(N18), 
	.S0(N19), 
	.O(n157), 
	.D(\reg_array[3][5] ), 
	.C(\reg_array[1][5] ), 
	.B(\reg_array[2][5] ), 
	.A(\reg_array[0][5] ));
   MUX4EHD U126 (.S1(N18), 
	.S0(N19), 
	.O(n158), 
	.D(\reg_array[7][6] ), 
	.C(\reg_array[5][6] ), 
	.B(\reg_array[6][6] ), 
	.A(\reg_array[4][6] ));
   MUX4EHD U127 (.S1(N18), 
	.S0(N19), 
	.O(n159), 
	.D(\reg_array[3][6] ), 
	.C(\reg_array[1][6] ), 
	.B(\reg_array[2][6] ), 
	.A(\reg_array[0][6] ));
   MUX4EHD U128 (.S1(N18), 
	.S0(N19), 
	.O(n160), 
	.D(\reg_array[7][7] ), 
	.C(\reg_array[5][7] ), 
	.B(\reg_array[6][7] ), 
	.A(\reg_array[4][7] ));
   MUX4EHD U129 (.S1(N18), 
	.S0(N19), 
	.O(n161), 
	.D(\reg_array[3][7] ), 
	.C(\reg_array[1][7] ), 
	.B(\reg_array[2][7] ), 
	.A(\reg_array[0][7] ));
   MUX4EHD U130 (.S1(N18), 
	.S0(N19), 
	.O(n162), 
	.D(\reg_array[7][8] ), 
	.C(\reg_array[5][8] ), 
	.B(\reg_array[6][8] ), 
	.A(\reg_array[4][8] ));
   MUX4EHD U131 (.S1(N18), 
	.S0(N19), 
	.O(n163), 
	.D(\reg_array[3][8] ), 
	.C(\reg_array[1][8] ), 
	.B(\reg_array[2][8] ), 
	.A(\reg_array[0][8] ));
   MUX4EHD U132 (.S1(N18), 
	.S0(N19), 
	.O(n164), 
	.D(\reg_array[7][9] ), 
	.C(\reg_array[5][9] ), 
	.B(\reg_array[6][9] ), 
	.A(\reg_array[4][9] ));
   MUX4EHD U133 (.S1(N18), 
	.S0(N19), 
	.O(n165), 
	.D(\reg_array[3][9] ), 
	.C(\reg_array[1][9] ), 
	.B(\reg_array[2][9] ), 
	.A(\reg_array[0][9] ));
   MUX4EHD U134 (.S1(N18), 
	.S0(N19), 
	.O(n166), 
	.D(\reg_array[7][10] ), 
	.C(\reg_array[5][10] ), 
	.B(\reg_array[6][10] ), 
	.A(\reg_array[4][10] ));
   MUX4EHD U135 (.S1(N18), 
	.S0(N19), 
	.O(n167), 
	.D(\reg_array[3][10] ), 
	.C(\reg_array[1][10] ), 
	.B(\reg_array[2][10] ), 
	.A(\reg_array[0][10] ));
   MUX4EHD U136 (.S1(N18), 
	.S0(N19), 
	.O(n168), 
	.D(\reg_array[7][11] ), 
	.C(\reg_array[5][11] ), 
	.B(\reg_array[6][11] ), 
	.A(\reg_array[4][11] ));
   MUX4EHD U137 (.S1(N18), 
	.S0(N19), 
	.O(n169), 
	.D(\reg_array[3][11] ), 
	.C(\reg_array[1][11] ), 
	.B(\reg_array[2][11] ), 
	.A(\reg_array[0][11] ));
   MUX4EHD U138 (.S1(N18), 
	.S0(N19), 
	.O(n170), 
	.D(\reg_array[7][12] ), 
	.C(\reg_array[5][12] ), 
	.B(\reg_array[6][12] ), 
	.A(\reg_array[4][12] ));
   MUX4EHD U139 (.S1(N18), 
	.S0(N19), 
	.O(n171), 
	.D(\reg_array[3][12] ), 
	.C(\reg_array[1][12] ), 
	.B(\reg_array[2][12] ), 
	.A(\reg_array[0][12] ));
   MUX4EHD U140 (.S1(N18), 
	.S0(N19), 
	.O(n172), 
	.D(\reg_array[7][13] ), 
	.C(\reg_array[5][13] ), 
	.B(\reg_array[6][13] ), 
	.A(\reg_array[4][13] ));
   MUX4EHD U141 (.S1(N18), 
	.S0(N19), 
	.O(n173), 
	.D(\reg_array[3][13] ), 
	.C(\reg_array[1][13] ), 
	.B(\reg_array[2][13] ), 
	.A(\reg_array[0][13] ));
   MUX4EHD U142 (.S1(N18), 
	.S0(N19), 
	.O(n174), 
	.D(\reg_array[7][14] ), 
	.C(\reg_array[5][14] ), 
	.B(\reg_array[6][14] ), 
	.A(\reg_array[4][14] ));
   MUX4EHD U143 (.S1(N18), 
	.S0(N19), 
	.O(n175), 
	.D(\reg_array[3][14] ), 
	.C(\reg_array[1][14] ), 
	.B(\reg_array[2][14] ), 
	.A(\reg_array[0][14] ));
   MUX4EHD U144 (.S1(N18), 
	.S0(N19), 
	.O(n176), 
	.D(\reg_array[7][15] ), 
	.C(\reg_array[5][15] ), 
	.B(\reg_array[6][15] ), 
	.A(\reg_array[4][15] ));
   MUX4EHD U145 (.S1(N18), 
	.S0(N19), 
	.O(n177), 
	.D(\reg_array[3][15] ), 
	.C(\reg_array[1][15] ), 
	.B(\reg_array[2][15] ), 
	.A(\reg_array[0][15] ));
   MUX4EHD U146 (.S1(N21), 
	.S0(N22), 
	.O(n178), 
	.D(\reg_array[7][0] ), 
	.C(\reg_array[5][0] ), 
	.B(\reg_array[6][0] ), 
	.A(\reg_array[4][0] ));
   MUX4EHD U147 (.S1(N21), 
	.S0(N22), 
	.O(n179), 
	.D(\reg_array[3][0] ), 
	.C(\reg_array[1][0] ), 
	.B(\reg_array[2][0] ), 
	.A(\reg_array[0][0] ));
   MUX4EHD U148 (.S1(N21), 
	.S0(N22), 
	.O(n180), 
	.D(\reg_array[7][1] ), 
	.C(\reg_array[5][1] ), 
	.B(\reg_array[6][1] ), 
	.A(\reg_array[4][1] ));
   MUX4EHD U149 (.S1(N21), 
	.S0(N22), 
	.O(n181), 
	.D(\reg_array[3][1] ), 
	.C(\reg_array[1][1] ), 
	.B(\reg_array[2][1] ), 
	.A(\reg_array[0][1] ));
   MUX4EHD U150 (.S1(N21), 
	.S0(N22), 
	.O(n182), 
	.D(\reg_array[7][2] ), 
	.C(\reg_array[5][2] ), 
	.B(\reg_array[6][2] ), 
	.A(\reg_array[4][2] ));
   MUX4EHD U151 (.S1(N21), 
	.S0(N22), 
	.O(n183), 
	.D(\reg_array[3][2] ), 
	.C(\reg_array[1][2] ), 
	.B(\reg_array[2][2] ), 
	.A(\reg_array[0][2] ));
   MUX4EHD U152 (.S1(N21), 
	.S0(N22), 
	.O(n184), 
	.D(\reg_array[7][3] ), 
	.C(\reg_array[5][3] ), 
	.B(\reg_array[6][3] ), 
	.A(\reg_array[4][3] ));
   MUX4EHD U153 (.S1(N21), 
	.S0(N22), 
	.O(n185), 
	.D(\reg_array[3][3] ), 
	.C(\reg_array[1][3] ), 
	.B(\reg_array[2][3] ), 
	.A(\reg_array[0][3] ));
   MUX4EHD U154 (.S1(N21), 
	.S0(N22), 
	.O(n186), 
	.D(\reg_array[7][4] ), 
	.C(\reg_array[5][4] ), 
	.B(\reg_array[6][4] ), 
	.A(\reg_array[4][4] ));
   MUX4EHD U155 (.S1(N21), 
	.S0(N22), 
	.O(n187), 
	.D(\reg_array[3][4] ), 
	.C(\reg_array[1][4] ), 
	.B(\reg_array[2][4] ), 
	.A(\reg_array[0][4] ));
   MUX4EHD U156 (.S1(N21), 
	.S0(N22), 
	.O(n188), 
	.D(\reg_array[7][5] ), 
	.C(\reg_array[5][5] ), 
	.B(\reg_array[6][5] ), 
	.A(\reg_array[4][5] ));
   MUX4EHD U157 (.S1(N21), 
	.S0(N22), 
	.O(n189), 
	.D(\reg_array[3][5] ), 
	.C(\reg_array[1][5] ), 
	.B(\reg_array[2][5] ), 
	.A(\reg_array[0][5] ));
   MUX4EHD U158 (.S1(N21), 
	.S0(N22), 
	.O(n190), 
	.D(\reg_array[7][6] ), 
	.C(\reg_array[5][6] ), 
	.B(\reg_array[6][6] ), 
	.A(\reg_array[4][6] ));
   MUX4EHD U159 (.S1(N21), 
	.S0(N22), 
	.O(n191), 
	.D(\reg_array[3][6] ), 
	.C(\reg_array[1][6] ), 
	.B(\reg_array[2][6] ), 
	.A(\reg_array[0][6] ));
   MUX4EHD U160 (.S1(N21), 
	.S0(N22), 
	.O(n192), 
	.D(\reg_array[7][7] ), 
	.C(\reg_array[5][7] ), 
	.B(\reg_array[6][7] ), 
	.A(\reg_array[4][7] ));
   MUX4EHD U161 (.S1(N21), 
	.S0(N22), 
	.O(n193), 
	.D(\reg_array[3][7] ), 
	.C(\reg_array[1][7] ), 
	.B(\reg_array[2][7] ), 
	.A(\reg_array[0][7] ));
   MUX4EHD U162 (.S1(N21), 
	.S0(N22), 
	.O(n194), 
	.D(\reg_array[7][8] ), 
	.C(\reg_array[5][8] ), 
	.B(\reg_array[6][8] ), 
	.A(\reg_array[4][8] ));
   MUX4EHD U163 (.S1(N21), 
	.S0(N22), 
	.O(n195), 
	.D(\reg_array[3][8] ), 
	.C(\reg_array[1][8] ), 
	.B(\reg_array[2][8] ), 
	.A(\reg_array[0][8] ));
   MUX4EHD U164 (.S1(N21), 
	.S0(N22), 
	.O(n196), 
	.D(\reg_array[7][9] ), 
	.C(\reg_array[5][9] ), 
	.B(\reg_array[6][9] ), 
	.A(\reg_array[4][9] ));
   MUX4EHD U165 (.S1(N21), 
	.S0(N22), 
	.O(n197), 
	.D(\reg_array[3][9] ), 
	.C(\reg_array[1][9] ), 
	.B(\reg_array[2][9] ), 
	.A(\reg_array[0][9] ));
   MUX4EHD U166 (.S1(N21), 
	.S0(N22), 
	.O(n198), 
	.D(\reg_array[7][10] ), 
	.C(\reg_array[5][10] ), 
	.B(\reg_array[6][10] ), 
	.A(\reg_array[4][10] ));
   MUX4EHD U167 (.S1(N21), 
	.S0(N22), 
	.O(n199), 
	.D(\reg_array[3][10] ), 
	.C(\reg_array[1][10] ), 
	.B(\reg_array[2][10] ), 
	.A(\reg_array[0][10] ));
   MUX4EHD U168 (.S1(N21), 
	.S0(N22), 
	.O(n200), 
	.D(\reg_array[7][11] ), 
	.C(\reg_array[5][11] ), 
	.B(\reg_array[6][11] ), 
	.A(\reg_array[4][11] ));
   MUX4EHD U169 (.S1(N21), 
	.S0(N22), 
	.O(n201), 
	.D(\reg_array[3][11] ), 
	.C(\reg_array[1][11] ), 
	.B(\reg_array[2][11] ), 
	.A(\reg_array[0][11] ));
   MUX4EHD U170 (.S1(N21), 
	.S0(N22), 
	.O(n202), 
	.D(\reg_array[7][12] ), 
	.C(\reg_array[5][12] ), 
	.B(\reg_array[6][12] ), 
	.A(\reg_array[4][12] ));
   MUX4EHD U171 (.S1(N21), 
	.S0(N22), 
	.O(n203), 
	.D(\reg_array[3][12] ), 
	.C(\reg_array[1][12] ), 
	.B(\reg_array[2][12] ), 
	.A(\reg_array[0][12] ));
   MUX4EHD U172 (.S1(N21), 
	.S0(N22), 
	.O(n204), 
	.D(\reg_array[7][13] ), 
	.C(\reg_array[5][13] ), 
	.B(\reg_array[6][13] ), 
	.A(\reg_array[4][13] ));
   MUX4EHD U173 (.S1(N21), 
	.S0(N22), 
	.O(n205), 
	.D(\reg_array[3][13] ), 
	.C(\reg_array[1][13] ), 
	.B(\reg_array[2][13] ), 
	.A(\reg_array[0][13] ));
   MUX4EHD U174 (.S1(N21), 
	.S0(N22), 
	.O(n206), 
	.D(\reg_array[7][14] ), 
	.C(\reg_array[5][14] ), 
	.B(\reg_array[6][14] ), 
	.A(\reg_array[4][14] ));
   MUX4EHD U175 (.S1(N21), 
	.S0(N22), 
	.O(n207), 
	.D(\reg_array[3][14] ), 
	.C(\reg_array[1][14] ), 
	.B(\reg_array[2][14] ), 
	.A(\reg_array[0][14] ));
   MUX4EHD U176 (.S1(N21), 
	.S0(N22), 
	.O(n208), 
	.D(\reg_array[7][15] ), 
	.C(\reg_array[5][15] ), 
	.B(\reg_array[6][15] ), 
	.A(\reg_array[4][15] ));
   MUX4EHD U177 (.S1(N21), 
	.S0(N22), 
	.O(n209), 
	.D(\reg_array[3][15] ), 
	.C(\reg_array[1][15] ), 
	.B(\reg_array[2][15] ), 
	.A(\reg_array[0][15] ));
endmodule

module control (
	opcode, 
	reset, 
	reg_dst, 
	mem_to_reg, 
	alu_op, 
	jump, 
	branch, 
	mem_read, 
	mem_write, 
	alu_src, 
	reg_write, 
	sign_or_zero, 
	n75);
   input [2:0] opcode;
   input reset;
   output [1:0] reg_dst;
   output [1:0] mem_to_reg;
   output [1:0] alu_op;
   output jump;
   output branch;
   output mem_read;
   output mem_write;
   output alu_src;
   output reg_write;
   output sign_or_zero;
   input n75;

   // Internal wires
   wire \mem_to_reg[1] ;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n1;
   wire n2;
   wire n3;

   assign reg_dst[1] = \mem_to_reg[1]  ;
   assign mem_to_reg[1] = \mem_to_reg[1]  ;
   assign mem_to_reg[0] = mem_read ;
   assign alu_op[1] = alu_src ;

   AO12EHD U4 (.O(reg_write), 
	.B2(n75), 
	.B1(n7), 
	.A1(\mem_to_reg[1] ));
   OA13EHD U11 (.O(alu_src), 
	.B3(n13), 
	.B2(n9), 
	.B1(n12), 
	.A1(n75));
   ND2DHD U3 (.O(n12), 
	.I2(n8), 
	.I1(n14));
   OR3EHD U5 (.O(alu_op[0]), 
	.I3(branch), 
	.I2(mem_write), 
	.I1(mem_read));
   AN2HHD U6 (.O(mem_write), 
	.I2(n75), 
	.I1(n13));
   AN2EHD U7 (.O(reg_dst[0]), 
	.I2(n6), 
	.I1(n3));
   ND2DHD U8 (.O(sign_or_zero), 
	.I2(n6), 
	.I1(opcode[0]));
   NR2CHD U10 (.O(mem_read), 
	.I2(reset), 
	.I1(n14));
   AN2EHD U12 (.O(branch), 
	.I2(opcode[2]), 
	.I1(n11));
   NR2CHD U13 (.O(n11), 
	.I2(reset), 
	.I1(n2));
   OAI112BHD U14 (.O(n7), 
	.C2(opcode[0]), 
	.C1(opcode[1]), 
	.B1(n8), 
	.A1(n1));
   INVDHD U15 (.O(n1), 
	.I(n9));
   AN3EHD U16 (.O(\mem_to_reg[1] ), 
	.I3(n10), 
	.I2(opcode[1]), 
	.I1(opcode[0]));
   NR2CHD U17 (.O(n10), 
	.I2(opcode[2]), 
	.I1(reset));
   NR3BHD U18 (.O(n6), 
	.I3(opcode[1]), 
	.I2(reset), 
	.I1(opcode[2]));
   AN2B1CHD U19 (.O(jump), 
	.I1(n11), 
	.B1(opcode[2]));
   INVDHD U20 (.O(n2), 
	.I(opcode[1]));
   ND3CHD U21 (.O(n14), 
	.I3(opcode[2]), 
	.I2(n2), 
	.I1(n3));
   ND3CHD U22 (.O(n8), 
	.I3(opcode[0]), 
	.I2(opcode[2]), 
	.I1(opcode[1]));
   NR3BHD U23 (.O(n9), 
	.I3(n3), 
	.I2(opcode[2]), 
	.I1(opcode[1]));
   INVDHD U24 (.O(n3), 
	.I(opcode[0]));
   AN3EHD U25 (.O(n13), 
	.I3(opcode[0]), 
	.I2(n2), 
	.I1(opcode[2]));
endmodule

module instr_mem (
	pc, 
	instruction);
   input [15:0] pc;
   output [15:0] instruction;

   // Internal wires
   wire \instruction[0] ;

   assign instruction[15] = \instruction[0]  ;
   assign instruction[14] = \instruction[0]  ;
   assign instruction[13] = \instruction[0]  ;
   assign instruction[12] = \instruction[0]  ;
   assign instruction[11] = \instruction[0]  ;
   assign instruction[10] = \instruction[0]  ;
   assign instruction[9] = \instruction[0]  ;
   assign instruction[8] = \instruction[0]  ;
   assign instruction[7] = \instruction[0]  ;
   assign instruction[6] = \instruction[0]  ;
   assign instruction[5] = \instruction[0]  ;
   assign instruction[4] = \instruction[0]  ;
   assign instruction[3] = \instruction[0]  ;
   assign instruction[2] = \instruction[0]  ;
   assign instruction[1] = \instruction[0]  ;
   assign instruction[0] = \instruction[0]  ;

   TIE0DHD U2 (.O(\instruction[0] ));
endmodule

module mips_16 (
	clk, 
	reset, 
	pc_out, 
	alu_result, 
	clk_m__L3_N1, 
	clk_m__L3_N10, 
	clk_m__L3_N100, 
	clk_m__L3_N101, 
	clk_m__L3_N102, 
	clk_m__L3_N103, 
	clk_m__L3_N104, 
	clk_m__L3_N105, 
	clk_m__L3_N106, 
	clk_m__L3_N107, 
	clk_m__L3_N108, 
	clk_m__L3_N109, 
	clk_m__L3_N11, 
	clk_m__L3_N110, 
	clk_m__L3_N111, 
	clk_m__L3_N112, 
	clk_m__L3_N113, 
	clk_m__L3_N114, 
	clk_m__L3_N115, 
	clk_m__L3_N116, 
	clk_m__L3_N117, 
	clk_m__L3_N118, 
	clk_m__L3_N119, 
	clk_m__L3_N12, 
	clk_m__L3_N120, 
	clk_m__L3_N121, 
	clk_m__L3_N122, 
	clk_m__L3_N123, 
	clk_m__L3_N124, 
	clk_m__L3_N125, 
	clk_m__L3_N126, 
	clk_m__L3_N127, 
	clk_m__L3_N128, 
	clk_m__L3_N129, 
	clk_m__L3_N13, 
	clk_m__L3_N130, 
	clk_m__L3_N131, 
	clk_m__L3_N132, 
	clk_m__L3_N133, 
	clk_m__L3_N134, 
	clk_m__L3_N135, 
	clk_m__L3_N136, 
	clk_m__L3_N137, 
	clk_m__L3_N138, 
	clk_m__L3_N139, 
	clk_m__L3_N14, 
	clk_m__L3_N140, 
	clk_m__L3_N141, 
	clk_m__L3_N142, 
	clk_m__L3_N143, 
	clk_m__L3_N144, 
	clk_m__L3_N145, 
	clk_m__L3_N146, 
	clk_m__L3_N147, 
	clk_m__L3_N148, 
	clk_m__L3_N149, 
	clk_m__L3_N15, 
	clk_m__L3_N150, 
	clk_m__L3_N151, 
	clk_m__L3_N152, 
	clk_m__L3_N153, 
	clk_m__L3_N154, 
	clk_m__L3_N155, 
	clk_m__L3_N156, 
	clk_m__L3_N157, 
	clk_m__L3_N158, 
	clk_m__L3_N159, 
	clk_m__L3_N16, 
	clk_m__L3_N160, 
	clk_m__L3_N161, 
	clk_m__L3_N162, 
	clk_m__L3_N163, 
	clk_m__L3_N164, 
	clk_m__L3_N165, 
	clk_m__L3_N166, 
	clk_m__L3_N167, 
	clk_m__L3_N168, 
	clk_m__L3_N169, 
	clk_m__L3_N17, 
	clk_m__L3_N170, 
	clk_m__L3_N171, 
	clk_m__L3_N172, 
	clk_m__L3_N173, 
	clk_m__L3_N174, 
	clk_m__L3_N175, 
	clk_m__L3_N176, 
	clk_m__L3_N177, 
	clk_m__L3_N18, 
	clk_m__L3_N19, 
	clk_m__L3_N2, 
	clk_m__L3_N20, 
	clk_m__L3_N21, 
	clk_m__L3_N22, 
	clk_m__L3_N23, 
	clk_m__L3_N24, 
	clk_m__L3_N25, 
	clk_m__L3_N26, 
	clk_m__L3_N27, 
	clk_m__L3_N28, 
	clk_m__L3_N29, 
	clk_m__L3_N3, 
	clk_m__L3_N30, 
	clk_m__L3_N31, 
	clk_m__L3_N32, 
	clk_m__L3_N33, 
	clk_m__L3_N34, 
	clk_m__L3_N35, 
	clk_m__L3_N36, 
	clk_m__L3_N37, 
	clk_m__L3_N38, 
	clk_m__L3_N39, 
	clk_m__L3_N4, 
	clk_m__L3_N40, 
	clk_m__L3_N41, 
	clk_m__L3_N42, 
	clk_m__L3_N43, 
	clk_m__L3_N44, 
	clk_m__L3_N45, 
	clk_m__L3_N46, 
	clk_m__L3_N47, 
	clk_m__L3_N48, 
	clk_m__L3_N49, 
	clk_m__L3_N5, 
	clk_m__L3_N50, 
	clk_m__L3_N51, 
	clk_m__L3_N52, 
	clk_m__L3_N53, 
	clk_m__L3_N54, 
	clk_m__L3_N55, 
	clk_m__L3_N56, 
	clk_m__L3_N57, 
	clk_m__L3_N58, 
	clk_m__L3_N59, 
	clk_m__L3_N6, 
	clk_m__L3_N60, 
	clk_m__L3_N61, 
	clk_m__L3_N62, 
	clk_m__L3_N63, 
	clk_m__L3_N64, 
	clk_m__L3_N65, 
	clk_m__L3_N66, 
	clk_m__L3_N67, 
	clk_m__L3_N68, 
	clk_m__L3_N69, 
	clk_m__L3_N7, 
	clk_m__L3_N70, 
	clk_m__L3_N71, 
	clk_m__L3_N72, 
	clk_m__L3_N73, 
	clk_m__L3_N74, 
	clk_m__L3_N75, 
	clk_m__L3_N76, 
	clk_m__L3_N77, 
	clk_m__L3_N78, 
	clk_m__L3_N79, 
	clk_m__L3_N8, 
	clk_m__L3_N80, 
	clk_m__L3_N81, 
	clk_m__L3_N82, 
	clk_m__L3_N83, 
	clk_m__L3_N84, 
	clk_m__L3_N85, 
	clk_m__L3_N86, 
	clk_m__L3_N87, 
	clk_m__L3_N88, 
	clk_m__L3_N89, 
	clk_m__L3_N9, 
	clk_m__L3_N90, 
	clk_m__L3_N91, 
	clk_m__L3_N92, 
	clk_m__L3_N93, 
	clk_m__L3_N94, 
	clk_m__L3_N95, 
	clk_m__L3_N96, 
	clk_m__L3_N97, 
	clk_m__L3_N98, 
	clk_m__L3_N99, 
	clk_m__N0);
   input clk;
   input reset;
   output [15:0] pc_out;
   output [15:0] alu_result;
   input clk_m__L3_N1;
   input clk_m__L3_N10;
   input clk_m__L3_N100;
   input clk_m__L3_N101;
   input clk_m__L3_N102;
   input clk_m__L3_N103;
   input clk_m__L3_N104;
   input clk_m__L3_N105;
   input clk_m__L3_N106;
   input clk_m__L3_N107;
   input clk_m__L3_N108;
   input clk_m__L3_N109;
   input clk_m__L3_N11;
   input clk_m__L3_N110;
   input clk_m__L3_N111;
   input clk_m__L3_N112;
   input clk_m__L3_N113;
   input clk_m__L3_N114;
   input clk_m__L3_N115;
   input clk_m__L3_N116;
   input clk_m__L3_N117;
   input clk_m__L3_N118;
   input clk_m__L3_N119;
   input clk_m__L3_N12;
   input clk_m__L3_N120;
   input clk_m__L3_N121;
   input clk_m__L3_N122;
   input clk_m__L3_N123;
   input clk_m__L3_N124;
   input clk_m__L3_N125;
   input clk_m__L3_N126;
   input clk_m__L3_N127;
   input clk_m__L3_N128;
   input clk_m__L3_N129;
   input clk_m__L3_N13;
   input clk_m__L3_N130;
   input clk_m__L3_N131;
   input clk_m__L3_N132;
   input clk_m__L3_N133;
   input clk_m__L3_N134;
   input clk_m__L3_N135;
   input clk_m__L3_N136;
   input clk_m__L3_N137;
   input clk_m__L3_N138;
   input clk_m__L3_N139;
   input clk_m__L3_N14;
   input clk_m__L3_N140;
   input clk_m__L3_N141;
   input clk_m__L3_N142;
   input clk_m__L3_N143;
   input clk_m__L3_N144;
   input clk_m__L3_N145;
   input clk_m__L3_N146;
   input clk_m__L3_N147;
   input clk_m__L3_N148;
   input clk_m__L3_N149;
   input clk_m__L3_N15;
   input clk_m__L3_N150;
   input clk_m__L3_N151;
   input clk_m__L3_N152;
   input clk_m__L3_N153;
   input clk_m__L3_N154;
   input clk_m__L3_N155;
   input clk_m__L3_N156;
   input clk_m__L3_N157;
   input clk_m__L3_N158;
   input clk_m__L3_N159;
   input clk_m__L3_N16;
   input clk_m__L3_N160;
   input clk_m__L3_N161;
   input clk_m__L3_N162;
   input clk_m__L3_N163;
   input clk_m__L3_N164;
   input clk_m__L3_N165;
   input clk_m__L3_N166;
   input clk_m__L3_N167;
   input clk_m__L3_N168;
   input clk_m__L3_N169;
   input clk_m__L3_N17;
   input clk_m__L3_N170;
   input clk_m__L3_N171;
   input clk_m__L3_N172;
   input clk_m__L3_N173;
   input clk_m__L3_N174;
   input clk_m__L3_N175;
   input clk_m__L3_N176;
   input clk_m__L3_N177;
   input clk_m__L3_N18;
   input clk_m__L3_N19;
   input clk_m__L3_N2;
   input clk_m__L3_N20;
   input clk_m__L3_N21;
   input clk_m__L3_N22;
   input clk_m__L3_N23;
   input clk_m__L3_N24;
   input clk_m__L3_N25;
   input clk_m__L3_N26;
   input clk_m__L3_N27;
   input clk_m__L3_N28;
   input clk_m__L3_N29;
   input clk_m__L3_N3;
   input clk_m__L3_N30;
   input clk_m__L3_N31;
   input clk_m__L3_N32;
   input clk_m__L3_N33;
   input clk_m__L3_N34;
   input clk_m__L3_N35;
   input clk_m__L3_N36;
   input clk_m__L3_N37;
   input clk_m__L3_N38;
   input clk_m__L3_N39;
   input clk_m__L3_N4;
   input clk_m__L3_N40;
   input clk_m__L3_N41;
   input clk_m__L3_N42;
   input clk_m__L3_N43;
   input clk_m__L3_N44;
   input clk_m__L3_N45;
   input clk_m__L3_N46;
   input clk_m__L3_N47;
   input clk_m__L3_N48;
   input clk_m__L3_N49;
   input clk_m__L3_N5;
   input clk_m__L3_N50;
   input clk_m__L3_N51;
   input clk_m__L3_N52;
   input clk_m__L3_N53;
   input clk_m__L3_N54;
   input clk_m__L3_N55;
   input clk_m__L3_N56;
   input clk_m__L3_N57;
   input clk_m__L3_N58;
   input clk_m__L3_N59;
   input clk_m__L3_N6;
   input clk_m__L3_N60;
   input clk_m__L3_N61;
   input clk_m__L3_N62;
   input clk_m__L3_N63;
   input clk_m__L3_N64;
   input clk_m__L3_N65;
   input clk_m__L3_N66;
   input clk_m__L3_N67;
   input clk_m__L3_N68;
   input clk_m__L3_N69;
   input clk_m__L3_N7;
   input clk_m__L3_N70;
   input clk_m__L3_N71;
   input clk_m__L3_N72;
   input clk_m__L3_N73;
   input clk_m__L3_N74;
   input clk_m__L3_N75;
   input clk_m__L3_N76;
   input clk_m__L3_N77;
   input clk_m__L3_N78;
   input clk_m__L3_N79;
   input clk_m__L3_N8;
   input clk_m__L3_N80;
   input clk_m__L3_N81;
   input clk_m__L3_N82;
   input clk_m__L3_N83;
   input clk_m__L3_N84;
   input clk_m__L3_N85;
   input clk_m__L3_N86;
   input clk_m__L3_N87;
   input clk_m__L3_N88;
   input clk_m__L3_N89;
   input clk_m__L3_N9;
   input clk_m__L3_N90;
   input clk_m__L3_N91;
   input clk_m__L3_N92;
   input clk_m__L3_N93;
   input clk_m__L3_N94;
   input clk_m__L3_N95;
   input clk_m__L3_N96;
   input clk_m__L3_N97;
   input clk_m__L3_N98;
   input clk_m__L3_N99;
   input clk_m__N0;

   // Internal wires
   wire FE_OFN97_n1;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire jump;
   wire branch;
   wire mem_read;
   wire mem_write;
   wire alu_src;
   wire reg_write;
   wire JRControl;
   wire zero_flag;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N67;
   wire N68;
   wire n31;
   wire n35;
   wire n36;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n69;
   wire \add_47/carry[15] ;
   wire \add_47/carry[14] ;
   wire \add_47/carry[13] ;
   wire \add_47/carry[12] ;
   wire \add_47/carry[11] ;
   wire \add_47/carry[10] ;
   wire \add_47/carry[9] ;
   wire \add_47/carry[8] ;
   wire \add_47/carry[7] ;
   wire \add_47/carry[6] ;
   wire \add_47/carry[5] ;
   wire \add_47/carry[4] ;
   wire \add_47/carry[3] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n32;
   wire n33;
   wire n34;
   wire n37;
   wire n68;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire [15:0] pc_next;
   wire [1:0] reg_dst;
   wire [1:0] mem_to_reg;
   wire [1:0] alu_op;
   wire [15:0] reg_write_data;
   wire [15:0] reg_read_data_1;
   wire [15:0] reg_read_data_2;
   wire [2:0] ALU_Control;
   wire [15:0] mem_read_data;

   assign pc_out[0] = N53 ;

   BUFKHD FE_OFC97_n1 (.O(n1), 
	.I(FE_OFN97_n1));
   AO222EHD U14 (.O(reg_write_data[9]), 
	.C2(n4), 
	.C1(N62), 
	.B2(n3), 
	.B1(alu_result[9]), 
	.A2(n31), 
	.A1(mem_read_data[9]));
   AO222EHD U15 (.O(reg_write_data[8]), 
	.C2(n4), 
	.C1(N61), 
	.B2(n3), 
	.B1(alu_result[8]), 
	.A2(n31), 
	.A1(mem_read_data[8]));
   AO222EHD U16 (.O(reg_write_data[7]), 
	.C2(n4), 
	.C1(N60), 
	.B2(n3), 
	.B1(alu_result[7]), 
	.A2(n31), 
	.A1(mem_read_data[7]));
   AO222EHD U17 (.O(reg_write_data[6]), 
	.C2(n4), 
	.C1(N59), 
	.B2(n3), 
	.B1(alu_result[6]), 
	.A2(n31), 
	.A1(mem_read_data[6]));
   AO222EHD U18 (.O(reg_write_data[5]), 
	.C2(n4), 
	.C1(N58), 
	.B2(n3), 
	.B1(alu_result[5]), 
	.A2(n31), 
	.A1(mem_read_data[5]));
   AO222EHD U19 (.O(reg_write_data[4]), 
	.C2(n4), 
	.C1(N57), 
	.B2(n3), 
	.B1(alu_result[4]), 
	.A2(n31), 
	.A1(mem_read_data[4]));
   AO222EHD U20 (.O(reg_write_data[3]), 
	.C2(n4), 
	.C1(N56), 
	.B2(n3), 
	.B1(alu_result[3]), 
	.A2(n31), 
	.A1(mem_read_data[3]));
   AO222EHD U21 (.O(reg_write_data[2]), 
	.C2(n4), 
	.C1(N55), 
	.B2(n3), 
	.B1(alu_result[2]), 
	.A2(n31), 
	.A1(mem_read_data[2]));
   AO222EHD U22 (.O(reg_write_data[1]), 
	.C2(n4), 
	.C1(N54), 
	.B2(n3), 
	.B1(alu_result[1]), 
	.A2(n31), 
	.A1(mem_read_data[1]));
   AO222EHD U23 (.O(reg_write_data[15]), 
	.C2(n4), 
	.C1(N68), 
	.B2(n3), 
	.B1(alu_result[15]), 
	.A2(n31), 
	.A1(mem_read_data[15]));
   AO222EHD U24 (.O(reg_write_data[14]), 
	.C2(n4), 
	.C1(N67), 
	.B2(n3), 
	.B1(alu_result[14]), 
	.A2(n31), 
	.A1(mem_read_data[14]));
   AO222EHD U25 (.O(reg_write_data[13]), 
	.C2(n4), 
	.C1(N66), 
	.B2(n3), 
	.B1(alu_result[13]), 
	.A2(n31), 
	.A1(mem_read_data[13]));
   AO222EHD U26 (.O(reg_write_data[12]), 
	.C2(n4), 
	.C1(N65), 
	.B2(n3), 
	.B1(alu_result[12]), 
	.A2(n31), 
	.A1(mem_read_data[12]));
   AO222EHD U27 (.O(reg_write_data[11]), 
	.C2(n4), 
	.C1(N64), 
	.B2(n3), 
	.B1(alu_result[11]), 
	.A2(n31), 
	.A1(mem_read_data[11]));
   AO222EHD U28 (.O(reg_write_data[10]), 
	.C2(n4), 
	.C1(N63), 
	.B2(n3), 
	.B1(alu_result[10]), 
	.A2(n31), 
	.A1(mem_read_data[10]));
   AO222EHD U29 (.O(reg_write_data[0]), 
	.C2(n4), 
	.C1(N53), 
	.B2(n3), 
	.B1(alu_result[0]), 
	.A2(n31), 
	.A1(mem_read_data[0]));
   OR2B1CHD U117 (.O(n57), 
	.I1(JRControl), 
	.B1(jump));
   instr_mem instrucion_memory (.pc({ pc_out[15],
		pc_out[14],
		pc_out[13],
		pc_out[12],
		pc_out[11],
		pc_out[10],
		pc_out[9],
		pc_out[8],
		pc_out[7],
		pc_out[6],
		pc_out[5],
		pc_out[4],
		pc_out[3],
		pc_out[2],
		pc_out[1],
		N53 }));
   control control_unit (.opcode({ n1,
		n1,
		n1 }), 
	.reset(reset), 
	.reg_dst({ reg_dst[1],
		reg_dst[0] }), 
	.mem_to_reg({ mem_to_reg[1],
		mem_to_reg[0] }), 
	.alu_op({ alu_op[1],
		alu_op[0] }), 
	.jump(jump), 
	.branch(branch), 
	.mem_read(mem_read), 
	.mem_write(mem_write), 
	.alu_src(alu_src), 
	.reg_write(reg_write), 
	.n75(n75));
   register_file reg_file (.clk(clk_m__L3_N122), 
	.rst(reset), 
	.reg_write_en(reg_write), 
	.reg_write_dest({ n2,
		n2,
		n2 }), 
	.reg_write_data({ reg_write_data[15],
		reg_write_data[14],
		reg_write_data[13],
		reg_write_data[12],
		reg_write_data[11],
		reg_write_data[10],
		reg_write_data[9],
		reg_write_data[8],
		reg_write_data[7],
		reg_write_data[6],
		reg_write_data[5],
		reg_write_data[4],
		reg_write_data[3],
		reg_write_data[2],
		reg_write_data[1],
		reg_write_data[0] }), 
	.reg_read_addr_1({ n1,
		n1,
		n1 }), 
	.reg_read_data_1({ reg_read_data_1[15],
		reg_read_data_1[14],
		reg_read_data_1[13],
		reg_read_data_1[12],
		reg_read_data_1[11],
		reg_read_data_1[10],
		reg_read_data_1[9],
		reg_read_data_1[8],
		reg_read_data_1[7],
		reg_read_data_1[6],
		reg_read_data_1[5],
		reg_read_data_1[4],
		reg_read_data_1[3],
		reg_read_data_1[2],
		reg_read_data_1[1],
		reg_read_data_1[0] }), 
	.reg_read_addr_2({ n1,
		n1,
		n1 }), 
	.reg_read_data_2({ reg_read_data_2[15],
		reg_read_data_2[14],
		reg_read_data_2[13],
		reg_read_data_2[12],
		reg_read_data_2[11],
		reg_read_data_2[10],
		reg_read_data_2[9],
		reg_read_data_2[8],
		reg_read_data_2[7],
		reg_read_data_2[6],
		reg_read_data_2[5],
		reg_read_data_2[4],
		reg_read_data_2[3],
		reg_read_data_2[2],
		reg_read_data_2[1],
		reg_read_data_2[0] }), 
	.clk_m__L3_N123(clk_m__L3_N123), 
	.clk_m__L3_N124(clk_m__L3_N124), 
	.clk_m__L3_N126(clk_m__L3_N126), 
	.clk_m__L3_N154(clk_m__L3_N154), 
	.clk_m__L3_N49(clk_m__L3_N49), 
	.clk_m__L3_N50(clk_m__L3_N50), 
	.clk_m__L3_N51(clk_m__L3_N51), 
	.clk_m__L3_N53(clk_m__L3_N53), 
	.clk_m__L3_N54(clk_m__L3_N54), 
	.clk_m__L3_N80(clk_m__L3_N80));
   JR_Control JRControl_unit (.alu_op({ alu_op[1],
		alu_op[0] }), 
	.funct({ n1,
		n1,
		n1,
		n1 }), 
	.JRControl(JRControl));
   ALUControl ALU_Control_unit (.ALU_Control({ ALU_Control[2],
		ALU_Control[1],
		ALU_Control[0] }), 
	.ALUOp({ alu_op[1],
		alu_op[0] }), 
	.Function({ n1,
		n1,
		n1,
		n1 }));
   alu alu_unit (.a({ reg_read_data_1[15],
		reg_read_data_1[14],
		reg_read_data_1[13],
		reg_read_data_1[12],
		reg_read_data_1[11],
		reg_read_data_1[10],
		reg_read_data_1[9],
		reg_read_data_1[8],
		reg_read_data_1[7],
		reg_read_data_1[6],
		reg_read_data_1[5],
		reg_read_data_1[4],
		reg_read_data_1[3],
		reg_read_data_1[2],
		reg_read_data_1[1],
		reg_read_data_1[0] }), 
	.b({ n16,
		n20,
		n18,
		n19,
		n17,
		n15,
		n14,
		n13,
		n12,
		n11,
		n7,
		n5,
		n6,
		n9,
		n8,
		n10 }), 
	.alu_control({ ALU_Control[2],
		ALU_Control[1],
		ALU_Control[0] }), 
	.result({ alu_result[15],
		alu_result[14],
		alu_result[13],
		alu_result[12],
		alu_result[11],
		alu_result[10],
		alu_result[9],
		alu_result[8],
		n76,
		n77,
		n78,
		n79,
		n80,
		n81,
		alu_result[1],
		alu_result[0] }), 
	.zero(zero_flag));
   data_memory datamem (.clk(clk), 
	.mem_access_addr({ alu_result[15],
		alu_result[14],
		alu_result[13],
		alu_result[12],
		alu_result[11],
		alu_result[10],
		alu_result[9],
		alu_result[8],
		alu_result[7],
		alu_result[6],
		alu_result[5],
		alu_result[4],
		alu_result[3],
		alu_result[2],
		alu_result[1],
		alu_result[0] }), 
	.mem_write_data({ reg_read_data_2[15],
		reg_read_data_2[14],
		reg_read_data_2[13],
		reg_read_data_2[12],
		reg_read_data_2[11],
		reg_read_data_2[10],
		reg_read_data_2[9],
		reg_read_data_2[8],
		reg_read_data_2[7],
		reg_read_data_2[6],
		reg_read_data_2[5],
		reg_read_data_2[4],
		reg_read_data_2[3],
		reg_read_data_2[2],
		reg_read_data_2[1],
		reg_read_data_2[0] }), 
	.mem_write_en(mem_write), 
	.mem_read(mem_read), 
	.mem_read_data({ mem_read_data[15],
		mem_read_data[14],
		mem_read_data[13],
		mem_read_data[12],
		mem_read_data[11],
		mem_read_data[10],
		mem_read_data[9],
		mem_read_data[8],
		mem_read_data[7],
		mem_read_data[6],
		mem_read_data[5],
		mem_read_data[4],
		mem_read_data[3],
		mem_read_data[2],
		mem_read_data[1],
		mem_read_data[0] }), 
	.clk_m__L3_N1(clk_m__L3_N1), 
	.clk_m__L3_N10(clk_m__L3_N10), 
	.clk_m__L3_N100(clk_m__L3_N100), 
	.clk_m__L3_N101(clk_m__L3_N101), 
	.clk_m__L3_N102(clk_m__L3_N102), 
	.clk_m__L3_N103(clk_m__L3_N103), 
	.clk_m__L3_N104(clk_m__L3_N104), 
	.clk_m__L3_N105(clk_m__L3_N105), 
	.clk_m__L3_N106(clk_m__L3_N106), 
	.clk_m__L3_N107(clk_m__L3_N107), 
	.clk_m__L3_N108(clk_m__L3_N108), 
	.clk_m__L3_N109(clk_m__L3_N109), 
	.clk_m__L3_N11(clk_m__L3_N11), 
	.clk_m__L3_N110(clk_m__L3_N110), 
	.clk_m__L3_N111(clk_m__L3_N111), 
	.clk_m__L3_N112(clk_m__L3_N112), 
	.clk_m__L3_N113(clk_m__L3_N113), 
	.clk_m__L3_N114(clk_m__L3_N114), 
	.clk_m__L3_N115(clk_m__L3_N115), 
	.clk_m__L3_N116(clk_m__L3_N116), 
	.clk_m__L3_N117(clk_m__L3_N117), 
	.clk_m__L3_N118(clk_m__L3_N118), 
	.clk_m__L3_N119(clk_m__L3_N119), 
	.clk_m__L3_N12(clk_m__L3_N12), 
	.clk_m__L3_N120(clk_m__L3_N120), 
	.clk_m__L3_N121(clk_m__L3_N121), 
	.clk_m__L3_N122(clk_m__L3_N122), 
	.clk_m__L3_N123(clk_m__L3_N123), 
	.clk_m__L3_N124(clk_m__L3_N124), 
	.clk_m__L3_N125(clk_m__L3_N125), 
	.clk_m__L3_N126(clk_m__L3_N126), 
	.clk_m__L3_N127(clk_m__L3_N127), 
	.clk_m__L3_N128(clk_m__L3_N128), 
	.clk_m__L3_N129(clk_m__L3_N129), 
	.clk_m__L3_N13(clk_m__L3_N13), 
	.clk_m__L3_N130(clk_m__L3_N130), 
	.clk_m__L3_N131(clk_m__L3_N131), 
	.clk_m__L3_N132(clk_m__L3_N132), 
	.clk_m__L3_N133(clk_m__L3_N133), 
	.clk_m__L3_N134(clk_m__L3_N134), 
	.clk_m__L3_N135(clk_m__L3_N135), 
	.clk_m__L3_N136(clk_m__L3_N136), 
	.clk_m__L3_N137(clk_m__L3_N137), 
	.clk_m__L3_N138(clk_m__L3_N138), 
	.clk_m__L3_N139(clk_m__L3_N139), 
	.clk_m__L3_N14(clk_m__L3_N14), 
	.clk_m__L3_N140(clk_m__L3_N140), 
	.clk_m__L3_N141(clk_m__L3_N141), 
	.clk_m__L3_N142(clk_m__L3_N142), 
	.clk_m__L3_N143(clk_m__L3_N143), 
	.clk_m__L3_N144(clk_m__L3_N144), 
	.clk_m__L3_N145(clk_m__L3_N145), 
	.clk_m__L3_N146(clk_m__L3_N146), 
	.clk_m__L3_N147(clk_m__L3_N147), 
	.clk_m__L3_N148(clk_m__L3_N148), 
	.clk_m__L3_N149(clk_m__L3_N149), 
	.clk_m__L3_N15(clk_m__L3_N15), 
	.clk_m__L3_N150(clk_m__L3_N150), 
	.clk_m__L3_N151(clk_m__L3_N151), 
	.clk_m__L3_N152(clk_m__L3_N152), 
	.clk_m__L3_N153(clk_m__L3_N153), 
	.clk_m__L3_N154(clk_m__L3_N154), 
	.clk_m__L3_N155(clk_m__L3_N155), 
	.clk_m__L3_N156(clk_m__L3_N156), 
	.clk_m__L3_N157(clk_m__L3_N157), 
	.clk_m__L3_N158(clk_m__L3_N158), 
	.clk_m__L3_N159(clk_m__L3_N159), 
	.clk_m__L3_N16(clk_m__L3_N16), 
	.clk_m__L3_N160(clk_m__L3_N160), 
	.clk_m__L3_N161(clk_m__L3_N161), 
	.clk_m__L3_N162(clk_m__L3_N162), 
	.clk_m__L3_N163(clk_m__L3_N163), 
	.clk_m__L3_N164(clk_m__L3_N164), 
	.clk_m__L3_N165(clk_m__L3_N165), 
	.clk_m__L3_N166(clk_m__L3_N166), 
	.clk_m__L3_N167(clk_m__L3_N167), 
	.clk_m__L3_N168(clk_m__L3_N168), 
	.clk_m__L3_N169(clk_m__L3_N169), 
	.clk_m__L3_N17(clk_m__L3_N17), 
	.clk_m__L3_N170(clk_m__L3_N170), 
	.clk_m__L3_N171(clk_m__L3_N171), 
	.clk_m__L3_N172(clk_m__L3_N172), 
	.clk_m__L3_N173(clk_m__L3_N173), 
	.clk_m__L3_N174(clk_m__L3_N174), 
	.clk_m__L3_N175(clk_m__L3_N175), 
	.clk_m__L3_N176(clk_m__L3_N176), 
	.clk_m__L3_N177(clk_m__L3_N177), 
	.clk_m__L3_N18(clk_m__L3_N18), 
	.clk_m__L3_N19(clk_m__L3_N19), 
	.clk_m__L3_N2(clk_m__L3_N2), 
	.clk_m__L3_N20(clk_m__L3_N20), 
	.clk_m__L3_N21(clk_m__L3_N21), 
	.clk_m__L3_N22(clk_m__L3_N22), 
	.clk_m__L3_N23(clk_m__L3_N23), 
	.clk_m__L3_N24(clk_m__L3_N24), 
	.clk_m__L3_N25(clk_m__L3_N25), 
	.clk_m__L3_N26(clk_m__L3_N26), 
	.clk_m__L3_N27(clk_m__L3_N27), 
	.clk_m__L3_N28(clk_m__L3_N28), 
	.clk_m__L3_N29(clk_m__L3_N29), 
	.clk_m__L3_N3(clk_m__L3_N3), 
	.clk_m__L3_N30(clk_m__L3_N30), 
	.clk_m__L3_N31(clk_m__L3_N31), 
	.clk_m__L3_N32(clk_m__L3_N32), 
	.clk_m__L3_N33(clk_m__L3_N33), 
	.clk_m__L3_N34(clk_m__L3_N34), 
	.clk_m__L3_N35(clk_m__L3_N35), 
	.clk_m__L3_N36(clk_m__L3_N36), 
	.clk_m__L3_N37(clk_m__L3_N37), 
	.clk_m__L3_N38(clk_m__L3_N38), 
	.clk_m__L3_N39(clk_m__L3_N39), 
	.clk_m__L3_N4(clk_m__L3_N4), 
	.clk_m__L3_N40(clk_m__L3_N40), 
	.clk_m__L3_N41(clk_m__L3_N41), 
	.clk_m__L3_N42(clk_m__L3_N42), 
	.clk_m__L3_N43(clk_m__L3_N43), 
	.clk_m__L3_N44(clk_m__L3_N44), 
	.clk_m__L3_N45(clk_m__L3_N45), 
	.clk_m__L3_N46(clk_m__L3_N46), 
	.clk_m__L3_N47(clk_m__L3_N47), 
	.clk_m__L3_N48(clk_m__L3_N48), 
	.clk_m__L3_N49(clk_m__L3_N49), 
	.clk_m__L3_N5(clk_m__L3_N5), 
	.clk_m__L3_N50(clk_m__L3_N50), 
	.clk_m__L3_N52(clk_m__L3_N52), 
	.clk_m__L3_N53(clk_m__L3_N53), 
	.clk_m__L3_N54(clk_m__L3_N54), 
	.clk_m__L3_N55(clk_m__L3_N55), 
	.clk_m__L3_N56(clk_m__L3_N56), 
	.clk_m__L3_N57(clk_m__L3_N57), 
	.clk_m__L3_N58(clk_m__L3_N58), 
	.clk_m__L3_N59(clk_m__L3_N59), 
	.clk_m__L3_N6(clk_m__L3_N6), 
	.clk_m__L3_N60(clk_m__L3_N60), 
	.clk_m__L3_N61(clk_m__L3_N61), 
	.clk_m__L3_N62(clk_m__L3_N62), 
	.clk_m__L3_N63(clk_m__L3_N63), 
	.clk_m__L3_N64(clk_m__L3_N64), 
	.clk_m__L3_N65(clk_m__L3_N65), 
	.clk_m__L3_N66(clk_m__L3_N66), 
	.clk_m__L3_N67(clk_m__L3_N67), 
	.clk_m__L3_N68(clk_m__L3_N68), 
	.clk_m__L3_N69(clk_m__L3_N69), 
	.clk_m__L3_N7(clk_m__L3_N7), 
	.clk_m__L3_N70(clk_m__L3_N70), 
	.clk_m__L3_N71(clk_m__L3_N71), 
	.clk_m__L3_N72(clk_m__L3_N72), 
	.clk_m__L3_N73(clk_m__L3_N73), 
	.clk_m__L3_N74(clk_m__L3_N74), 
	.clk_m__L3_N75(clk_m__L3_N75), 
	.clk_m__L3_N76(clk_m__L3_N76), 
	.clk_m__L3_N77(clk_m__L3_N77), 
	.clk_m__L3_N78(clk_m__L3_N78), 
	.clk_m__L3_N79(clk_m__L3_N79), 
	.clk_m__L3_N8(clk_m__L3_N8), 
	.clk_m__L3_N80(clk_m__L3_N80), 
	.clk_m__L3_N81(clk_m__L3_N81), 
	.clk_m__L3_N82(clk_m__L3_N82), 
	.clk_m__L3_N83(clk_m__L3_N83), 
	.clk_m__L3_N84(clk_m__L3_N84), 
	.clk_m__L3_N85(clk_m__L3_N85), 
	.clk_m__L3_N86(clk_m__L3_N86), 
	.clk_m__L3_N87(clk_m__L3_N87), 
	.clk_m__L3_N88(clk_m__L3_N88), 
	.clk_m__L3_N89(clk_m__L3_N89), 
	.clk_m__L3_N9(clk_m__L3_N9), 
	.clk_m__L3_N90(clk_m__L3_N90), 
	.clk_m__L3_N91(clk_m__L3_N91), 
	.clk_m__L3_N92(clk_m__L3_N92), 
	.clk_m__L3_N93(clk_m__L3_N93), 
	.clk_m__L3_N94(clk_m__L3_N94), 
	.clk_m__L3_N95(clk_m__L3_N95), 
	.clk_m__L3_N96(clk_m__L3_N96), 
	.clk_m__L3_N97(clk_m__L3_N97), 
	.clk_m__L3_N98(clk_m__L3_N98), 
	.clk_m__L3_N99(clk_m__L3_N99), 
	.clk_m__N0(clk_m__N0));
   QDFFRBEHD \pc_current_reg[15]  (.RB(n75), 
	.Q(pc_out[15]), 
	.D(pc_next[15]), 
	.CK(clk_m__L3_N124));
   QDFFRBEHD \pc_current_reg[9]  (.RB(n75), 
	.Q(pc_out[9]), 
	.D(pc_next[9]), 
	.CK(clk_m__L3_N126));
   QDFFRBEHD \pc_current_reg[8]  (.RB(n75), 
	.Q(pc_out[8]), 
	.D(pc_next[8]), 
	.CK(clk_m__L3_N126));
   QDFFRBEHD \pc_current_reg[7]  (.RB(n75), 
	.Q(pc_out[7]), 
	.D(pc_next[7]), 
	.CK(clk_m__L3_N50));
   QDFFRBEHD \pc_current_reg[6]  (.RB(n75), 
	.Q(pc_out[6]), 
	.D(pc_next[6]), 
	.CK(clk_m__L3_N50));
   QDFFRBEHD \pc_current_reg[5]  (.RB(n75), 
	.Q(pc_out[5]), 
	.D(pc_next[5]), 
	.CK(clk_m__L3_N50));
   QDFFRBEHD \pc_current_reg[4]  (.RB(n75), 
	.Q(pc_out[4]), 
	.D(pc_next[4]), 
	.CK(clk_m__L3_N51));
   QDFFRBEHD \pc_current_reg[3]  (.RB(n75), 
	.Q(pc_out[3]), 
	.D(pc_next[3]), 
	.CK(clk_m__L3_N51));
   QDFFRBEHD \pc_current_reg[2]  (.RB(n75), 
	.Q(pc_out[2]), 
	.D(pc_next[2]), 
	.CK(clk_m__L3_N154));
   QDFFRBEHD \pc_current_reg[14]  (.RB(n75), 
	.Q(pc_out[14]), 
	.D(pc_next[14]), 
	.CK(clk_m__L3_N124));
   QDFFRBEHD \pc_current_reg[13]  (.RB(n75), 
	.Q(pc_out[13]), 
	.D(pc_next[13]), 
	.CK(clk_m__L3_N123));
   QDFFRBEHD \pc_current_reg[12]  (.RB(n75), 
	.Q(pc_out[12]), 
	.D(pc_next[12]), 
	.CK(clk_m__L3_N123));
   QDFFRBEHD \pc_current_reg[11]  (.RB(n75), 
	.Q(pc_out[11]), 
	.D(pc_next[11]), 
	.CK(clk_m__L3_N122));
   QDFFRBEHD \pc_current_reg[10]  (.RB(n75), 
	.Q(pc_out[10]), 
	.D(pc_next[10]), 
	.CK(clk_m__L3_N122));
   QDFFRBEHD \pc_current_reg[1]  (.RB(n75), 
	.Q(pc_out[1]), 
	.D(pc_next[1]), 
	.CK(clk_m__L3_N51));
   QDFFRBEHD \pc_current_reg[0]  (.RB(n75), 
	.Q(N53), 
	.D(pc_next[0]), 
	.CK(clk_m__L3_N154));
   TIE0KHD U3 (.O(FE_OFN97_n1));
   AN2EHD U4 (.O(n2), 
	.I2(n74), 
	.I1(reg_dst[1]));
   XNR2EHD U5 (.O(n3), 
	.I2(mem_to_reg[1]), 
	.I1(mem_to_reg[0]));
   AN2EHD U6 (.O(n4), 
	.I2(n72), 
	.I1(mem_to_reg[1]));
   INVDHD U7 (.O(n73), 
	.I(alu_src));
   BUFEHD U8 (.O(alu_result[6]), 
	.I(n77));
   BUFEHD U9 (.O(alu_result[7]), 
	.I(n76));
   BUFEHD U10 (.O(alu_result[4]), 
	.I(n79));
   BUFEHD U11 (.O(alu_result[2]), 
	.I(n81));
   BUFEHD U12 (.O(alu_result[5]), 
	.I(n78));
   BUFEHD U13 (.O(alu_result[3]), 
	.I(n80));
   INVDHD U30 (.O(n71), 
	.I(n69));
   AN2EHD U31 (.O(n5), 
	.I2(reg_read_data_2[4]), 
	.I1(n73));
   AN2EHD U32 (.O(n6), 
	.I2(reg_read_data_2[3]), 
	.I1(n73));
   AN2EHD U33 (.O(n7), 
	.I2(reg_read_data_2[5]), 
	.I1(n73));
   AN2EHD U34 (.O(n8), 
	.I2(reg_read_data_2[1]), 
	.I1(n73));
   AN2EHD U35 (.O(n9), 
	.I2(reg_read_data_2[2]), 
	.I1(n73));
   AN2EHD U36 (.O(n10), 
	.I2(reg_read_data_2[0]), 
	.I1(n73));
   AN2EHD U37 (.O(n11), 
	.I2(reg_read_data_2[6]), 
	.I1(n73));
   AN2EHD U38 (.O(n12), 
	.I2(n73), 
	.I1(reg_read_data_2[7]));
   AN2EHD U39 (.O(n13), 
	.I2(n73), 
	.I1(reg_read_data_2[8]));
   AN2EHD U40 (.O(n14), 
	.I2(n73), 
	.I1(reg_read_data_2[9]));
   AN2EHD U41 (.O(n15), 
	.I2(n73), 
	.I1(reg_read_data_2[10]));
   AN2EHD U42 (.O(n16), 
	.I2(n73), 
	.I1(reg_read_data_2[15]));
   AN2EHD U43 (.O(n17), 
	.I2(n73), 
	.I1(reg_read_data_2[11]));
   AN2EHD U44 (.O(n18), 
	.I2(n73), 
	.I1(reg_read_data_2[13]));
   AN2EHD U45 (.O(n19), 
	.I2(n73), 
	.I1(reg_read_data_2[12]));
   AN2EHD U46 (.O(n20), 
	.I2(n73), 
	.I1(reg_read_data_2[14]));
   NR3HHD U48 (.O(n38), 
	.I3(n69), 
	.I2(jump), 
	.I1(JRControl));
   ND3CHD U49 (.O(pc_next[15]), 
	.I3(n34), 
	.I2(n33), 
	.I1(n32));
   ND2DHD U50 (.O(n34), 
	.I2(JRControl), 
	.I1(reg_read_data_1[15]));
   ND2DHD U51 (.O(n33), 
	.I2(n56), 
	.I1(N68));
   ND2DHD U52 (.O(n32), 
	.I2(n38), 
	.I1(N68));
   OAI12CHD U53 (.O(n56), 
	.B2(n71), 
	.B1(JRControl), 
	.A1(n57));
   ND2DHD U54 (.O(n69), 
	.I2(branch), 
	.I1(zero_flag));
   NR3BHD U56 (.O(n39), 
	.I3(n71), 
	.I2(jump), 
	.I1(JRControl));
   ND2DHD U57 (.O(pc_next[10]), 
	.I2(n67), 
	.I1(n66));
   ND2DHD U58 (.O(n67), 
	.I2(n38), 
	.I1(N63));
   AOI22BHD U59 (.O(n66), 
	.B2(JRControl), 
	.B1(reg_read_data_1[10]), 
	.A2(N63), 
	.A1(n39));
   ND2DHD U60 (.O(pc_next[11]), 
	.I2(n65), 
	.I1(n64));
   ND2DHD U61 (.O(n65), 
	.I2(n38), 
	.I1(N64));
   AOI22BHD U62 (.O(n64), 
	.B2(JRControl), 
	.B1(reg_read_data_1[11]), 
	.A2(N64), 
	.A1(n39));
   ND2DHD U63 (.O(pc_next[12]), 
	.I2(n63), 
	.I1(n62));
   ND2DHD U64 (.O(n63), 
	.I2(n38), 
	.I1(N65));
   AOI22BHD U65 (.O(n62), 
	.B2(JRControl), 
	.B1(reg_read_data_1[12]), 
	.A2(N65), 
	.A1(n39));
   ND2DHD U66 (.O(pc_next[13]), 
	.I2(n61), 
	.I1(n60));
   ND2DHD U67 (.O(n61), 
	.I2(n38), 
	.I1(N66));
   AOI22BHD U68 (.O(n60), 
	.B2(JRControl), 
	.B1(reg_read_data_1[13]), 
	.A2(N66), 
	.A1(n39));
   ND2DHD U69 (.O(pc_next[14]), 
	.I2(n59), 
	.I1(n58));
   ND2DHD U70 (.O(n59), 
	.I2(n38), 
	.I1(N67));
   AOI22BHD U71 (.O(n58), 
	.B2(JRControl), 
	.B1(reg_read_data_1[14]), 
	.A2(N67), 
	.A1(n39));
   ND2DHD U72 (.O(pc_next[2]), 
	.I2(n53), 
	.I1(n52));
   ND2DHD U73 (.O(n53), 
	.I2(n38), 
	.I1(N55));
   AOI22BHD U74 (.O(n52), 
	.B2(JRControl), 
	.B1(reg_read_data_1[2]), 
	.A2(N55), 
	.A1(n39));
   ND2DHD U75 (.O(pc_next[3]), 
	.I2(n51), 
	.I1(n50));
   ND2DHD U76 (.O(n51), 
	.I2(n38), 
	.I1(N56));
   AOI22BHD U77 (.O(n50), 
	.B2(JRControl), 
	.B1(reg_read_data_1[3]), 
	.A2(N56), 
	.A1(n39));
   ND2DHD U78 (.O(pc_next[4]), 
	.I2(n49), 
	.I1(n48));
   ND2DHD U79 (.O(n49), 
	.I2(n38), 
	.I1(N57));
   AOI22BHD U80 (.O(n48), 
	.B2(JRControl), 
	.B1(reg_read_data_1[4]), 
	.A2(N57), 
	.A1(n39));
   ND2DHD U81 (.O(pc_next[5]), 
	.I2(n47), 
	.I1(n46));
   ND2DHD U82 (.O(n47), 
	.I2(n38), 
	.I1(N58));
   AOI22BHD U83 (.O(n46), 
	.B2(JRControl), 
	.B1(reg_read_data_1[5]), 
	.A2(N58), 
	.A1(n39));
   ND2DHD U84 (.O(pc_next[6]), 
	.I2(n45), 
	.I1(n44));
   ND2DHD U85 (.O(n45), 
	.I2(n38), 
	.I1(N59));
   AOI22BHD U86 (.O(n44), 
	.B2(JRControl), 
	.B1(reg_read_data_1[6]), 
	.A2(N59), 
	.A1(n39));
   ND2DHD U87 (.O(pc_next[7]), 
	.I2(n43), 
	.I1(n42));
   ND2DHD U88 (.O(n43), 
	.I2(n38), 
	.I1(N60));
   AOI22BHD U89 (.O(n42), 
	.B2(JRControl), 
	.B1(reg_read_data_1[7]), 
	.A2(N60), 
	.A1(n39));
   ND2DHD U90 (.O(pc_next[8]), 
	.I2(n41), 
	.I1(n40));
   ND2DHD U91 (.O(n41), 
	.I2(n38), 
	.I1(N61));
   AOI22BHD U92 (.O(n40), 
	.B2(JRControl), 
	.B1(reg_read_data_1[8]), 
	.A2(N61), 
	.A1(n39));
   ND2DHD U93 (.O(pc_next[9]), 
	.I2(n36), 
	.I1(n35));
   ND2DHD U94 (.O(n36), 
	.I2(n38), 
	.I1(N62));
   AOI22BHD U95 (.O(n35), 
	.B2(JRControl), 
	.B1(reg_read_data_1[9]), 
	.A2(N62), 
	.A1(n39));
   ND2DHD U96 (.O(pc_next[1]), 
	.I2(n55), 
	.I1(n54));
   ND2DHD U97 (.O(n55), 
	.I2(n38), 
	.I1(N54));
   AOI22BHD U98 (.O(n54), 
	.B2(JRControl), 
	.B1(reg_read_data_1[1]), 
	.A2(N54), 
	.A1(n39));
   NR2CHD U100 (.O(n31), 
	.I2(mem_to_reg[1]), 
	.I1(n72));
   INVDHD U101 (.O(n72), 
	.I(mem_to_reg[0]));
   INVDHD U102 (.O(n74), 
	.I(reg_dst[0]));
   ND3CHD U103 (.O(pc_next[0]), 
	.I3(n70), 
	.I2(n68), 
	.I1(n37));
   ND2DHD U104 (.O(n70), 
	.I2(JRControl), 
	.I1(reg_read_data_1[0]));
   ND2DHD U105 (.O(n37), 
	.I2(N53), 
	.I1(n39));
   ND2DHD U106 (.O(n68), 
	.I2(n38), 
	.I1(N53));
   INVDHD U108 (.O(N54), 
	.I(pc_out[1]));
   INVDHD U109 (.O(n75), 
	.I(reset));
   XOR2CHD U110 (.O(N68), 
	.I2(\add_47/carry[15] ), 
	.I1(pc_out[15]));
   AN2CHD U111 (.O(\add_47/carry[15] ), 
	.I2(\add_47/carry[14] ), 
	.I1(pc_out[14]));
   XOR2CHD U112 (.O(N67), 
	.I2(\add_47/carry[14] ), 
	.I1(pc_out[14]));
   AN2CHD U113 (.O(\add_47/carry[14] ), 
	.I2(\add_47/carry[13] ), 
	.I1(pc_out[13]));
   XOR2CHD U114 (.O(N66), 
	.I2(\add_47/carry[13] ), 
	.I1(pc_out[13]));
   AN2CHD U115 (.O(\add_47/carry[13] ), 
	.I2(\add_47/carry[12] ), 
	.I1(pc_out[12]));
   XOR2CHD U116 (.O(N65), 
	.I2(\add_47/carry[12] ), 
	.I1(pc_out[12]));
   AN2CHD U118 (.O(\add_47/carry[12] ), 
	.I2(\add_47/carry[11] ), 
	.I1(pc_out[11]));
   XOR2CHD U119 (.O(N64), 
	.I2(\add_47/carry[11] ), 
	.I1(pc_out[11]));
   AN2CHD U120 (.O(\add_47/carry[11] ), 
	.I2(\add_47/carry[10] ), 
	.I1(pc_out[10]));
   XOR2CHD U121 (.O(N63), 
	.I2(\add_47/carry[10] ), 
	.I1(pc_out[10]));
   AN2CHD U122 (.O(\add_47/carry[10] ), 
	.I2(\add_47/carry[9] ), 
	.I1(pc_out[9]));
   XOR2CHD U123 (.O(N62), 
	.I2(\add_47/carry[9] ), 
	.I1(pc_out[9]));
   AN2CHD U124 (.O(\add_47/carry[9] ), 
	.I2(\add_47/carry[8] ), 
	.I1(pc_out[8]));
   XOR2CHD U125 (.O(N61), 
	.I2(\add_47/carry[8] ), 
	.I1(pc_out[8]));
   AN2CHD U126 (.O(\add_47/carry[8] ), 
	.I2(\add_47/carry[7] ), 
	.I1(pc_out[7]));
   XOR2CHD U127 (.O(N60), 
	.I2(\add_47/carry[7] ), 
	.I1(pc_out[7]));
   AN2CHD U128 (.O(\add_47/carry[7] ), 
	.I2(\add_47/carry[6] ), 
	.I1(pc_out[6]));
   XOR2CHD U129 (.O(N59), 
	.I2(\add_47/carry[6] ), 
	.I1(pc_out[6]));
   AN2CHD U130 (.O(\add_47/carry[6] ), 
	.I2(\add_47/carry[5] ), 
	.I1(pc_out[5]));
   XOR2CHD U131 (.O(N58), 
	.I2(\add_47/carry[5] ), 
	.I1(pc_out[5]));
   AN2CHD U132 (.O(\add_47/carry[5] ), 
	.I2(\add_47/carry[4] ), 
	.I1(pc_out[4]));
   XOR2CHD U133 (.O(N57), 
	.I2(\add_47/carry[4] ), 
	.I1(pc_out[4]));
   AN2CHD U134 (.O(\add_47/carry[4] ), 
	.I2(\add_47/carry[3] ), 
	.I1(pc_out[3]));
   XOR2CHD U135 (.O(N56), 
	.I2(\add_47/carry[3] ), 
	.I1(pc_out[3]));
   AN2CHD U136 (.O(\add_47/carry[3] ), 
	.I2(pc_out[1]), 
	.I1(pc_out[2]));
   XOR2CHD U137 (.O(N55), 
	.I2(pc_out[1]), 
	.I1(pc_out[2]));
endmodule

module mips (
	vdd, 
	vddio, 
	gnd, 
	vss, 
	clk, 
	reset, 
	pc_out, 
	alu_result);
   inout vdd;
   inout vddio;
   inout gnd;
   inout vss;
   input clk;
   input reset;
   output [15:0] pc_out;
   output [15:0] alu_result;

   // Internal wires
   wire clk_m__N0;
   wire clk_m__L3_N177;
   wire clk_m__L3_N176;
   wire clk_m__L3_N175;
   wire clk_m__L3_N174;
   wire clk_m__L3_N173;
   wire clk_m__L3_N172;
   wire clk_m__L3_N171;
   wire clk_m__L3_N170;
   wire clk_m__L3_N169;
   wire clk_m__L3_N168;
   wire clk_m__L3_N167;
   wire clk_m__L3_N166;
   wire clk_m__L3_N165;
   wire clk_m__L3_N164;
   wire clk_m__L3_N163;
   wire clk_m__L3_N162;
   wire clk_m__L3_N161;
   wire clk_m__L3_N160;
   wire clk_m__L3_N159;
   wire clk_m__L3_N158;
   wire clk_m__L3_N157;
   wire clk_m__L3_N156;
   wire clk_m__L3_N155;
   wire clk_m__L3_N154;
   wire clk_m__L3_N153;
   wire clk_m__L3_N152;
   wire clk_m__L3_N151;
   wire clk_m__L3_N150;
   wire clk_m__L3_N149;
   wire clk_m__L3_N148;
   wire clk_m__L3_N147;
   wire clk_m__L3_N146;
   wire clk_m__L3_N145;
   wire clk_m__L3_N144;
   wire clk_m__L3_N143;
   wire clk_m__L3_N142;
   wire clk_m__L3_N141;
   wire clk_m__L3_N140;
   wire clk_m__L3_N139;
   wire clk_m__L3_N138;
   wire clk_m__L3_N137;
   wire clk_m__L3_N136;
   wire clk_m__L3_N135;
   wire clk_m__L3_N134;
   wire clk_m__L3_N133;
   wire clk_m__L3_N132;
   wire clk_m__L3_N131;
   wire clk_m__L3_N130;
   wire clk_m__L3_N129;
   wire clk_m__L3_N128;
   wire clk_m__L3_N127;
   wire clk_m__L3_N126;
   wire clk_m__L3_N125;
   wire clk_m__L3_N124;
   wire clk_m__L3_N123;
   wire clk_m__L3_N122;
   wire clk_m__L3_N121;
   wire clk_m__L3_N120;
   wire clk_m__L3_N119;
   wire clk_m__L3_N118;
   wire clk_m__L3_N117;
   wire clk_m__L3_N116;
   wire clk_m__L3_N115;
   wire clk_m__L3_N114;
   wire clk_m__L3_N113;
   wire clk_m__L3_N112;
   wire clk_m__L3_N111;
   wire clk_m__L3_N110;
   wire clk_m__L3_N109;
   wire clk_m__L3_N108;
   wire clk_m__L3_N107;
   wire clk_m__L3_N106;
   wire clk_m__L3_N105;
   wire clk_m__L3_N104;
   wire clk_m__L3_N103;
   wire clk_m__L3_N102;
   wire clk_m__L3_N101;
   wire clk_m__L3_N100;
   wire clk_m__L3_N99;
   wire clk_m__L3_N98;
   wire clk_m__L3_N97;
   wire clk_m__L3_N96;
   wire clk_m__L3_N95;
   wire clk_m__L3_N94;
   wire clk_m__L3_N93;
   wire clk_m__L3_N92;
   wire clk_m__L3_N91;
   wire clk_m__L3_N90;
   wire clk_m__L3_N89;
   wire clk_m__L3_N88;
   wire clk_m__L3_N87;
   wire clk_m__L3_N86;
   wire clk_m__L3_N85;
   wire clk_m__L3_N84;
   wire clk_m__L3_N83;
   wire clk_m__L3_N82;
   wire clk_m__L3_N81;
   wire clk_m__L3_N80;
   wire clk_m__L3_N79;
   wire clk_m__L3_N78;
   wire clk_m__L3_N77;
   wire clk_m__L3_N76;
   wire clk_m__L3_N75;
   wire clk_m__L3_N74;
   wire clk_m__L3_N73;
   wire clk_m__L3_N72;
   wire clk_m__L3_N71;
   wire clk_m__L3_N70;
   wire clk_m__L3_N69;
   wire clk_m__L3_N68;
   wire clk_m__L3_N67;
   wire clk_m__L3_N66;
   wire clk_m__L3_N65;
   wire clk_m__L3_N64;
   wire clk_m__L3_N63;
   wire clk_m__L3_N62;
   wire clk_m__L3_N61;
   wire clk_m__L3_N60;
   wire clk_m__L3_N59;
   wire clk_m__L3_N58;
   wire clk_m__L3_N57;
   wire clk_m__L3_N56;
   wire clk_m__L3_N55;
   wire clk_m__L3_N54;
   wire clk_m__L3_N53;
   wire clk_m__L3_N52;
   wire clk_m__L3_N51;
   wire clk_m__L3_N50;
   wire clk_m__L3_N49;
   wire clk_m__L3_N48;
   wire clk_m__L3_N47;
   wire clk_m__L3_N46;
   wire clk_m__L3_N45;
   wire clk_m__L3_N44;
   wire clk_m__L3_N43;
   wire clk_m__L3_N42;
   wire clk_m__L3_N41;
   wire clk_m__L3_N40;
   wire clk_m__L3_N39;
   wire clk_m__L3_N38;
   wire clk_m__L3_N37;
   wire clk_m__L3_N36;
   wire clk_m__L3_N35;
   wire clk_m__L3_N34;
   wire clk_m__L3_N33;
   wire clk_m__L3_N32;
   wire clk_m__L3_N31;
   wire clk_m__L3_N30;
   wire clk_m__L3_N29;
   wire clk_m__L3_N28;
   wire clk_m__L3_N27;
   wire clk_m__L3_N26;
   wire clk_m__L3_N25;
   wire clk_m__L3_N24;
   wire clk_m__L3_N23;
   wire clk_m__L3_N22;
   wire clk_m__L3_N21;
   wire clk_m__L3_N20;
   wire clk_m__L3_N19;
   wire clk_m__L3_N18;
   wire clk_m__L3_N17;
   wire clk_m__L3_N16;
   wire clk_m__L3_N15;
   wire clk_m__L3_N14;
   wire clk_m__L3_N13;
   wire clk_m__L3_N12;
   wire clk_m__L3_N11;
   wire clk_m__L3_N10;
   wire clk_m__L3_N9;
   wire clk_m__L3_N8;
   wire clk_m__L3_N7;
   wire clk_m__L3_N6;
   wire clk_m__L3_N5;
   wire clk_m__L3_N4;
   wire clk_m__L3_N3;
   wire clk_m__L3_N2;
   wire clk_m__L3_N1;
   wire clk_m__L3_N0;
   wire clk_m__L2_N17;
   wire clk_m__L2_N16;
   wire clk_m__L2_N15;
   wire clk_m__L2_N14;
   wire clk_m__L2_N13;
   wire clk_m__L2_N12;
   wire clk_m__L2_N11;
   wire clk_m__L2_N10;
   wire clk_m__L2_N9;
   wire clk_m__L2_N8;
   wire clk_m__L2_N7;
   wire clk_m__L2_N6;
   wire clk_m__L2_N5;
   wire clk_m__L2_N4;
   wire clk_m__L2_N3;
   wire clk_m__L2_N2;
   wire clk_m__L2_N1;
   wire clk_m__L2_N0;
   wire clk_m__L1_N5;
   wire clk_m__L1_N4;
   wire clk_m__L1_N3;
   wire clk_m__L1_N2;
   wire clk_m__L1_N1;
   wire clk_m__L1_N0;
   wire FE_OFN96_n1;
   wire clk_m;
   wire reset_m;
   wire n1;
   wire n2;
   wire [15:0] pc_out_m;
   wire [15:0] alu_result_m;

   BUFCKGHD clk_m__I0 (.O(clk_m__N0), 
	.I(clk_m__L2_N10));
   BUFCKGHD clk_m__L3_I177 (.O(clk_m__L3_N177), 
	.I(clk_m__L2_N17));
   BUFCKHHD clk_m__L3_I176 (.O(clk_m__L3_N176), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I175 (.O(clk_m__L3_N175), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I174 (.O(clk_m__L3_N174), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I173 (.O(clk_m__L3_N173), 
	.I(clk_m__L2_N17));
   BUFCKHHD clk_m__L3_I172 (.O(clk_m__L3_N172), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I171 (.O(clk_m__L3_N171), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I170 (.O(clk_m__L3_N170), 
	.I(clk_m__L2_N17));
   BUFCKHHD clk_m__L3_I169 (.O(clk_m__L3_N169), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I168 (.O(clk_m__L3_N168), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I167 (.O(clk_m__L3_N167), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I166 (.O(clk_m__L3_N166), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I165 (.O(clk_m__L3_N165), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I164 (.O(clk_m__L3_N164), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I163 (.O(clk_m__L3_N163), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I162 (.O(clk_m__L3_N162), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I161 (.O(clk_m__L3_N161), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I160 (.O(clk_m__L3_N160), 
	.I(clk_m__L2_N16));
   BUFCKHHD clk_m__L3_I159 (.O(clk_m__L3_N159), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I158 (.O(clk_m__L3_N158), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I157 (.O(clk_m__L3_N157), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I156 (.O(clk_m__L3_N156), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I155 (.O(clk_m__L3_N155), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I154 (.O(clk_m__L3_N154), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I153 (.O(clk_m__L3_N153), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I152 (.O(clk_m__L3_N152), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I151 (.O(clk_m__L3_N151), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I150 (.O(clk_m__L3_N150), 
	.I(clk_m__L2_N15));
   BUFCKHHD clk_m__L3_I149 (.O(clk_m__L3_N149), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I148 (.O(clk_m__L3_N148), 
	.I(clk_m__L2_N15));
   BUFCKHHD clk_m__L3_I147 (.O(clk_m__L3_N147), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I146 (.O(clk_m__L3_N146), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I145 (.O(clk_m__L3_N145), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I144 (.O(clk_m__L3_N144), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I143 (.O(clk_m__L3_N143), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I142 (.O(clk_m__L3_N142), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I141 (.O(clk_m__L3_N141), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I140 (.O(clk_m__L3_N140), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I139 (.O(clk_m__L3_N139), 
	.I(clk_m__L2_N14));
   BUFCKHHD clk_m__L3_I138 (.O(clk_m__L3_N138), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I137 (.O(clk_m__L3_N137), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I136 (.O(clk_m__L3_N136), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I135 (.O(clk_m__L3_N135), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I134 (.O(clk_m__L3_N134), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I133 (.O(clk_m__L3_N133), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I132 (.O(clk_m__L3_N132), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I131 (.O(clk_m__L3_N131), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I130 (.O(clk_m__L3_N130), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I129 (.O(clk_m__L3_N129), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I128 (.O(clk_m__L3_N128), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I127 (.O(clk_m__L3_N127), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I126 (.O(clk_m__L3_N126), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I125 (.O(clk_m__L3_N125), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I124 (.O(clk_m__L3_N124), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I123 (.O(clk_m__L3_N123), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I122 (.O(clk_m__L3_N122), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I121 (.O(clk_m__L3_N121), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I120 (.O(clk_m__L3_N120), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I119 (.O(clk_m__L3_N119), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I118 (.O(clk_m__L3_N118), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I117 (.O(clk_m__L3_N117), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I116 (.O(clk_m__L3_N116), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I115 (.O(clk_m__L3_N115), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I114 (.O(clk_m__L3_N114), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I113 (.O(clk_m__L3_N113), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I112 (.O(clk_m__L3_N112), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I111 (.O(clk_m__L3_N111), 
	.I(clk_m__L2_N11));
   BUFCKHHD clk_m__L3_I110 (.O(clk_m__L3_N110), 
	.I(clk_m__L2_N11));
   BUFCKHHD clk_m__L3_I109 (.O(clk_m__L3_N109), 
	.I(clk_m__L2_N11));
   BUFCKHHD clk_m__L3_I108 (.O(clk_m__L3_N108), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I107 (.O(clk_m__L3_N107), 
	.I(clk_m__L2_N10));
   BUFCKGHD clk_m__L3_I106 (.O(clk_m__L3_N106), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I105 (.O(clk_m__L3_N105), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I104 (.O(clk_m__L3_N104), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I103 (.O(clk_m__L3_N103), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I102 (.O(clk_m__L3_N102), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I101 (.O(clk_m__L3_N101), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I100 (.O(clk_m__L3_N100), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I99 (.O(clk_m__L3_N99), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I98 (.O(clk_m__L3_N98), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I97 (.O(clk_m__L3_N97), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I96 (.O(clk_m__L3_N96), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I95 (.O(clk_m__L3_N95), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I94 (.O(clk_m__L3_N94), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I93 (.O(clk_m__L3_N93), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I92 (.O(clk_m__L3_N92), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I91 (.O(clk_m__L3_N91), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I90 (.O(clk_m__L3_N90), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I89 (.O(clk_m__L3_N89), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I88 (.O(clk_m__L3_N88), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I87 (.O(clk_m__L3_N87), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I86 (.O(clk_m__L3_N86), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I85 (.O(clk_m__L3_N85), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I84 (.O(clk_m__L3_N84), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I83 (.O(clk_m__L3_N83), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I82 (.O(clk_m__L3_N82), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I81 (.O(clk_m__L3_N81), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I80 (.O(clk_m__L3_N80), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I79 (.O(clk_m__L3_N79), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I78 (.O(clk_m__L3_N78), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I77 (.O(clk_m__L3_N77), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I76 (.O(clk_m__L3_N76), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I75 (.O(clk_m__L3_N75), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I74 (.O(clk_m__L3_N74), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I73 (.O(clk_m__L3_N73), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I72 (.O(clk_m__L3_N72), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I71 (.O(clk_m__L3_N71), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I70 (.O(clk_m__L3_N70), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I69 (.O(clk_m__L3_N69), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I68 (.O(clk_m__L3_N68), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I67 (.O(clk_m__L3_N67), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I66 (.O(clk_m__L3_N66), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I65 (.O(clk_m__L3_N65), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I64 (.O(clk_m__L3_N64), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I63 (.O(clk_m__L3_N63), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I62 (.O(clk_m__L3_N62), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I61 (.O(clk_m__L3_N61), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I60 (.O(clk_m__L3_N60), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I59 (.O(clk_m__L3_N59), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I58 (.O(clk_m__L3_N58), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I57 (.O(clk_m__L3_N57), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I56 (.O(clk_m__L3_N56), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I55 (.O(clk_m__L3_N55), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I54 (.O(clk_m__L3_N54), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I53 (.O(clk_m__L3_N53), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I52 (.O(clk_m__L3_N52), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I51 (.O(clk_m__L3_N51), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I50 (.O(clk_m__L3_N50), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I49 (.O(clk_m__L3_N49), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I48 (.O(clk_m__L3_N48), 
	.I(clk_m__L2_N4));
   BUFCKGHD clk_m__L3_I47 (.O(clk_m__L3_N47), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I46 (.O(clk_m__L3_N46), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I45 (.O(clk_m__L3_N45), 
	.I(clk_m__L2_N4));
   BUFCKGHD clk_m__L3_I44 (.O(clk_m__L3_N44), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I43 (.O(clk_m__L3_N43), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I42 (.O(clk_m__L3_N42), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I41 (.O(clk_m__L3_N41), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I40 (.O(clk_m__L3_N40), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I39 (.O(clk_m__L3_N39), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I38 (.O(clk_m__L3_N38), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I37 (.O(clk_m__L3_N37), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I36 (.O(clk_m__L3_N36), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I35 (.O(clk_m__L3_N35), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I34 (.O(clk_m__L3_N34), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I33 (.O(clk_m__L3_N33), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I32 (.O(clk_m__L3_N32), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I31 (.O(clk_m__L3_N31), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I30 (.O(clk_m__L3_N30), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I29 (.O(clk_m__L3_N29), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I28 (.O(clk_m__L3_N28), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I27 (.O(clk_m__L3_N27), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I26 (.O(clk_m__L3_N26), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I25 (.O(clk_m__L3_N25), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I24 (.O(clk_m__L3_N24), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I23 (.O(clk_m__L3_N23), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I22 (.O(clk_m__L3_N22), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I21 (.O(clk_m__L3_N21), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I20 (.O(clk_m__L3_N20), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I19 (.O(clk_m__L3_N19), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I18 (.O(clk_m__L3_N18), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I17 (.O(clk_m__L3_N17), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I16 (.O(clk_m__L3_N16), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I15 (.O(clk_m__L3_N15), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I14 (.O(clk_m__L3_N14), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I13 (.O(clk_m__L3_N13), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I12 (.O(clk_m__L3_N12), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I11 (.O(clk_m__L3_N11), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I10 (.O(clk_m__L3_N10), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I9 (.O(clk_m__L3_N9), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I8 (.O(clk_m__L3_N8), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I7 (.O(clk_m__L3_N7), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I6 (.O(clk_m__L3_N6), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I5 (.O(clk_m__L3_N5), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I4 (.O(clk_m__L3_N4), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I3 (.O(clk_m__L3_N3), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I2 (.O(clk_m__L3_N2), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I1 (.O(clk_m__L3_N1), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I0 (.O(clk_m__L3_N0), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L2_I17 (.O(clk_m__L2_N17), 
	.I(clk_m__L1_N5));
   BUFCKHHD clk_m__L2_I16 (.O(clk_m__L2_N16), 
	.I(clk_m__L1_N5));
   BUFCKHHD clk_m__L2_I15 (.O(clk_m__L2_N15), 
	.I(clk_m__L1_N5));
   BUFCKHHD clk_m__L2_I14 (.O(clk_m__L2_N14), 
	.I(clk_m__L1_N4));
   BUFCKHHD clk_m__L2_I13 (.O(clk_m__L2_N13), 
	.I(clk_m__L1_N4));
   BUFCKHHD clk_m__L2_I12 (.O(clk_m__L2_N12), 
	.I(clk_m__L1_N4));
   BUFCKHHD clk_m__L2_I11 (.O(clk_m__L2_N11), 
	.I(clk_m__L1_N3));
   BUFCKHHD clk_m__L2_I10 (.O(clk_m__L2_N10), 
	.I(clk_m__L1_N3));
   BUFCKHHD clk_m__L2_I9 (.O(clk_m__L2_N9), 
	.I(clk_m__L1_N3));
   BUFCKHHD clk_m__L2_I8 (.O(clk_m__L2_N8), 
	.I(clk_m__L1_N2));
   BUFCKHHD clk_m__L2_I7 (.O(clk_m__L2_N7), 
	.I(clk_m__L1_N2));
   BUFCKHHD clk_m__L2_I6 (.O(clk_m__L2_N6), 
	.I(clk_m__L1_N2));
   BUFCKHHD clk_m__L2_I5 (.O(clk_m__L2_N5), 
	.I(clk_m__L1_N1));
   BUFCKHHD clk_m__L2_I4 (.O(clk_m__L2_N4), 
	.I(clk_m__L1_N1));
   BUFCKHHD clk_m__L2_I3 (.O(clk_m__L2_N3), 
	.I(clk_m__L1_N1));
   BUFCKHHD clk_m__L2_I2 (.O(clk_m__L2_N2), 
	.I(clk_m__L1_N0));
   BUFCKHHD clk_m__L2_I1 (.O(clk_m__L2_N1), 
	.I(clk_m__L1_N0));
   BUFCKHHD clk_m__L2_I0 (.O(clk_m__L2_N0), 
	.I(clk_m__L1_N0));
   BUFCKHHD clk_m__L1_I5 (.O(clk_m__L1_N5), 
	.I(clk_m));
   BUFCKGHD clk_m__L1_I4 (.O(clk_m__L1_N4), 
	.I(clk_m));
   BUFCKHHD clk_m__L1_I3 (.O(clk_m__L1_N3), 
	.I(clk_m));
   BUFCKHHD clk_m__L1_I2 (.O(clk_m__L1_N2), 
	.I(clk_m));
   BUFCKGHD clk_m__L1_I1 (.O(clk_m__L1_N1), 
	.I(clk_m));
   BUFCKHHD clk_m__L1_I0 (.O(clk_m__L1_N0), 
	.I(clk_m));
   BUFCKIHD FE_OFC96_n1 (.O(FE_OFN96_n1), 
	.I(n1));
   XMHA in1 (.SMT(n1), 
	.PU(n1), 
	.PD(n1), 
	.O(clk_m), 
	.I(clk));
   XMHA in2 (.SMT(n1), 
	.PU(n1), 
	.PD(n1), 
	.O(reset_m), 
	.I(reset));
   YA28SHA out1 (.SR(n1), 
	.O(pc_out[0]), 
	.I(pc_out_m[0]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out2 (.SR(n1), 
	.O(pc_out[1]), 
	.I(pc_out_m[1]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out3 (.SR(n1), 
	.O(pc_out[2]), 
	.I(pc_out_m[2]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out4 (.SR(n1), 
	.O(pc_out[3]), 
	.I(pc_out_m[3]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out5 (.SR(n1), 
	.O(pc_out[4]), 
	.I(pc_out_m[4]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out6 (.SR(FE_OFN96_n1), 
	.O(pc_out[5]), 
	.I(pc_out_m[5]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out7 (.SR(FE_OFN96_n1), 
	.O(pc_out[6]), 
	.I(pc_out_m[6]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out8 (.SR(n1), 
	.O(pc_out[7]), 
	.I(pc_out_m[7]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out9 (.SR(n1), 
	.O(pc_out[8]), 
	.I(pc_out_m[8]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out10 (.SR(n1), 
	.O(pc_out[9]), 
	.I(pc_out_m[9]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out11 (.SR(n1), 
	.O(pc_out[10]), 
	.I(pc_out_m[10]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out12 (.SR(n1), 
	.O(pc_out[11]), 
	.I(pc_out_m[11]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out13 (.SR(n1), 
	.O(pc_out[12]), 
	.I(pc_out_m[12]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out14 (.SR(n1), 
	.O(pc_out[13]), 
	.I(pc_out_m[13]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out15 (.SR(n1), 
	.O(pc_out[14]), 
	.I(pc_out_m[14]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out16 (.SR(n1), 
	.O(pc_out[15]), 
	.I(pc_out_m[15]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out17 (.SR(n1), 
	.O(alu_result[0]), 
	.I(alu_result_m[0]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out18 (.SR(n1), 
	.O(alu_result[1]), 
	.I(alu_result_m[1]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out19 (.SR(n1), 
	.O(alu_result[2]), 
	.I(alu_result_m[2]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out20 (.SR(n1), 
	.O(alu_result[3]), 
	.I(alu_result_m[3]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out21 (.SR(n1), 
	.O(alu_result[4]), 
	.I(alu_result_m[4]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out22 (.SR(n1), 
	.O(alu_result[5]), 
	.I(alu_result_m[5]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out23 (.SR(FE_OFN96_n1), 
	.O(alu_result[6]), 
	.I(alu_result_m[6]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out24 (.SR(FE_OFN96_n1), 
	.O(alu_result[7]), 
	.I(alu_result_m[7]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out25 (.SR(FE_OFN96_n1), 
	.O(alu_result[8]), 
	.I(alu_result_m[8]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out26 (.SR(FE_OFN96_n1), 
	.O(alu_result[9]), 
	.I(alu_result_m[9]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out27 (.SR(FE_OFN96_n1), 
	.O(alu_result[10]), 
	.I(alu_result_m[10]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out28 (.SR(FE_OFN96_n1), 
	.O(alu_result[11]), 
	.I(alu_result_m[11]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out29 (.SR(FE_OFN96_n1), 
	.O(alu_result[12]), 
	.I(alu_result_m[12]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out30 (.SR(FE_OFN96_n1), 
	.O(alu_result[13]), 
	.I(alu_result_m[13]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out31 (.SR(FE_OFN96_n1), 
	.O(alu_result[14]), 
	.I(alu_result_m[14]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out32 (.SR(FE_OFN96_n1), 
	.O(alu_result[15]), 
	.I(alu_result_m[15]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   VCCKHA pwr_1 (.VCC(vdd));
   VCCKHA pwr_2 (.VCC(vdd));
   VCCKHA pwr_3 (.VCC(vdd));
   VCCKHA pwr_4 (.VCC(vdd));
   VCC3IHA pwr_5 (.VCC3I(vddio));
   VCC3IHA pwr_6 (.VCC3I(vddio));
   VCC3IHA pwr_7 (.VCC3I(vddio));
   VCC3IHA pwr_8 (.VCC3I(vddio));
   GND3IHA gnd_1 (.GND3I(vss));
   GND3IHA gnd_2 (.GND3I(vss));
   GND3IHA gnd_3 (.GND3I(vss));
   GND3IHA gnd_4 (.GND3I(vss));
   GNDKHA gnd_5 (.GND(gnd));
   GNDKHA gnd_6 (.GND(gnd));
   GNDKHA gnd_7 (.GND(gnd));
   GNDKHA gnd_8 (.GND(gnd));
   CORNERHA corner_1 ();
   CORNERHA corner_2 ();
   CORNERHA corner_3 ();
   CORNERHA corner_4 ();
   mips_16 mips_core (.clk(clk_m__L3_N0), 
	.reset(reset_m), 
	.pc_out({ pc_out_m[15],
		pc_out_m[14],
		pc_out_m[13],
		pc_out_m[12],
		pc_out_m[11],
		pc_out_m[10],
		pc_out_m[9],
		pc_out_m[8],
		pc_out_m[7],
		pc_out_m[6],
		pc_out_m[5],
		pc_out_m[4],
		pc_out_m[3],
		pc_out_m[2],
		pc_out_m[1],
		pc_out_m[0] }), 
	.alu_result({ alu_result_m[15],
		alu_result_m[14],
		alu_result_m[13],
		alu_result_m[12],
		alu_result_m[11],
		alu_result_m[10],
		alu_result_m[9],
		alu_result_m[8],
		alu_result_m[7],
		alu_result_m[6],
		alu_result_m[5],
		alu_result_m[4],
		alu_result_m[3],
		alu_result_m[2],
		alu_result_m[1],
		alu_result_m[0] }), 
	.clk_m__L3_N1(clk_m__L3_N1), 
	.clk_m__L3_N10(clk_m__L3_N10), 
	.clk_m__L3_N100(clk_m__L3_N100), 
	.clk_m__L3_N101(clk_m__L3_N101), 
	.clk_m__L3_N102(clk_m__L3_N102), 
	.clk_m__L3_N103(clk_m__L3_N103), 
	.clk_m__L3_N104(clk_m__L3_N104), 
	.clk_m__L3_N105(clk_m__L3_N105), 
	.clk_m__L3_N106(clk_m__L3_N106), 
	.clk_m__L3_N107(clk_m__L3_N107), 
	.clk_m__L3_N108(clk_m__L3_N108), 
	.clk_m__L3_N109(clk_m__L3_N109), 
	.clk_m__L3_N11(clk_m__L3_N11), 
	.clk_m__L3_N110(clk_m__L3_N110), 
	.clk_m__L3_N111(clk_m__L3_N111), 
	.clk_m__L3_N112(clk_m__L3_N112), 
	.clk_m__L3_N113(clk_m__L3_N113), 
	.clk_m__L3_N114(clk_m__L3_N114), 
	.clk_m__L3_N115(clk_m__L3_N115), 
	.clk_m__L3_N116(clk_m__L3_N116), 
	.clk_m__L3_N117(clk_m__L3_N117), 
	.clk_m__L3_N118(clk_m__L3_N118), 
	.clk_m__L3_N119(clk_m__L3_N119), 
	.clk_m__L3_N12(clk_m__L3_N12), 
	.clk_m__L3_N120(clk_m__L3_N120), 
	.clk_m__L3_N121(clk_m__L3_N121), 
	.clk_m__L3_N122(clk_m__L3_N122), 
	.clk_m__L3_N123(clk_m__L3_N123), 
	.clk_m__L3_N124(clk_m__L3_N124), 
	.clk_m__L3_N125(clk_m__L3_N125), 
	.clk_m__L3_N126(clk_m__L3_N126), 
	.clk_m__L3_N127(clk_m__L3_N127), 
	.clk_m__L3_N128(clk_m__L3_N128), 
	.clk_m__L3_N129(clk_m__L3_N129), 
	.clk_m__L3_N13(clk_m__L3_N13), 
	.clk_m__L3_N130(clk_m__L3_N130), 
	.clk_m__L3_N131(clk_m__L3_N131), 
	.clk_m__L3_N132(clk_m__L3_N132), 
	.clk_m__L3_N133(clk_m__L3_N133), 
	.clk_m__L3_N134(clk_m__L3_N134), 
	.clk_m__L3_N135(clk_m__L3_N135), 
	.clk_m__L3_N136(clk_m__L3_N136), 
	.clk_m__L3_N137(clk_m__L3_N137), 
	.clk_m__L3_N138(clk_m__L3_N138), 
	.clk_m__L3_N139(clk_m__L3_N139), 
	.clk_m__L3_N14(clk_m__L3_N14), 
	.clk_m__L3_N140(clk_m__L3_N140), 
	.clk_m__L3_N141(clk_m__L3_N141), 
	.clk_m__L3_N142(clk_m__L3_N142), 
	.clk_m__L3_N143(clk_m__L3_N143), 
	.clk_m__L3_N144(clk_m__L3_N144), 
	.clk_m__L3_N145(clk_m__L3_N145), 
	.clk_m__L3_N146(clk_m__L3_N146), 
	.clk_m__L3_N147(clk_m__L3_N147), 
	.clk_m__L3_N148(clk_m__L3_N148), 
	.clk_m__L3_N149(clk_m__L3_N149), 
	.clk_m__L3_N15(clk_m__L3_N15), 
	.clk_m__L3_N150(clk_m__L3_N150), 
	.clk_m__L3_N151(clk_m__L3_N151), 
	.clk_m__L3_N152(clk_m__L3_N152), 
	.clk_m__L3_N153(clk_m__L3_N153), 
	.clk_m__L3_N154(clk_m__L3_N154), 
	.clk_m__L3_N155(clk_m__L3_N155), 
	.clk_m__L3_N156(clk_m__L3_N156), 
	.clk_m__L3_N157(clk_m__L3_N157), 
	.clk_m__L3_N158(clk_m__L3_N158), 
	.clk_m__L3_N159(clk_m__L3_N159), 
	.clk_m__L3_N16(clk_m__L3_N16), 
	.clk_m__L3_N160(clk_m__L3_N160), 
	.clk_m__L3_N161(clk_m__L3_N161), 
	.clk_m__L3_N162(clk_m__L3_N162), 
	.clk_m__L3_N163(clk_m__L3_N163), 
	.clk_m__L3_N164(clk_m__L3_N164), 
	.clk_m__L3_N165(clk_m__L3_N165), 
	.clk_m__L3_N166(clk_m__L3_N166), 
	.clk_m__L3_N167(clk_m__L3_N167), 
	.clk_m__L3_N168(clk_m__L3_N168), 
	.clk_m__L3_N169(clk_m__L3_N169), 
	.clk_m__L3_N17(clk_m__L3_N17), 
	.clk_m__L3_N170(clk_m__L3_N170), 
	.clk_m__L3_N171(clk_m__L3_N171), 
	.clk_m__L3_N172(clk_m__L3_N172), 
	.clk_m__L3_N173(clk_m__L3_N173), 
	.clk_m__L3_N174(clk_m__L3_N174), 
	.clk_m__L3_N175(clk_m__L3_N175), 
	.clk_m__L3_N176(clk_m__L3_N176), 
	.clk_m__L3_N177(clk_m__L3_N177), 
	.clk_m__L3_N18(clk_m__L3_N18), 
	.clk_m__L3_N19(clk_m__L3_N19), 
	.clk_m__L3_N2(clk_m__L3_N2), 
	.clk_m__L3_N20(clk_m__L3_N20), 
	.clk_m__L3_N21(clk_m__L3_N21), 
	.clk_m__L3_N22(clk_m__L3_N22), 
	.clk_m__L3_N23(clk_m__L3_N23), 
	.clk_m__L3_N24(clk_m__L3_N24), 
	.clk_m__L3_N25(clk_m__L3_N25), 
	.clk_m__L3_N26(clk_m__L3_N26), 
	.clk_m__L3_N27(clk_m__L3_N27), 
	.clk_m__L3_N28(clk_m__L3_N28), 
	.clk_m__L3_N29(clk_m__L3_N29), 
	.clk_m__L3_N3(clk_m__L3_N3), 
	.clk_m__L3_N30(clk_m__L3_N30), 
	.clk_m__L3_N31(clk_m__L3_N31), 
	.clk_m__L3_N32(clk_m__L3_N32), 
	.clk_m__L3_N33(clk_m__L3_N33), 
	.clk_m__L3_N34(clk_m__L3_N34), 
	.clk_m__L3_N35(clk_m__L3_N35), 
	.clk_m__L3_N36(clk_m__L3_N36), 
	.clk_m__L3_N37(clk_m__L3_N37), 
	.clk_m__L3_N38(clk_m__L3_N38), 
	.clk_m__L3_N39(clk_m__L3_N39), 
	.clk_m__L3_N4(clk_m__L3_N4), 
	.clk_m__L3_N40(clk_m__L3_N40), 
	.clk_m__L3_N41(clk_m__L3_N41), 
	.clk_m__L3_N42(clk_m__L3_N42), 
	.clk_m__L3_N43(clk_m__L3_N43), 
	.clk_m__L3_N44(clk_m__L3_N44), 
	.clk_m__L3_N45(clk_m__L3_N45), 
	.clk_m__L3_N46(clk_m__L3_N46), 
	.clk_m__L3_N47(clk_m__L3_N47), 
	.clk_m__L3_N48(clk_m__L3_N48), 
	.clk_m__L3_N49(clk_m__L3_N49), 
	.clk_m__L3_N5(clk_m__L3_N5), 
	.clk_m__L3_N50(clk_m__L3_N50), 
	.clk_m__L3_N51(clk_m__L3_N51), 
	.clk_m__L3_N52(clk_m__L3_N52), 
	.clk_m__L3_N53(clk_m__L3_N53), 
	.clk_m__L3_N54(clk_m__L3_N54), 
	.clk_m__L3_N55(clk_m__L3_N55), 
	.clk_m__L3_N56(clk_m__L3_N56), 
	.clk_m__L3_N57(clk_m__L3_N57), 
	.clk_m__L3_N58(clk_m__L3_N58), 
	.clk_m__L3_N59(clk_m__L3_N59), 
	.clk_m__L3_N6(clk_m__L3_N6), 
	.clk_m__L3_N60(clk_m__L3_N60), 
	.clk_m__L3_N61(clk_m__L3_N61), 
	.clk_m__L3_N62(clk_m__L3_N62), 
	.clk_m__L3_N63(clk_m__L3_N63), 
	.clk_m__L3_N64(clk_m__L3_N64), 
	.clk_m__L3_N65(clk_m__L3_N65), 
	.clk_m__L3_N66(clk_m__L3_N66), 
	.clk_m__L3_N67(clk_m__L3_N67), 
	.clk_m__L3_N68(clk_m__L3_N68), 
	.clk_m__L3_N69(clk_m__L3_N69), 
	.clk_m__L3_N7(clk_m__L3_N7), 
	.clk_m__L3_N70(clk_m__L3_N70), 
	.clk_m__L3_N71(clk_m__L3_N71), 
	.clk_m__L3_N72(clk_m__L3_N72), 
	.clk_m__L3_N73(clk_m__L3_N73), 
	.clk_m__L3_N74(clk_m__L3_N74), 
	.clk_m__L3_N75(clk_m__L3_N75), 
	.clk_m__L3_N76(clk_m__L3_N76), 
	.clk_m__L3_N77(clk_m__L3_N77), 
	.clk_m__L3_N78(clk_m__L3_N78), 
	.clk_m__L3_N79(clk_m__L3_N79), 
	.clk_m__L3_N8(clk_m__L3_N8), 
	.clk_m__L3_N80(clk_m__L3_N80), 
	.clk_m__L3_N81(clk_m__L3_N81), 
	.clk_m__L3_N82(clk_m__L3_N82), 
	.clk_m__L3_N83(clk_m__L3_N83), 
	.clk_m__L3_N84(clk_m__L3_N84), 
	.clk_m__L3_N85(clk_m__L3_N85), 
	.clk_m__L3_N86(clk_m__L3_N86), 
	.clk_m__L3_N87(clk_m__L3_N87), 
	.clk_m__L3_N88(clk_m__L3_N88), 
	.clk_m__L3_N89(clk_m__L3_N89), 
	.clk_m__L3_N9(clk_m__L3_N9), 
	.clk_m__L3_N90(clk_m__L3_N90), 
	.clk_m__L3_N91(clk_m__L3_N91), 
	.clk_m__L3_N92(clk_m__L3_N92), 
	.clk_m__L3_N93(clk_m__L3_N93), 
	.clk_m__L3_N94(clk_m__L3_N94), 
	.clk_m__L3_N95(clk_m__L3_N95), 
	.clk_m__L3_N96(clk_m__L3_N96), 
	.clk_m__L3_N97(clk_m__L3_N97), 
	.clk_m__L3_N98(clk_m__L3_N98), 
	.clk_m__L3_N99(clk_m__L3_N99), 
	.clk_m__N0(clk_m__N0));
   TIE1DHD U3 (.O(n2));
   TIE0DHD U4 (.O(n1));
endmodule

