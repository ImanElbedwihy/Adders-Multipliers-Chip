/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May  5 23:55:48 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2065577432 */

/* blackbox module full_adder_bbox__0_12 */

/* blackbox module full_adder_bbox_0__0_11 */

/* blackbox module full_adder_bbox_1__0_10 */

/* blackbox module full_adder_bbox_2__0_9 */

module four_bit_adder__0_13(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_12 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(Cin), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_11 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_10 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_9 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_17 */

/* blackbox module full_adder_bbox_0__0_16 */

/* blackbox module full_adder_bbox_1__0_15 */

/* blackbox module full_adder_bbox_2__0_14 */

module four_bit_adder__0_18(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_17 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b0), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_16 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_15 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_14 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_22 */

/* blackbox module full_adder_bbox_0__0_21 */

/* blackbox module full_adder_bbox_1__0_20 */

/* blackbox module full_adder_bbox_2__0_19 */

module four_bit_adder__0_23(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_22 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b1), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_21 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_20 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_19 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_27 */

/* blackbox module full_adder_bbox_0__0_26 */

/* blackbox module full_adder_bbox_1__0_25 */

/* blackbox module full_adder_bbox_2__0_24 */

module four_bit_adder__0_28(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_27 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b0), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_26 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_25 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_24 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_32 */

/* blackbox module full_adder_bbox_0__0_31 */

/* blackbox module full_adder_bbox_1__0_30 */

/* blackbox module full_adder_bbox_2__0_29 */

module four_bit_adder__0_33(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_32 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b1), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_31 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_30 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_29 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_37 */

/* blackbox module full_adder_bbox_0__0_36 */

/* blackbox module full_adder_bbox_1__0_35 */

/* blackbox module full_adder_bbox_2__0_34 */

module four_bit_adder__0_38(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_37 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b0), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_36 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_35 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_34 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_42 */

/* blackbox module full_adder_bbox_0__0_41 */

/* blackbox module full_adder_bbox_1__0_40 */

/* blackbox module full_adder_bbox_2__0_39 */

module four_bit_adder__0_43(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_42 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b1), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_41 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_40 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_39 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_47 */

/* blackbox module full_adder_bbox_0__0_46 */

/* blackbox module full_adder_bbox_1__0_45 */

/* blackbox module full_adder_bbox_2__0_44 */

module four_bit_adder__0_48(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_47 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b0), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_46 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_45 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_44 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_52 */

/* blackbox module full_adder_bbox_0__0_51 */

/* blackbox module full_adder_bbox_1__0_50 */

/* blackbox module full_adder_bbox_2__0_49 */

module four_bit_adder__0_53(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_52 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b1), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_51 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_50 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_49 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_57 */

/* blackbox module full_adder_bbox_0__0_56 */

/* blackbox module full_adder_bbox_1__0_55 */

/* blackbox module full_adder_bbox_2__0_54 */

module four_bit_adder__0_58(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_57 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b0), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_56 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_55 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_54 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_62 */

/* blackbox module full_adder_bbox_0__0_61 */

/* blackbox module full_adder_bbox_1__0_60 */

/* blackbox module full_adder_bbox_2__0_59 */

module four_bit_adder__0_63(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_62 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b1), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_61 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_60 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_59 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_67 */

/* blackbox module full_adder_bbox_0__0_66 */

/* blackbox module full_adder_bbox_1__0_65 */

/* blackbox module full_adder_bbox_2__0_64 */

module four_bit_adder__0_68(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_67 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b0), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_66 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_65 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_64 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_72 */

/* blackbox module full_adder_bbox_0__0_71 */

/* blackbox module full_adder_bbox_1__0_70 */

/* blackbox module full_adder_bbox_2__0_69 */

module four_bit_adder__0_73(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_72 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b1), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_71 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_70 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_69 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox__0_77 */

/* blackbox module full_adder_bbox_0__0_76 */

/* blackbox module full_adder_bbox_1__0_75 */

/* blackbox module full_adder_bbox_2__0_74 */

module four_bit_adder__0_78(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox__0_77 loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b0), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0__0_76 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1__0_75 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2__0_74 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

/* blackbox module full_adder_bbox */

/* blackbox module full_adder_bbox_0 */

/* blackbox module full_adder_bbox_1 */

/* blackbox module full_adder_bbox_2 */

module four_bit_adder(A, B, Cin, Sum, Cout);
   input [3:0]A;
   input [3:0]B;
   input Cin;
   output [3:0]Sum;
   output Cout;

   full_adder_bbox loop_0_FA (.i_bit1(A[0]), .i_bit2(B[0]), .i_carry(1'b1), 
      .o_sum(Sum[0]), .o_carry(n_0));
   full_adder_bbox_0 loop_1_FA (.i_bit1(A[1]), .i_bit2(B[1]), .i_carry(n_0), 
      .o_sum(Sum[1]), .o_carry(n_1));
   full_adder_bbox_1 loop_2_FA (.i_bit1(A[2]), .i_bit2(B[2]), .i_carry(n_1), 
      .o_sum(Sum[2]), .o_carry(n_2));
   full_adder_bbox_2 loop_3_FA (.i_bit1(A[3]), .i_bit2(B[3]), .i_carry(n_2), 
      .o_sum(Sum[3]), .o_carry(Cout));
endmodule

module CSA(A, B, Cin, Sum, Cout, Overflow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]Sum;
   output Cout;
   output Overflow;

   wire C;
   wire C0;
   wire C1;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;

   four_bit_adder__0_13 A_inst (.A({A[3], A[2], A[1], A[0]}), .B({B[3], B[2], 
      B[1], B[0]}), .Cin(Cin), .Sum({Sum[3], Sum[2], Sum[1], Sum[0]}), .Cout(C));
   four_bit_adder__0_18 loop1_6_A0 (.A({A[31], A[30], A[29], A[28]}), .B({B[31], 
      B[30], B[29], B[28]}), .Cin(), .Sum({n_3, n_2, n_1, n_0}), .Cout(C0));
   four_bit_adder__0_23 loop1_6_A1 (.A({A[31], A[30], A[29], A[28]}), .B({B[31], 
      B[30], B[29], B[28]}), .Cin(), .Sum({n_7, n_6, n_5, n_4}), .Cout(C1));
   four_bit_adder__0_28 loop1_5_A0 (.A({A[27], A[26], A[25], A[24]}), .B({B[27], 
      B[26], B[25], B[24]}), .Cin(), .Sum({n_12, n_11, n_10, n_9}), .Cout(n_8));
   four_bit_adder__0_33 loop1_5_A1 (.A({A[27], A[26], A[25], A[24]}), .B({B[27], 
      B[26], B[25], B[24]}), .Cin(), .Sum({n_17, n_16, n_15, n_14}), .Cout(n_13));
   four_bit_adder__0_38 loop1_4_A0 (.A({A[23], A[22], A[21], A[20]}), .B({B[23], 
      B[22], B[21], B[20]}), .Cin(), .Sum({n_22, n_21, n_20, n_19}), .Cout(n_18));
   four_bit_adder__0_43 loop1_4_A1 (.A({A[23], A[22], A[21], A[20]}), .B({B[23], 
      B[22], B[21], B[20]}), .Cin(), .Sum({n_27, n_26, n_25, n_24}), .Cout(n_23));
   four_bit_adder__0_48 loop1_3_A0 (.A({A[19], A[18], A[17], A[16]}), .B({B[19], 
      B[18], B[17], B[16]}), .Cin(), .Sum({n_32, n_31, n_30, n_29}), .Cout(n_28));
   four_bit_adder__0_53 loop1_3_A1 (.A({A[19], A[18], A[17], A[16]}), .B({B[19], 
      B[18], B[17], B[16]}), .Cin(), .Sum({n_37, n_36, n_35, n_34}), .Cout(n_33));
   four_bit_adder__0_58 loop1_2_A0 (.A({A[15], A[14], A[13], A[12]}), .B({B[15], 
      B[14], B[13], B[12]}), .Cin(), .Sum({n_42, n_41, n_40, n_39}), .Cout(n_38));
   four_bit_adder__0_63 loop1_2_A1 (.A({A[15], A[14], A[13], A[12]}), .B({B[15], 
      B[14], B[13], B[12]}), .Cin(), .Sum({n_47, n_46, n_45, n_44}), .Cout(n_43));
   four_bit_adder__0_68 loop1_1_A0 (.A({A[11], A[10], A[9], A[8]}), .B({B[11], 
      B[10], B[9], B[8]}), .Cin(), .Sum({n_52, n_51, n_50, n_49}), .Cout(n_48));
   four_bit_adder__0_73 loop1_1_A1 (.A({A[11], A[10], A[9], A[8]}), .B({B[11], 
      B[10], B[9], B[8]}), .Cin(), .Sum({n_57, n_56, n_55, n_54}), .Cout(n_53));
   four_bit_adder__0_78 loop1_0_A0 (.A({A[7], A[6], A[5], A[4]}), .B({B[7], B[6], 
      B[5], B[4]}), .Cin(), .Sum({n_62, n_61, n_60, n_59}), .Cout(n_58));
   four_bit_adder loop1_0_A1 (.A({A[7], A[6], A[5], A[4]}), .B({B[7], B[6], B[5], 
      B[4]}), .Cin(), .Sum({n_67, n_66, n_65, n_64}), .Cout(n_63));
   MUX2_X1_LVT i_0_0_0 (.A(C0), .B(C1), .S(n_0_0_3), .Z(Cout));
   OAI21_X1_LVT i_0_0_1 (.A(n_0_0_0), .B1(n_0_0_1), .B2(Sum[31]), .ZN(Overflow));
   NAND2_X1_LVT i_0_0_2 (.A1(Sum[31]), .A2(n_0_0_2), .ZN(n_0_0_0));
   NAND2_X1_LVT i_0_0_3 (.A1(A[31]), .A2(B[31]), .ZN(n_0_0_1));
   NOR2_X1_LVT i_0_0_4 (.A1(A[31]), .A2(B[31]), .ZN(n_0_0_2));
   MUX2_X1_LVT i_0_0_5 (.A(n_59), .B(n_64), .S(C), .Z(Sum[4]));
   MUX2_X1_LVT i_0_0_6 (.A(n_60), .B(n_65), .S(C), .Z(Sum[5]));
   MUX2_X1_LVT i_0_0_7 (.A(n_61), .B(n_66), .S(C), .Z(Sum[6]));
   MUX2_X1_LVT i_0_0_8 (.A(n_62), .B(n_67), .S(C), .Z(Sum[7]));
   MUX2_X1_LVT i_0_0_9 (.A(n_49), .B(n_54), .S(n_0_0_8), .Z(Sum[8]));
   MUX2_X1_LVT i_0_0_10 (.A(n_50), .B(n_55), .S(n_0_0_8), .Z(Sum[9]));
   MUX2_X1_LVT i_0_0_11 (.A(n_51), .B(n_56), .S(n_0_0_8), .Z(Sum[10]));
   MUX2_X1_LVT i_0_0_12 (.A(n_52), .B(n_57), .S(n_0_0_8), .Z(Sum[11]));
   MUX2_X1_LVT i_0_0_13 (.A(n_39), .B(n_44), .S(n_0_0_7), .Z(Sum[12]));
   MUX2_X1_LVT i_0_0_14 (.A(n_40), .B(n_45), .S(n_0_0_7), .Z(Sum[13]));
   MUX2_X1_LVT i_0_0_15 (.A(n_41), .B(n_46), .S(n_0_0_7), .Z(Sum[14]));
   MUX2_X1_LVT i_0_0_16 (.A(n_42), .B(n_47), .S(n_0_0_7), .Z(Sum[15]));
   MUX2_X1_LVT i_0_0_17 (.A(n_29), .B(n_34), .S(n_0_0_6), .Z(Sum[16]));
   MUX2_X1_LVT i_0_0_18 (.A(n_30), .B(n_35), .S(n_0_0_6), .Z(Sum[17]));
   MUX2_X1_LVT i_0_0_19 (.A(n_31), .B(n_36), .S(n_0_0_6), .Z(Sum[18]));
   MUX2_X1_LVT i_0_0_20 (.A(n_32), .B(n_37), .S(n_0_0_6), .Z(Sum[19]));
   MUX2_X1_LVT i_0_0_21 (.A(n_19), .B(n_24), .S(n_0_0_5), .Z(Sum[20]));
   MUX2_X1_LVT i_0_0_22 (.A(n_20), .B(n_25), .S(n_0_0_5), .Z(Sum[21]));
   MUX2_X1_LVT i_0_0_23 (.A(n_21), .B(n_26), .S(n_0_0_5), .Z(Sum[22]));
   MUX2_X1_LVT i_0_0_24 (.A(n_22), .B(n_27), .S(n_0_0_5), .Z(Sum[23]));
   MUX2_X1_LVT i_0_0_25 (.A(n_9), .B(n_14), .S(n_0_0_4), .Z(Sum[24]));
   MUX2_X1_LVT i_0_0_26 (.A(n_10), .B(n_15), .S(n_0_0_4), .Z(Sum[25]));
   MUX2_X1_LVT i_0_0_27 (.A(n_11), .B(n_16), .S(n_0_0_4), .Z(Sum[26]));
   MUX2_X1_LVT i_0_0_28 (.A(n_12), .B(n_17), .S(n_0_0_4), .Z(Sum[27]));
   MUX2_X1_LVT i_0_0_29 (.A(n_0), .B(n_4), .S(n_0_0_3), .Z(Sum[28]));
   MUX2_X1_LVT i_0_0_30 (.A(n_1), .B(n_5), .S(n_0_0_3), .Z(Sum[29]));
   MUX2_X1_LVT i_0_0_31 (.A(n_2), .B(n_6), .S(n_0_0_3), .Z(Sum[30]));
   MUX2_X1_LVT i_0_0_32 (.A(n_3), .B(n_7), .S(n_0_0_3), .Z(Sum[31]));
   MUX2_X1_LVT i_0_0_33 (.A(n_8), .B(n_13), .S(n_0_0_4), .Z(n_0_0_3));
   MUX2_X1_LVT i_0_0_34 (.A(n_18), .B(n_23), .S(n_0_0_5), .Z(n_0_0_4));
   MUX2_X1_LVT i_0_0_35 (.A(n_28), .B(n_33), .S(n_0_0_6), .Z(n_0_0_5));
   MUX2_X1_LVT i_0_0_36 (.A(n_38), .B(n_43), .S(n_0_0_7), .Z(n_0_0_6));
   MUX2_X1_LVT i_0_0_37 (.A(n_48), .B(n_53), .S(n_0_0_8), .Z(n_0_0_7));
   MUX2_X1_LVT i_0_0_38 (.A(n_58), .B(n_63), .S(C), .Z(n_0_0_8));
endmodule
