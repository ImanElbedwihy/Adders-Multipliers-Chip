module alu_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [15:0] A;
   input [15:0] B;
   input CI;
   output [15:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [15:1] carry;

   FA1DHD U1_0 (.S(SUM[0]), 
	.CO(carry[1]), 
	.CI(n1), 
	.B(B[0]), 
	.A(A[0]));
   FA1DHD U1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.CI(carry[1]), 
	.B(B[1]), 
	.A(A[1]));
   FA1DHD U1_13 (.S(SUM[13]), 
	.CO(carry[14]), 
	.CI(carry[13]), 
	.B(B[13]), 
	.A(A[13]));
   FA1DHD U1_11 (.S(SUM[11]), 
	.CO(carry[12]), 
	.CI(carry[11]), 
	.B(B[11]), 
	.A(A[11]));
   FA1DHD U1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.CI(carry[7]), 
	.B(B[7]), 
	.A(A[7]));
   FA1DHD U1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(B[5]), 
	.A(A[5]));
   FA1DHD U1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(B[3]), 
	.A(A[3]));
   FA1DHD U1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(B[2]), 
	.A(A[2]));
   FA1DHD U1_9 (.S(SUM[9]), 
	.CO(carry[10]), 
	.CI(carry[9]), 
	.B(B[9]), 
	.A(A[9]));
   FA1DHD U1_14 (.S(SUM[14]), 
	.CO(carry[15]), 
	.CI(carry[14]), 
	.B(B[14]), 
	.A(A[14]));
   FA1DHD U1_12 (.S(SUM[12]), 
	.CO(carry[13]), 
	.CI(carry[12]), 
	.B(B[12]), 
	.A(A[12]));
   FA1DHD U1_10 (.S(SUM[10]), 
	.CO(carry[11]), 
	.CI(carry[10]), 
	.B(B[10]), 
	.A(A[10]));
   FA1DHD U1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.CI(carry[8]), 
	.B(B[8]), 
	.A(A[8]));
   FA1DHD U1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(B[6]), 
	.A(A[6]));
   FA1DHD U1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(B[4]), 
	.A(A[4]));
   XOR3EHD U1_15 (.O(SUM[15]), 
	.I3(carry[15]), 
	.I2(B[15]), 
	.I1(A[15]));
   TIE0DHD U1 (.O(n1));
endmodule

module alu_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [15:0] A;
   input [15:0] B;
   input CI;
   output [15:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire [16:0] carry;

   FA1DHD U2_0 (.S(DIFF[0]), 
	.CO(carry[1]), 
	.CI(n17), 
	.B(n16), 
	.A(A[0]));
   FA1DHD U2_1 (.S(DIFF[1]), 
	.CO(carry[2]), 
	.CI(carry[1]), 
	.B(n15), 
	.A(A[1]));
   FA1DHD U2_13 (.S(DIFF[13]), 
	.CO(carry[14]), 
	.CI(carry[13]), 
	.B(n3), 
	.A(A[13]));
   FA1DHD U2_11 (.S(DIFF[11]), 
	.CO(carry[12]), 
	.CI(carry[11]), 
	.B(n5), 
	.A(A[11]));
   FA1DHD U2_7 (.S(DIFF[7]), 
	.CO(carry[8]), 
	.CI(carry[7]), 
	.B(n9), 
	.A(A[7]));
   FA1DHD U2_5 (.S(DIFF[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(n11), 
	.A(A[5]));
   FA1DHD U2_3 (.S(DIFF[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(n13), 
	.A(A[3]));
   FA1DHD U2_2 (.S(DIFF[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(n14), 
	.A(A[2]));
   FA1DHD U2_9 (.S(DIFF[9]), 
	.CO(carry[10]), 
	.CI(carry[9]), 
	.B(n7), 
	.A(A[9]));
   FA1DHD U2_14 (.S(DIFF[14]), 
	.CO(carry[15]), 
	.CI(carry[14]), 
	.B(n2), 
	.A(A[14]));
   FA1DHD U2_12 (.S(DIFF[12]), 
	.CO(carry[13]), 
	.CI(carry[12]), 
	.B(n4), 
	.A(A[12]));
   FA1DHD U2_10 (.S(DIFF[10]), 
	.CO(carry[11]), 
	.CI(carry[10]), 
	.B(n6), 
	.A(A[10]));
   FA1DHD U2_8 (.S(DIFF[8]), 
	.CO(carry[9]), 
	.CI(carry[8]), 
	.B(n8), 
	.A(A[8]));
   FA1DHD U2_6 (.S(DIFF[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(n10), 
	.A(A[6]));
   FA1DHD U2_4 (.S(DIFF[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(n12), 
	.A(A[4]));
   XOR3EHD U2_15 (.O(DIFF[15]), 
	.I3(carry[15]), 
	.I2(n1), 
	.I1(A[15]));
   INVDHD U1 (.O(n1), 
	.I(B[15]));
   INVDHD U2 (.O(n12), 
	.I(B[4]));
   INVDHD U3 (.O(n10), 
	.I(B[6]));
   INVDHD U4 (.O(n8), 
	.I(B[8]));
   INVDHD U5 (.O(n6), 
	.I(B[10]));
   INVDHD U6 (.O(n4), 
	.I(B[12]));
   INVDHD U7 (.O(n2), 
	.I(B[14]));
   INVDHD U8 (.O(n7), 
	.I(B[9]));
   INVDHD U9 (.O(n14), 
	.I(B[2]));
   INVDHD U10 (.O(n13), 
	.I(B[3]));
   INVDHD U11 (.O(n11), 
	.I(B[5]));
   INVDHD U12 (.O(n9), 
	.I(B[7]));
   INVDHD U13 (.O(n5), 
	.I(B[11]));
   INVDHD U14 (.O(n3), 
	.I(B[13]));
   INVDHD U15 (.O(n15), 
	.I(B[1]));
   INVDHD U16 (.O(n16), 
	.I(B[0]));
   TIE1DHD U17 (.O(n17));
endmodule

module data_memory (
	clk, 
	mem_access_addr, 
	mem_write_data, 
	mem_write_en, 
	mem_read, 
	mem_read_data, 
	clk_m__L3_N1, 
	clk_m__L3_N10, 
	clk_m__L3_N100, 
	clk_m__L3_N101, 
	clk_m__L3_N102, 
	clk_m__L3_N103, 
	clk_m__L3_N104, 
	clk_m__L3_N105, 
	clk_m__L3_N106, 
	clk_m__L3_N107, 
	clk_m__L3_N108, 
	clk_m__L3_N109, 
	clk_m__L3_N11, 
	clk_m__L3_N110, 
	clk_m__L3_N111, 
	clk_m__L3_N112, 
	clk_m__L3_N113, 
	clk_m__L3_N114, 
	clk_m__L3_N115, 
	clk_m__L3_N116, 
	clk_m__L3_N117, 
	clk_m__L3_N118, 
	clk_m__L3_N119, 
	clk_m__L3_N12, 
	clk_m__L3_N120, 
	clk_m__L3_N121, 
	clk_m__L3_N122, 
	clk_m__L3_N123, 
	clk_m__L3_N124, 
	clk_m__L3_N125, 
	clk_m__L3_N126, 
	clk_m__L3_N127, 
	clk_m__L3_N128, 
	clk_m__L3_N129, 
	clk_m__L3_N13, 
	clk_m__L3_N130, 
	clk_m__L3_N131, 
	clk_m__L3_N132, 
	clk_m__L3_N133, 
	clk_m__L3_N134, 
	clk_m__L3_N135, 
	clk_m__L3_N136, 
	clk_m__L3_N137, 
	clk_m__L3_N138, 
	clk_m__L3_N139, 
	clk_m__L3_N14, 
	clk_m__L3_N140, 
	clk_m__L3_N141, 
	clk_m__L3_N142, 
	clk_m__L3_N143, 
	clk_m__L3_N144, 
	clk_m__L3_N145, 
	clk_m__L3_N146, 
	clk_m__L3_N147, 
	clk_m__L3_N148, 
	clk_m__L3_N149, 
	clk_m__L3_N15, 
	clk_m__L3_N150, 
	clk_m__L3_N151, 
	clk_m__L3_N152, 
	clk_m__L3_N153, 
	clk_m__L3_N154, 
	clk_m__L3_N155, 
	clk_m__L3_N156, 
	clk_m__L3_N157, 
	clk_m__L3_N158, 
	clk_m__L3_N159, 
	clk_m__L3_N16, 
	clk_m__L3_N160, 
	clk_m__L3_N161, 
	clk_m__L3_N162, 
	clk_m__L3_N163, 
	clk_m__L3_N164, 
	clk_m__L3_N165, 
	clk_m__L3_N166, 
	clk_m__L3_N167, 
	clk_m__L3_N168, 
	clk_m__L3_N169, 
	clk_m__L3_N17, 
	clk_m__L3_N170, 
	clk_m__L3_N171, 
	clk_m__L3_N172, 
	clk_m__L3_N173, 
	clk_m__L3_N174, 
	clk_m__L3_N175, 
	clk_m__L3_N176, 
	clk_m__L3_N177, 
	clk_m__L3_N18, 
	clk_m__L3_N19, 
	clk_m__L3_N2, 
	clk_m__L3_N20, 
	clk_m__L3_N21, 
	clk_m__L3_N22, 
	clk_m__L3_N23, 
	clk_m__L3_N24, 
	clk_m__L3_N25, 
	clk_m__L3_N26, 
	clk_m__L3_N27, 
	clk_m__L3_N28, 
	clk_m__L3_N29, 
	clk_m__L3_N3, 
	clk_m__L3_N30, 
	clk_m__L3_N31, 
	clk_m__L3_N32, 
	clk_m__L3_N33, 
	clk_m__L3_N34, 
	clk_m__L3_N35, 
	clk_m__L3_N36, 
	clk_m__L3_N37, 
	clk_m__L3_N38, 
	clk_m__L3_N39, 
	clk_m__L3_N4, 
	clk_m__L3_N40, 
	clk_m__L3_N41, 
	clk_m__L3_N42, 
	clk_m__L3_N43, 
	clk_m__L3_N44, 
	clk_m__L3_N45, 
	clk_m__L3_N46, 
	clk_m__L3_N47, 
	clk_m__L3_N48, 
	clk_m__L3_N49, 
	clk_m__L3_N5, 
	clk_m__L3_N50, 
	clk_m__L3_N52, 
	clk_m__L3_N53, 
	clk_m__L3_N54, 
	clk_m__L3_N55, 
	clk_m__L3_N56, 
	clk_m__L3_N57, 
	clk_m__L3_N58, 
	clk_m__L3_N59, 
	clk_m__L3_N6, 
	clk_m__L3_N60, 
	clk_m__L3_N61, 
	clk_m__L3_N62, 
	clk_m__L3_N63, 
	clk_m__L3_N64, 
	clk_m__L3_N65, 
	clk_m__L3_N66, 
	clk_m__L3_N67, 
	clk_m__L3_N68, 
	clk_m__L3_N69, 
	clk_m__L3_N7, 
	clk_m__L3_N70, 
	clk_m__L3_N71, 
	clk_m__L3_N72, 
	clk_m__L3_N73, 
	clk_m__L3_N74, 
	clk_m__L3_N75, 
	clk_m__L3_N76, 
	clk_m__L3_N77, 
	clk_m__L3_N78, 
	clk_m__L3_N79, 
	clk_m__L3_N8, 
	clk_m__L3_N80, 
	clk_m__L3_N81, 
	clk_m__L3_N82, 
	clk_m__L3_N83, 
	clk_m__L3_N84, 
	clk_m__L3_N85, 
	clk_m__L3_N86, 
	clk_m__L3_N87, 
	clk_m__L3_N88, 
	clk_m__L3_N89, 
	clk_m__L3_N9, 
	clk_m__L3_N90, 
	clk_m__L3_N91, 
	clk_m__L3_N92, 
	clk_m__L3_N93, 
	clk_m__L3_N94, 
	clk_m__L3_N95, 
	clk_m__L3_N96, 
	clk_m__L3_N97, 
	clk_m__L3_N98, 
	clk_m__L3_N99, 
	clk_m__N0);
   input clk;
   input [15:0] mem_access_addr;
   input [15:0] mem_write_data;
   input mem_write_en;
   input mem_read;
   output [15:0] mem_read_data;
   input clk_m__L3_N1;
   input clk_m__L3_N10;
   input clk_m__L3_N100;
   input clk_m__L3_N101;
   input clk_m__L3_N102;
   input clk_m__L3_N103;
   input clk_m__L3_N104;
   input clk_m__L3_N105;
   input clk_m__L3_N106;
   input clk_m__L3_N107;
   input clk_m__L3_N108;
   input clk_m__L3_N109;
   input clk_m__L3_N11;
   input clk_m__L3_N110;
   input clk_m__L3_N111;
   input clk_m__L3_N112;
   input clk_m__L3_N113;
   input clk_m__L3_N114;
   input clk_m__L3_N115;
   input clk_m__L3_N116;
   input clk_m__L3_N117;
   input clk_m__L3_N118;
   input clk_m__L3_N119;
   input clk_m__L3_N12;
   input clk_m__L3_N120;
   input clk_m__L3_N121;
   input clk_m__L3_N122;
   input clk_m__L3_N123;
   input clk_m__L3_N124;
   input clk_m__L3_N125;
   input clk_m__L3_N126;
   input clk_m__L3_N127;
   input clk_m__L3_N128;
   input clk_m__L3_N129;
   input clk_m__L3_N13;
   input clk_m__L3_N130;
   input clk_m__L3_N131;
   input clk_m__L3_N132;
   input clk_m__L3_N133;
   input clk_m__L3_N134;
   input clk_m__L3_N135;
   input clk_m__L3_N136;
   input clk_m__L3_N137;
   input clk_m__L3_N138;
   input clk_m__L3_N139;
   input clk_m__L3_N14;
   input clk_m__L3_N140;
   input clk_m__L3_N141;
   input clk_m__L3_N142;
   input clk_m__L3_N143;
   input clk_m__L3_N144;
   input clk_m__L3_N145;
   input clk_m__L3_N146;
   input clk_m__L3_N147;
   input clk_m__L3_N148;
   input clk_m__L3_N149;
   input clk_m__L3_N15;
   input clk_m__L3_N150;
   input clk_m__L3_N151;
   input clk_m__L3_N152;
   input clk_m__L3_N153;
   input clk_m__L3_N154;
   input clk_m__L3_N155;
   input clk_m__L3_N156;
   input clk_m__L3_N157;
   input clk_m__L3_N158;
   input clk_m__L3_N159;
   input clk_m__L3_N16;
   input clk_m__L3_N160;
   input clk_m__L3_N161;
   input clk_m__L3_N162;
   input clk_m__L3_N163;
   input clk_m__L3_N164;
   input clk_m__L3_N165;
   input clk_m__L3_N166;
   input clk_m__L3_N167;
   input clk_m__L3_N168;
   input clk_m__L3_N169;
   input clk_m__L3_N17;
   input clk_m__L3_N170;
   input clk_m__L3_N171;
   input clk_m__L3_N172;
   input clk_m__L3_N173;
   input clk_m__L3_N174;
   input clk_m__L3_N175;
   input clk_m__L3_N176;
   input clk_m__L3_N177;
   input clk_m__L3_N18;
   input clk_m__L3_N19;
   input clk_m__L3_N2;
   input clk_m__L3_N20;
   input clk_m__L3_N21;
   input clk_m__L3_N22;
   input clk_m__L3_N23;
   input clk_m__L3_N24;
   input clk_m__L3_N25;
   input clk_m__L3_N26;
   input clk_m__L3_N27;
   input clk_m__L3_N28;
   input clk_m__L3_N29;
   input clk_m__L3_N3;
   input clk_m__L3_N30;
   input clk_m__L3_N31;
   input clk_m__L3_N32;
   input clk_m__L3_N33;
   input clk_m__L3_N34;
   input clk_m__L3_N35;
   input clk_m__L3_N36;
   input clk_m__L3_N37;
   input clk_m__L3_N38;
   input clk_m__L3_N39;
   input clk_m__L3_N4;
   input clk_m__L3_N40;
   input clk_m__L3_N41;
   input clk_m__L3_N42;
   input clk_m__L3_N43;
   input clk_m__L3_N44;
   input clk_m__L3_N45;
   input clk_m__L3_N46;
   input clk_m__L3_N47;
   input clk_m__L3_N48;
   input clk_m__L3_N49;
   input clk_m__L3_N5;
   input clk_m__L3_N50;
   input clk_m__L3_N52;
   input clk_m__L3_N53;
   input clk_m__L3_N54;
   input clk_m__L3_N55;
   input clk_m__L3_N56;
   input clk_m__L3_N57;
   input clk_m__L3_N58;
   input clk_m__L3_N59;
   input clk_m__L3_N6;
   input clk_m__L3_N60;
   input clk_m__L3_N61;
   input clk_m__L3_N62;
   input clk_m__L3_N63;
   input clk_m__L3_N64;
   input clk_m__L3_N65;
   input clk_m__L3_N66;
   input clk_m__L3_N67;
   input clk_m__L3_N68;
   input clk_m__L3_N69;
   input clk_m__L3_N7;
   input clk_m__L3_N70;
   input clk_m__L3_N71;
   input clk_m__L3_N72;
   input clk_m__L3_N73;
   input clk_m__L3_N74;
   input clk_m__L3_N75;
   input clk_m__L3_N76;
   input clk_m__L3_N77;
   input clk_m__L3_N78;
   input clk_m__L3_N79;
   input clk_m__L3_N8;
   input clk_m__L3_N80;
   input clk_m__L3_N81;
   input clk_m__L3_N82;
   input clk_m__L3_N83;
   input clk_m__L3_N84;
   input clk_m__L3_N85;
   input clk_m__L3_N86;
   input clk_m__L3_N87;
   input clk_m__L3_N88;
   input clk_m__L3_N89;
   input clk_m__L3_N9;
   input clk_m__L3_N90;
   input clk_m__L3_N91;
   input clk_m__L3_N92;
   input clk_m__L3_N93;
   input clk_m__L3_N94;
   input clk_m__L3_N95;
   input clk_m__L3_N96;
   input clk_m__L3_N97;
   input clk_m__L3_N98;
   input clk_m__L3_N99;
   input clk_m__N0;

   // Internal wires
   wire FE_PHN7506_n2582;
   wire FE_PHN7505_n2417;
   wire FE_PHN7504_n2582;
   wire FE_PHN7503_n1001;
   wire FE_PHN7502_n1014;
   wire FE_PHN7501_n2890;
   wire FE_PHN7500_n2180;
   wire FE_PHN7499_n4102;
   wire FE_PHN7498_n2395;
   wire FE_PHN7497_n2417;
   wire FE_PHN7496_n2582;
   wire FE_PHN7495_n1013;
   wire FE_PHN7494_n1001;
   wire FE_PHN7493_n3964;
   wire FE_PHN7492_n1017;
   wire FE_PHN7491_n974;
   wire FE_PHN7490_n1014;
   wire FE_PHN7489_n2394;
   wire FE_PHN7488_n3953;
   wire FE_PHN7487_n3934;
   wire FE_PHN7486_n2132;
   wire FE_PHN7485_n2168;
   wire FE_PHN7484_n3960;
   wire FE_PHN7483_n2571;
   wire FE_PHN7482_n3923;
   wire FE_PHN7481_n2892;
   wire FE_PHN7480_n2155;
   wire FE_PHN7479_n2175;
   wire FE_PHN7478_n3968;
   wire FE_PHN7477_n2628;
   wire FE_PHN7476_n2159;
   wire FE_PHN7475_n2592;
   wire FE_PHN7474_n4155;
   wire FE_PHN7473_n2170;
   wire FE_PHN7472_n4137;
   wire FE_PHN7471_n4147;
   wire FE_PHN7470_n2166;
   wire FE_PHN7469_n3230;
   wire FE_PHN7468_n2614;
   wire FE_PHN7467_n2395;
   wire FE_PHN7466_n2130;
   wire FE_PHN7465_n2890;
   wire FE_PHN7464_n4102;
   wire FE_PHN7463_n2180;
   wire FE_PHN7462_n2417;
   wire FE_PHN7461_n2582;
   wire FE_PHN7460_n979;
   wire FE_PHN7459_n1154;
   wire FE_PHN7458_n938;
   wire FE_PHN7457_n1001;
   wire FE_PHN7456_n4215;
   wire FE_PHN7455_n3129;
   wire FE_PHN7454_n4229;
   wire FE_PHN7453_n3964;
   wire FE_PHN7452_n3028;
   wire FE_PHN7451_n974;
   wire FE_PHN7450_n1017;
   wire FE_PHN7449_n1014;
   wire FE_PHN7448_n2426;
   wire FE_PHN7447_n4013;
   wire FE_PHN7446_n2119;
   wire FE_PHN7445_n2393;
   wire FE_PHN7444_n2133;
   wire FE_PHN7443_n2604;
   wire FE_PHN7442_n3068;
   wire FE_PHN7441_n2164;
   wire FE_PHN7440_n2126;
   wire FE_PHN7439_n2378;
   wire FE_PHN7438_n2151;
   wire FE_PHN7437_n2610;
   wire FE_PHN7436_n2165;
   wire FE_PHN7435_n2379;
   wire FE_PHN7434_n2118;
   wire FE_PHN7433_n2167;
   wire FE_PHN7432_n2603;
   wire FE_PHN7431_n2135;
   wire FE_PHN7430_n2887;
   wire FE_PHN7429_n2169;
   wire FE_PHN7428_n3953;
   wire FE_PHN7427_n2179;
   wire FE_PHN7426_n3934;
   wire FE_PHN7425_n2154;
   wire FE_PHN7424_n2168;
   wire FE_PHN7423_n2892;
   wire FE_PHN7422_n2570;
   wire FE_PHN7421_n2434;
   wire FE_PHN7420_n3968;
   wire FE_PHN7419_n4155;
   wire FE_PHN7418_n2410;
   wire FE_PHN7417_n2152;
   wire FE_PHN7416_n2132;
   wire FE_PHN7415_n2175;
   wire FE_PHN7414_n2394;
   wire FE_PHN7413_n2170;
   wire FE_PHN7412_n2120;
   wire FE_PHN7411_n2628;
   wire FE_PHN7410_n4121;
   wire FE_PHN7409_n4137;
   wire FE_PHN7408_n2402;
   wire FE_PHN7407_n2571;
   wire FE_PHN7406_n3960;
   wire FE_PHN7405_n2155;
   wire FE_PHN7404_n3923;
   wire FE_PHN7403_n2625;
   wire FE_PHN7402_n2578;
   wire FE_PHN7401_n1863;
   wire FE_PHN7400_n2159;
   wire FE_PHN7399_n4139;
   wire FE_PHN7398_n2166;
   wire FE_PHN7397_n2395;
   wire FE_PHN7396_n2592;
   wire FE_PHN7395_n3230;
   wire FE_PHN7394_n4163;
   wire FE_PHN7393_n2614;
   wire FE_PHN7392_n4147;
   wire FE_PHN7391_n2130;
   wire FE_PHN7390_n2890;
   wire FE_PHN7389_n4102;
   wire FE_PHN7388_n2180;
   wire FE_PHN7387_n2417;
   wire FE_PHN7386_n2582;
   wire FE_PHN7385_n914;
   wire FE_PHN7384_n2857;
   wire FE_PHN7383_n901;
   wire FE_PHN7382_n1007;
   wire FE_PHN7381_n2594;
   wire FE_PHN7380_n996;
   wire FE_PHN7379_n2380;
   wire FE_PHN7378_n2398;
   wire FE_PHN7377_n4027;
   wire FE_PHN7376_n4210;
   wire FE_PHN7375_n1054;
   wire FE_PHN7374_n2696;
   wire FE_PHN7373_n2172;
   wire FE_PHN7372_n3965;
   wire FE_PHN7371_n3212;
   wire FE_PHN7370_n1922;
   wire FE_PHN7369_n4308;
   wire FE_PHN7368_n4274;
   wire FE_PHN7367_n1880;
   wire FE_PHN7366_n985;
   wire FE_PHN7365_n2587;
   wire FE_PHN7364_n2619;
   wire FE_PHN7363_n2181;
   wire FE_PHN7362_n933;
   wire FE_PHN7361_n2163;
   wire FE_PHN7360_n4142;
   wire FE_PHN7359_n1918;
   wire FE_PHN7358_n2876;
   wire FE_PHN7357_n1094;
   wire FE_PHN7356_n1031;
   wire FE_PHN7355_n3955;
   wire FE_PHN7354_n3971;
   wire FE_PHN7353_n2566;
   wire FE_PHN7352_n3932;
   wire FE_PHN7351_n4110;
   wire FE_PHN7350_n4018;
   wire FE_PHN7349_n2428;
   wire FE_PHN7348_n2388;
   wire FE_PHN7347_n4273;
   wire FE_PHN7346_n3970;
   wire FE_PHN7345_n1874;
   wire FE_PHN7344_n2747;
   wire FE_PHN7343_n2618;
   wire FE_PHN7342_n2432;
   wire FE_PHN7341_n2695;
   wire FE_PHN7340_n4116;
   wire FE_PHN7339_n2121;
   wire FE_PHN7338_n2149;
   wire FE_PHN7337_n1015;
   wire FE_PHN7336_n4294;
   wire FE_PHN7335_n2611;
   wire FE_PHN7334_n953;
   wire FE_PHN7333_n1190;
   wire FE_PHN7332_n2412;
   wire FE_PHN7331_n2750;
   wire FE_PHN7330_n1919;
   wire FE_PHN7329_n1872;
   wire FE_PHN7328_n1906;
   wire FE_PHN7327_n2602;
   wire FE_PHN7326_n950;
   wire FE_PHN7325_n2576;
   wire FE_PHN7324_n1178;
   wire FE_PHN7323_n2124;
   wire FE_PHN7322_n4148;
   wire FE_PHN7321_n906;
   wire FE_PHN7320_n964;
   wire FE_PHN7319_n979;
   wire FE_PHN7318_n2622;
   wire FE_PHN7317_n2572;
   wire FE_PHN7316_n2138;
   wire FE_PHN7315_n2612;
   wire FE_PHN7314_n4114;
   wire FE_PHN7313_n1154;
   wire FE_PHN7312_n2251;
   wire FE_PHN7311_n938;
   wire FE_PHN7310_n1001;
   wire FE_PHN7309_n4046;
   wire FE_PHN7308_n3072;
   wire FE_PHN7307_n3052;
   wire FE_PHN7306_n2564;
   wire FE_PHN7305_n4180;
   wire FE_PHN7304_n928;
   wire FE_PHN7303_n905;
   wire FE_PHN7302_n3919;
   wire FE_PHN7301_n4215;
   wire FE_PHN7300_n4219;
   wire FE_PHN7299_n2574;
   wire FE_PHN7298_n4174;
   wire FE_PHN7297_n975;
   wire FE_PHN7296_n2599;
   wire FE_PHN7295_n1082;
   wire FE_PHN7294_n948;
   wire FE_PHN7293_n3129;
   wire FE_PHN7292_n2580;
   wire FE_PHN7291_n3028;
   wire FE_PHN7290_n1017;
   wire FE_PHN7289_n4229;
   wire FE_PHN7288_n1014;
   wire FE_PHN7287_n3964;
   wire FE_PHN7286_n974;
   wire FE_PHN7285_n1013;
   wire FE_PHN7284_n4365;
   wire FE_PHN7283_n2972;
   wire FE_PHN7282_n4409;
   wire FE_PHN7281_n3068;
   wire FE_PHN7280_n2887;
   wire FE_PHN7279_n2426;
   wire FE_PHN7278_n4013;
   wire FE_PHN7277_n2133;
   wire FE_PHN7276_n2892;
   wire FE_PHN7275_n2425;
   wire FE_PHN7274_n2379;
   wire FE_PHN7273_n2377;
   wire FE_PHN7272_n4011;
   wire FE_PHN7271_n2119;
   wire FE_PHN7270_n2151;
   wire FE_PHN7269_n2427;
   wire FE_PHN7268_n2126;
   wire FE_PHN7267_n2395;
   wire FE_PHN7266_n4002;
   wire FE_PHN7265_n2603;
   wire FE_PHN7264_n2434;
   wire FE_PHN7263_n2610;
   wire FE_PHN7262_n3953;
   wire FE_PHN7261_n2570;
   wire FE_PHN7260_n2135;
   wire FE_PHN7259_n2179;
   wire FE_PHN7258_n2378;
   wire FE_PHN7257_n2165;
   wire FE_PHN7256_n2168;
   wire FE_PHN7255_n2175;
   wire FE_PHN7254_n2118;
   wire FE_PHN7253_n2393;
   wire FE_PHN7252_n2169;
   wire FE_PHN7251_n2152;
   wire FE_PHN7250_n2164;
   wire FE_PHN7249_n2890;
   wire FE_PHN7248_n2120;
   wire FE_PHN7247_n3934;
   wire FE_PHN7246_n2571;
   wire FE_PHN7245_n4153;
   wire FE_PHN7244_n2410;
   wire FE_PHN7243_n3960;
   wire FE_PHN7242_n4137;
   wire FE_PHN7241_n2578;
   wire FE_PHN7240_n3923;
   wire FE_PHN7239_n2132;
   wire FE_PHN7238_n3230;
   wire FE_PHN7237_n3968;
   wire FE_PHN7236_n2417;
   wire FE_PHN7235_n4155;
   wire FE_PHN7234_n2167;
   wire FE_PHN7233_n4121;
   wire FE_PHN7232_n2155;
   wire FE_PHN7231_n2154;
   wire FE_PHN7230_n2180;
   wire FE_PHN7229_n2394;
   wire FE_PHN7228_n2402;
   wire FE_PHN7227_n2625;
   wire FE_PHN7226_n2159;
   wire FE_PHN7225_n2170;
   wire FE_PHN7224_n2582;
   wire FE_PHN7223_n4139;
   wire FE_PHN7222_n4147;
   wire FE_PHN7221_n2166;
   wire FE_PHN7220_n2592;
   wire FE_PHN7219_n2628;
   wire FE_PHN7218_n1863;
   wire FE_PHN7217_n2614;
   wire FE_PHN7216_n4102;
   wire FE_PHN7215_n4163;
   wire FE_PHN7214_n2130;
   wire FE_PHN7213_n2604;
   wire FE_PHN7212_n3150;
   wire FE_PHN7211_n4135;
   wire FE_PHN7210_n880;
   wire FE_PHN7209_n1913;
   wire FE_PHN7208_n2422;
   wire FE_PHN7207_n4107;
   wire FE_PHN7206_n3017;
   wire FE_PHN7205_n1086;
   wire FE_PHN7204_n4016;
   wire FE_PHN7203_n2697;
   wire FE_PHN7202_n3944;
   wire FE_PHN7201_n3962;
   wire FE_PHN7200_n921;
   wire FE_PHN7199_n2609;
   wire FE_PHN7198_n2123;
   wire FE_PHN7197_n2177;
   wire FE_PHN7196_n2589;
   wire FE_PHN7195_n2743;
   wire FE_PHN7194_n2873;
   wire FE_PHN7193_n1028;
   wire FE_PHN7192_n973;
   wire FE_PHN7191_n2749;
   wire FE_PHN7190_n3047;
   wire FE_PHN7189_n3021;
   wire FE_PHN7188_n2171;
   wire FE_PHN7187_n1908;
   wire FE_PHN7186_n2590;
   wire FE_PHN7185_n2381;
   wire FE_PHN7184_n2122;
   wire FE_PHN7183_n2935;
   wire FE_PHN7182_n4151;
   wire FE_PHN7181_n1375;
   wire FE_PHN7180_n2616;
   wire FE_PHN7179_n1012;
   wire FE_PHN7178_n967;
   wire FE_PHN7177_n981;
   wire FE_PHN7176_n2624;
   wire FE_PHN7175_n2919;
   wire FE_PHN7174_n4008;
   wire FE_PHN7173_n4158;
   wire FE_PHN7172_n2176;
   wire FE_PHN7171_n2904;
   wire FE_PHN7170_n2701;
   wire FE_PHN7169_n4404;
   wire FE_PHN7168_n4331;
   wire FE_PHN7167_n1865;
   wire FE_PHN7166_n2908;
   wire FE_PHN7165_n3033;
   wire FE_PHN7164_n2889;
   wire FE_PHN7163_n4259;
   wire FE_PHN7162_n3965;
   wire FE_PHN7161_n4358;
   wire FE_PHN7160_n1158;
   wire FE_PHN7159_n4035;
   wire FE_PHN7158_n4150;
   wire FE_PHN7157_n4062;
   wire FE_PHN7156_n2386;
   wire FE_PHN7155_n3945;
   wire FE_PHN7154_n2922;
   wire FE_PHN7153_n3212;
   wire FE_PHN7152_n2390;
   wire FE_PHN7151_n1007;
   wire FE_PHN7150_n2893;
   wire FE_PHN7149_n1286;
   wire FE_PHN7148_n2907;
   wire FE_PHN7147_n1019;
   wire FE_PHN7146_n2626;
   wire FE_PHN7145_n1003;
   wire FE_PHN7144_n888;
   wire FE_PHN7143_n4308;
   wire FE_PHN7142_n2161;
   wire FE_PHN7141_n4034;
   wire FE_PHN7140_n2925;
   wire FE_PHN7139_n2144;
   wire FE_PHN7138_n2432;
   wire FE_PHN7137_n3979;
   wire FE_PHN7136_n4210;
   wire FE_PHN7135_n4032;
   wire FE_PHN7134_n2938;
   wire FE_PHN7133_n4012;
   wire FE_PHN7132_n2403;
   wire FE_PHN7131_n2941;
   wire FE_PHN7130_n901;
   wire FE_PHN7129_n985;
   wire FE_PHN7128_n2375;
   wire FE_PHN7127_n983;
   wire FE_PHN7126_n996;
   wire FE_PHN7125_n2125;
   wire FE_PHN7124_n4242;
   wire FE_PHN7123_n2696;
   wire FE_PHN7122_n4274;
   wire FE_PHN7121_n2857;
   wire FE_PHN7120_n3983;
   wire FE_PHN7119_n2587;
   wire FE_PHN7118_n917;
   wire FE_PHN7117_n3260;
   wire FE_PHN7116_n2257;
   wire FE_PHN7115_n3980;
   wire FE_PHN7114_n1906;
   wire FE_PHN7113_n4031;
   wire FE_PHN7112_n2398;
   wire FE_PHN7111_n2876;
   wire FE_PHN7110_n962;
   wire FE_PHN7109_n930;
   wire FE_PHN7108_n933;
   wire FE_PHN7107_n914;
   wire FE_PHN7106_n2577;
   wire FE_PHN7105_n2424;
   wire FE_PHN7104_n949;
   wire FE_PHN7103_n2407;
   wire FE_PHN7102_n2148;
   wire FE_PHN7101_n2695;
   wire FE_PHN7100_n1054;
   wire FE_PHN7099_n2566;
   wire FE_PHN7098_n4273;
   wire FE_PHN7097_n1031;
   wire FE_PHN7096_n2419;
   wire FE_PHN7095_n2181;
   wire FE_PHN7094_n980;
   wire FE_PHN7093_n2615;
   wire FE_PHN7092_n3981;
   wire FE_PHN7091_n2747;
   wire FE_PHN7090_n4027;
   wire FE_PHN7089_n3971;
   wire FE_PHN7088_n2163;
   wire FE_PHN7087_n3966;
   wire FE_PHN7086_n2750;
   wire FE_PHN7085_n4294;
   wire FE_PHN7084_n2406;
   wire FE_PHN7083_n2429;
   wire FE_PHN7082_n2382;
   wire FE_PHN7081_n2172;
   wire FE_PHN7080_n3970;
   wire FE_PHN7079_n2121;
   wire FE_PHN7078_n2131;
   wire FE_PHN7077_n3955;
   wire FE_PHN7076_n2619;
   wire FE_PHN7075_n4018;
   wire FE_PHN7074_n979;
   wire FE_PHN7073_n2401;
   wire FE_PHN7072_n2156;
   wire FE_PHN7071_n1015;
   wire FE_PHN7070_n2376;
   wire FE_PHN7069_n1190;
   wire FE_PHN7068_n2380;
   wire FE_PHN7067_n927;
   wire FE_PHN7066_n2428;
   wire FE_PHN7065_n944;
   wire FE_PHN7064_n1094;
   wire FE_PHN7063_n1874;
   wire FE_PHN7062_n2611;
   wire FE_PHN7061_n1178;
   wire FE_PHN7060_n1872;
   wire FE_PHN7059_n4116;
   wire FE_PHN7058_n2411;
   wire FE_PHN7057_n4148;
   wire FE_PHN7056_n1918;
   wire FE_PHN7055_n964;
   wire FE_PHN7054_n2423;
   wire FE_PHN7053_n3932;
   wire FE_PHN7052_n950;
   wire FE_PHN7051_n2594;
   wire FE_PHN7050_n906;
   wire FE_PHN7049_n2137;
   wire FE_PHN7048_n2138;
   wire FE_PHN7047_n2149;
   wire FE_PHN7046_n2618;
   wire FE_PHN7045_n2124;
   wire FE_PHN7044_n4142;
   wire FE_PHN7043_n1880;
   wire FE_PHN7042_n1154;
   wire FE_PHN7041_n2622;
   wire FE_PHN7040_n953;
   wire FE_PHN7039_n2598;
   wire FE_PHN7038_n1922;
   wire FE_PHN7037_n2602;
   wire FE_PHN7036_n1919;
   wire FE_PHN7035_n2576;
   wire FE_PHN7034_n938;
   wire FE_PHN7033_n4110;
   wire FE_PHN7032_n2388;
   wire FE_PHN7031_n1001;
   wire FE_PHN7030_n2412;
   wire FE_PHN7029_n4114;
   wire FE_PHN7028_n2572;
   wire FE_PHN7027_n2251;
   wire FE_PHN7026_n2612;
   wire FE_PHN7025_n844;
   wire FE_PHN7024_n3131;
   wire FE_PHN7023_n3924;
   wire FE_PHN7022_n4204;
   wire FE_PHN7021_n2995;
   wire FE_PHN7020_n1021;
   wire FE_PHN7019_n3112;
   wire FE_PHN7018_ram_229__12_;
   wire FE_PHN7017_n882;
   wire FE_PHN7016_n2928;
   wire FE_PHN7015_n1030;
   wire FE_PHN7014_n3078;
   wire FE_PHN7013_n2970;
   wire FE_PHN7012_n4243;
   wire FE_PHN7011_n2980;
   wire FE_PHN7010_n3087;
   wire FE_PHN7009_n2896;
   wire FE_PHN7008_n4245;
   wire FE_PHN7007_n4238;
   wire FE_PHN7006_n870;
   wire FE_PHN7005_ram_145__7_;
   wire FE_PHN7004_n4359;
   wire FE_PHN7003_n4094;
   wire FE_PHN7002_n4196;
   wire FE_PHN7001_n4262;
   wire FE_PHN7000_n3921;
   wire FE_PHN6999_n999;
   wire FE_PHN6998_n2906;
   wire FE_PHN6997_n891;
   wire FE_PHN6996_n4281;
   wire FE_PHN6995_n3075;
   wire FE_PHN6994_n4251;
   wire FE_PHN6993_n3926;
   wire FE_PHN6992_n3056;
   wire FE_PHN6991_n4134;
   wire FE_PHN6990_n3099;
   wire FE_PHN6989_n2997;
   wire FE_PHN6988_n969;
   wire FE_PHN6987_n3918;
   wire FE_PHN6986_n1068;
   wire FE_PHN6985_n3969;
   wire FE_PHN6984_n3265;
   wire FE_PHN6983_n3940;
   wire FE_PHN6982_n884;
   wire FE_PHN6981_n4201;
   wire FE_PHN6980_n951;
   wire FE_PHN6979_n890;
   wire FE_PHN6978_n4333;
   wire FE_PHN6977_n3108;
   wire FE_PHN6976_ram_214__13_;
   wire FE_PHN6975_n4266;
   wire FE_PHN6974_n1006;
   wire FE_PHN6973_n2926;
   wire FE_PHN6972_n4269;
   wire FE_PHN6971_n2994;
   wire FE_PHN6970_n3098;
   wire FE_PHN6969_n2897;
   wire FE_PHN6968_n3024;
   wire FE_PHN6967_n2933;
   wire FE_PHN6966_n3076;
   wire FE_PHN6965_n3084;
   wire FE_PHN6964_n3958;
   wire FE_PHN6963_n4271;
   wire FE_PHN6962_n4339;
   wire FE_PHN6961_n3994;
   wire FE_PHN6960_n1110;
   wire FE_PHN6959_n2934;
   wire FE_PHN6958_n892;
   wire FE_PHN6957_n4355;
   wire FE_PHN6956_n4003;
   wire FE_PHN6955_n2978;
   wire FE_PHN6954_n2946;
   wire FE_PHN6953_n4362;
   wire FE_PHN6952_n3103;
   wire FE_PHN6951_n3931;
   wire FE_PHN6950_n4410;
   wire FE_PHN6949_n4361;
   wire FE_PHN6948_n2987;
   wire FE_PHN6947_n4233;
   wire FE_PHN6946_n4387;
   wire FE_PHN6945_ram_153__11_;
   wire FE_PHN6944_n2399;
   wire FE_PHN6943_n3079;
   wire FE_PHN6942_n919;
   wire FE_PHN6941_n1020;
   wire FE_PHN6940_n2413;
   wire FE_PHN6939_n957;
   wire FE_PHN6938_n2992;
   wire FE_PHN6937_n3952;
   wire FE_PHN6936_n3910;
   wire FE_PHN6935_n1093;
   wire FE_PHN6934_n4076;
   wire FE_PHN6933_ram_221__1_;
   wire FE_PHN6932_n4222;
   wire FE_PHN6931_n2916;
   wire FE_PHN6930_n3915;
   wire FE_PHN6929_n4295;
   wire FE_PHN6928_n1087;
   wire FE_PHN6927_n4169;
   wire FE_PHN6926_n4291;
   wire FE_PHN6925_n4202;
   wire FE_PHN6924_n3956;
   wire FE_PHN6923_n3060;
   wire FE_PHN6922_n3976;
   wire FE_PHN6921_n3996;
   wire FE_PHN6920_n3947;
   wire FE_PHN6919_n848;
   wire FE_PHN6918_n4183;
   wire FE_PHN6917_n2621;
   wire FE_PHN6916_n4111;
   wire FE_PHN6915_n4021;
   wire FE_PHN6914_n936;
   wire FE_PHN6913_ram_144__8_;
   wire FE_PHN6912_n3954;
   wire FE_PHN6911_n846;
   wire FE_PHN6910_n994;
   wire FE_PHN6909_n2936;
   wire FE_PHN6908_n4371;
   wire FE_PHN6907_n3936;
   wire FE_PHN6906_n2735;
   wire FE_PHN6905_n1899;
   wire FE_PHN6904_n4311;
   wire FE_PHN6903_n3984;
   wire FE_PHN6902_n876;
   wire FE_PHN6901_n2437;
   wire FE_PHN6900_n4239;
   wire FE_PHN6899_n872;
   wire FE_PHN6898_n3951;
   wire FE_PHN6897_n3959;
   wire FE_PHN6896_n3998;
   wire FE_PHN6895_n840;
   wire FE_PHN6894_n4252;
   wire FE_PHN6893_n988;
   wire FE_PHN6892_n961;
   wire FE_PHN6891_n4172;
   wire FE_PHN6890_n1106;
   wire FE_PHN6889_n3948;
   wire FE_PHN6888_n2158;
   wire FE_PHN6887_n3027;
   wire FE_PHN6886_n4033;
   wire FE_PHN6885_n958;
   wire FE_PHN6884_n2967;
   wire FE_PHN6883_n4324;
   wire FE_PHN6882_n4017;
   wire FE_PHN6881_n2374;
   wire FE_PHN6880_n4028;
   wire FE_PHN6879_n3972;
   wire FE_PHN6878_n3914;
   wire FE_PHN6877_n1056;
   wire FE_PHN6876_n3063;
   wire FE_PHN6875_n3025;
   wire FE_PHN6874_n4005;
   wire FE_PHN6873_n1066;
   wire FE_PHN6872_n3257;
   wire FE_PHN6871_n4185;
   wire FE_PHN6870_n4166;
   wire FE_PHN6869_n4188;
   wire FE_PHN6868_n839;
   wire FE_PHN6867_n4327;
   wire FE_PHN6866_n851;
   wire FE_PHN6865_n3937;
   wire FE_PHN6864_n989;
   wire FE_PHN6863_n1078;
   wire FE_PHN6862_ram_133__9_;
   wire FE_PHN6861_n3987;
   wire FE_PHN6860_n2943;
   wire FE_PHN6859_n2998;
   wire FE_PHN6858_n902;
   wire FE_PHN6857_n4211;
   wire FE_PHN6856_n4377;
   wire FE_PHN6855_n3943;
   wire FE_PHN6854_n4226;
   wire FE_PHN6853_n855;
   wire FE_PHN6852_n1051;
   wire FE_PHN6851_n3029;
   wire FE_PHN6850_n3930;
   wire FE_PHN6849_n2971;
   wire FE_PHN6848_n852;
   wire FE_PHN6847_n3116;
   wire FE_PHN6846_n857;
   wire FE_PHN6845_n3963;
   wire FE_PHN6844_n1069;
   wire FE_PHN6843_n2258;
   wire FE_PHN6842_n4217;
   wire FE_PHN6841_n3043;
   wire FE_PHN6840_n4323;
   wire FE_PHN6839_n2396;
   wire FE_PHN6838_n2930;
   wire FE_PHN6837_n3207;
   wire FE_PHN6836_n2433;
   wire FE_PHN6835_n3052;
   wire FE_PHN6834_n887;
   wire FE_PHN6833_n945;
   wire FE_PHN6832_n1896;
   wire FE_PHN6831_n965;
   wire FE_PHN6830_n2722;
   wire FE_PHN6829_n941;
   wire FE_PHN6828_n2127;
   wire FE_PHN6827_n1034;
   wire FE_PHN6826_n2623;
   wire FE_PHN6825_n858;
   wire FE_PHN6824_n4220;
   wire FE_PHN6823_n3927;
   wire FE_PHN6822_n866;
   wire FE_PHN6821_n889;
   wire FE_PHN6820_n4393;
   wire FE_PHN6819_n4278;
   wire FE_PHN6818_n4036;
   wire FE_PHN6817_n1037;
   wire FE_PHN6816_n2932;
   wire FE_PHN6815_n920;
   wire FE_PHN6814_n4307;
   wire FE_PHN6813_n4029;
   wire FE_PHN6812_n864;
   wire FE_PHN6811_n2754;
   wire FE_PHN6810_n3988;
   wire FE_PHN6809_n3023;
   wire FE_PHN6808_n4195;
   wire FE_PHN6807_n972;
   wire FE_PHN6806_n878;
   wire FE_PHN6805_n856;
   wire FE_PHN6804_n2430;
   wire FE_PHN6803_n4299;
   wire FE_PHN6802_n3073;
   wire FE_PHN6801_n894;
   wire FE_PHN6800_n2141;
   wire FE_PHN6799_n3916;
   wire FE_PHN6798_n4014;
   wire FE_PHN6797_n913;
   wire FE_PHN6796_n3055;
   wire FE_PHN6795_n861;
   wire FE_PHN6794_n943;
   wire FE_PHN6793_n4340;
   wire FE_PHN6792_n3071;
   wire FE_PHN6791_n929;
   wire FE_PHN6790_n2900;
   wire FE_PHN6789_n1079;
   wire FE_PHN6788_n4232;
   wire FE_PHN6787_n4209;
   wire FE_PHN6786_n1022;
   wire FE_PHN6785_n2178;
   wire FE_PHN6784_n4225;
   wire FE_PHN6783_n935;
   wire FE_PHN6782_n4001;
   wire FE_PHN6781_n4277;
   wire FE_PHN6780_n842;
   wire FE_PHN6779_n2927;
   wire FE_PHN6778_n925;
   wire FE_PHN6777_n2400;
   wire FE_PHN6776_n910;
   wire FE_PHN6775_n4240;
   wire FE_PHN6774_n2383;
   wire FE_PHN6773_n3992;
   wire FE_PHN6772_n4203;
   wire FE_PHN6771_n1038;
   wire FE_PHN6770_n4000;
   wire FE_PHN6769_n4350;
   wire FE_PHN6768_n4194;
   wire FE_PHN6767_n4164;
   wire FE_PHN6766_n911;
   wire FE_PHN6765_n2405;
   wire FE_PHN6764_n3258;
   wire FE_PHN6763_n2945;
   wire FE_PHN6762_n4174;
   wire FE_PHN6761_n3129;
   wire FE_PHN6760_n3219;
   wire FE_PHN6759_n1920;
   wire FE_PHN6758_n2389;
   wire FE_PHN6757_n959;
   wire FE_PHN6756_n2564;
   wire FE_PHN6755_n3028;
   wire FE_PHN6754_n2420;
   wire FE_PHN6753_n928;
   wire FE_PHN6752_n905;
   wire FE_PHN6751_n3077;
   wire FE_PHN6750_n2385;
   wire FE_PHN6749_n4178;
   wire FE_PHN6748_n1014;
   wire FE_PHN6747_n4049;
   wire FE_PHN6746_n1870;
   wire FE_PHN6745_n1017;
   wire FE_PHN6744_n3072;
   wire FE_PHN6743_n4248;
   wire FE_PHN6742_n4214;
   wire FE_PHN6741_n2574;
   wire FE_PHN6740_n4334;
   wire FE_PHN6739_n2431;
   wire FE_PHN6738_n1902;
   wire FE_PHN6737_n3919;
   wire FE_PHN6736_n2415;
   wire FE_PHN6735_n4046;
   wire FE_PHN6734_n4255;
   wire FE_PHN6733_n3263;
   wire FE_PHN6732_n4343;
   wire FE_PHN6731_n3964;
   wire FE_PHN6730_n975;
   wire FE_PHN6729_n1905;
   wire FE_PHN6728_n4215;
   wire FE_PHN6727_n4180;
   wire FE_PHN6726_n946;
   wire FE_PHN6725_n2408;
   wire FE_PHN6724_n2580;
   wire FE_PHN6723_n3040;
   wire FE_PHN6722_n2599;
   wire FE_PHN6721_n948;
   wire FE_PHN6720_n954;
   wire FE_PHN6719_n1013;
   wire FE_PHN6718_n4219;
   wire FE_PHN6717_n2964;
   wire FE_PHN6716_n4229;
   wire FE_PHN6715_n1873;
   wire FE_PHN6714_n1082;
   wire FE_PHN6713_n974;
   wire FE_PHN6712_n3068;
   wire FE_PHN6711_n2133;
   wire FE_PHN6710_n2610;
   wire FE_PHN6709_n2180;
   wire FE_PHN6708_n2166;
   wire FE_PHN6707_n2167;
   wire FE_PHN6706_n2890;
   wire FE_PHN6705_n4409;
   wire FE_PHN6704_n2887;
   wire FE_PHN6703_n2126;
   wire FE_PHN6702_n4013;
   wire FE_PHN6701_n4137;
   wire FE_PHN6700_n3953;
   wire FE_PHN6699_n2120;
   wire FE_PHN6698_n3230;
   wire FE_PHN6697_n2614;
   wire FE_PHN6696_n2570;
   wire FE_PHN6695_n2179;
   wire FE_PHN6694_n2175;
   wire FE_PHN6693_n2154;
   wire FE_PHN6692_n2972;
   wire FE_PHN6691_n2155;
   wire FE_PHN6690_n2135;
   wire FE_PHN6689_n2164;
   wire FE_PHN6688_n2592;
   wire FE_PHN6687_n2394;
   wire FE_PHN6686_n4155;
   wire FE_PHN6685_n2379;
   wire FE_PHN6684_n4002;
   wire FE_PHN6683_n2604;
   wire FE_PHN6682_n2165;
   wire FE_PHN6681_n2625;
   wire FE_PHN6680_n2159;
   wire FE_PHN6679_n2132;
   wire FE_PHN6678_n4102;
   wire FE_PHN6677_n2603;
   wire FE_PHN6676_n3934;
   wire FE_PHN6675_n3960;
   wire FE_PHN6674_n1863;
   wire FE_PHN6673_n2582;
   wire FE_PHN6672_n2151;
   wire FE_PHN6671_n2119;
   wire FE_PHN6670_n2427;
   wire FE_PHN6669_n4147;
   wire FE_PHN6668_n4163;
   wire FE_PHN6667_n2628;
   wire FE_PHN6666_n4365;
   wire FE_PHN6665_n2417;
   wire FE_PHN6664_n2892;
   wire FE_PHN6663_n2393;
   wire FE_PHN6662_n2169;
   wire FE_PHN6661_n4153;
   wire FE_PHN6660_n2170;
   wire FE_PHN6659_n4139;
   wire FE_PHN6658_n2130;
   wire FE_PHN6657_n2434;
   wire FE_PHN6656_n2118;
   wire FE_PHN6655_n2426;
   wire FE_PHN6654_n3968;
   wire FE_PHN6653_n2378;
   wire FE_PHN6652_n2578;
   wire FE_PHN6651_n3923;
   wire FE_PHN6650_n2571;
   wire FE_PHN6649_n2402;
   wire FE_PHN6648_n4121;
   wire FE_PHN6647_n2425;
   wire FE_PHN6646_n2395;
   wire FE_PHN6645_n2410;
   wire FE_PHN6644_n2168;
   wire FE_PHN6643_n2377;
   wire FE_PHN6642_n4011;
   wire FE_PHN6641_n2152;
   wire FE_PHN6640_n2414;
   wire FE_PHN6639_n2397;
   wire FE_PHN6638_n2921;
   wire FE_PHN6637_n2743;
   wire FE_PHN6636_n2749;
   wire FE_PHN6635_n2122;
   wire FE_PHN6634_n2176;
   wire FE_PHN6633_n2589;
   wire FE_PHN6632_n4158;
   wire FE_PHN6631_n4062;
   wire FE_PHN6630_n3965;
   wire FE_PHN6629_n1913;
   wire FE_PHN6628_n4135;
   wire FE_PHN6627_n2697;
   wire FE_PHN6626_n3033;
   wire FE_PHN6625_n2609;
   wire FE_PHN6624_n4107;
   wire FE_PHN6623_n3944;
   wire FE_PHN6622_n2123;
   wire FE_PHN6621_n3034;
   wire FE_PHN6620_n921;
   wire FE_PHN6619_n1908;
   wire FE_PHN6618_n1375;
   wire FE_PHN6617_n2908;
   wire FE_PHN6616_n2257;
   wire FE_PHN6615_n4151;
   wire FE_PHN6614_n2624;
   wire FE_PHN6613_n1865;
   wire FE_PHN6612_n2386;
   wire FE_PHN6611_n3004;
   wire FE_PHN6610_n4150;
   wire FE_PHN6609_n2390;
   wire FE_PHN6608_n3017;
   wire FE_PHN6607_n2626;
   wire FE_PHN6606_n2422;
   wire FE_PHN6605_n2876;
   wire FE_PHN6604_n2577;
   wire FE_PHN6603_n3150;
   wire FE_PHN6602_n3047;
   wire FE_PHN6601_n2177;
   wire FE_PHN6600_n2406;
   wire FE_PHN6599_n2587;
   wire FE_PHN6598_n1012;
   wire FE_PHN6597_n985;
   wire FE_PHN6596_n973;
   wire FE_PHN6595_n2701;
   wire FE_PHN6594_n1007;
   wire FE_PHN6593_n2873;
   wire FE_PHN6592_n2919;
   wire FE_PHN6591_n2398;
   wire FE_PHN6590_n2171;
   wire FE_PHN6589_n2938;
   wire FE_PHN6588_n1003;
   wire FE_PHN6587_n1286;
   wire FE_PHN6586_n2889;
   wire FE_PHN6585_n2161;
   wire FE_PHN6584_n3021;
   wire FE_PHN6583_n1028;
   wire FE_PHN6582_n2619;
   wire FE_PHN6581_n981;
   wire FE_PHN6580_n2590;
   wire FE_PHN6579_n977;
   wire FE_PHN6578_n2893;
   wire FE_PHN6577_n2616;
   wire FE_PHN6576_n2857;
   wire FE_PHN6575_n983;
   wire FE_PHN6574_n2428;
   wire FE_PHN6573_n2907;
   wire FE_PHN6572_n1086;
   wire FE_PHN6571_n2381;
   wire FE_PHN6570_n2925;
   wire FE_PHN6569_n2941;
   wire FE_PHN6568_n896;
   wire FE_PHN6567_n2750;
   wire FE_PHN6566_n2375;
   wire FE_PHN6565_n2696;
   wire FE_PHN6564_n1158;
   wire FE_PHN6563_n4012;
   wire FE_PHN6562_n1019;
   wire FE_PHN6561_n2407;
   wire FE_PHN6560_n2181;
   wire FE_PHN6559_n996;
   wire FE_PHN6558_n1031;
   wire FE_PHN6557_n1094;
   wire FE_PHN6556_n2429;
   wire FE_PHN6555_n2566;
   wire FE_PHN6554_n2695;
   wire FE_PHN6553_n980;
   wire FE_PHN6552_n2144;
   wire FE_PHN6551_n2172;
   wire FE_PHN6550_n2125;
   wire FE_PHN6549_n2411;
   wire FE_PHN6548_n1015;
   wire FE_PHN6547_n967;
   wire FE_PHN6546_n979;
   wire FE_PHN6545_n880;
   wire FE_PHN6544_n2611;
   wire FE_PHN6543_n3945;
   wire FE_PHN6542_n4210;
   wire FE_PHN6541_n2148;
   wire FE_PHN6540_n1001;
   wire FE_PHN6539_n2747;
   wire FE_PHN6538_n2594;
   wire FE_PHN6537_n4018;
   wire FE_PHN6536_n2618;
   wire FE_PHN6535_n2424;
   wire FE_PHN6534_n1054;
   wire FE_PHN6533_n898;
   wire FE_PHN6532_n4403;
   wire FE_PHN6531_n3980;
   wire FE_PHN6530_n1154;
   wire FE_PHN6529_n3981;
   wire FE_PHN6528_n2602;
   wire FE_PHN6527_n1190;
   wire FE_PHN6526_n4016;
   wire FE_PHN6525_n962;
   wire FE_PHN6524_n2376;
   wire FE_PHN6523_n2576;
   wire FE_PHN6522_n2423;
   wire FE_PHN6521_n3932;
   wire FE_PHN6520_n4358;
   wire FE_PHN6519_n4259;
   wire FE_PHN6518_n1178;
   wire FE_PHN6517_n953;
   wire FE_PHN6516_n917;
   wire FE_PHN6515_n3962;
   wire FE_PHN6514_n2622;
   wire FE_PHN6513_n3971;
   wire FE_PHN6512_n2380;
   wire FE_PHN6511_n4274;
   wire FE_PHN6510_n2572;
   wire FE_PHN6509_n2156;
   wire FE_PHN6508_n888;
   wire FE_PHN6507_n4294;
   wire FE_PHN6506_n4114;
   wire FE_PHN6505_n949;
   wire FE_PHN6504_n4391;
   wire FE_PHN6503_n2251;
   wire FE_PHN6502_n3212;
   wire FE_PHN6501_n2412;
   wire FE_PHN6500_n4035;
   wire FE_PHN6499_n2615;
   wire FE_PHN6498_n2131;
   wire FE_PHN6497_n1872;
   wire FE_PHN6496_n4308;
   wire FE_PHN6495_n1874;
   wire FE_PHN6494_n2388;
   wire FE_PHN6493_n3970;
   wire FE_PHN6492_n4034;
   wire FE_PHN6491_n1922;
   wire FE_PHN6490_n3955;
   wire FE_PHN6489_n4404;
   wire FE_PHN6488_n4273;
   wire FE_PHN6487_n2935;
   wire FE_PHN6486_n2968;
   wire FE_PHN6485_n4374;
   wire FE_PHN6484_n3260;
   wire FE_PHN6483_n2138;
   wire FE_PHN6482_n4242;
   wire FE_PHN6481_n1906;
   wire FE_PHN6480_n1918;
   wire FE_PHN6479_n938;
   wire FE_PHN6478_n4370;
   wire FE_PHN6477_n964;
   wire FE_PHN6476_n906;
   wire FE_PHN6475_n2163;
   wire FE_PHN6474_n2598;
   wire FE_PHN6473_n950;
   wire FE_PHN6472_n901;
   wire FE_PHN6471_n2612;
   wire FE_PHN6470_n944;
   wire FE_PHN6469_n2121;
   wire FE_PHN6468_n933;
   wire FE_PHN6467_n2419;
   wire FE_PHN6466_n3983;
   wire FE_PHN6465_n2124;
   wire FE_PHN6464_n4116;
   wire FE_PHN6463_n1880;
   wire FE_PHN6462_n4032;
   wire FE_PHN6461_n3966;
   wire FE_PHN6460_n2137;
   wire FE_PHN6459_n3979;
   wire FE_PHN6458_n4148;
   wire FE_PHN6457_n2403;
   wire FE_PHN6456_n1919;
   wire FE_PHN6455_n927;
   wire FE_PHN6454_n4008;
   wire FE_PHN6453_n2904;
   wire FE_PHN6452_n2922;
   wire FE_PHN6451_n3000;
   wire FE_PHN6450_n4027;
   wire FE_PHN6449_n2985;
   wire FE_PHN6448_n2382;
   wire FE_PHN6447_n2149;
   wire FE_PHN6446_n4331;
   wire FE_PHN6445_n2401;
   wire FE_PHN6444_n2432;
   wire FE_PHN6443_n4142;
   wire FE_PHN6442_n4110;
   wire FE_PHN6441_n930;
   wire FE_PHN6440_n914;
   wire FE_PHN6439_n4031;
   wire FE_PHN6438_n2605;
   wire FE_PHN6437_n1904;
   wire FE_PHN6436_n904;
   wire FE_PHN6435_n3109;
   wire FE_PHN6434_n4123;
   wire FE_PHN6433_n4244;
   wire FE_PHN6432_n3066;
   wire FE_PHN6431_n3911;
   wire FE_PHN6430_n3005;
   wire FE_PHN6429_n4285;
   wire FE_PHN6428_n3119;
   wire FE_PHN6427_ram_98__3_;
   wire FE_PHN6426_n3030;
   wire FE_PHN6425_n2262;
   wire FE_PHN6424_n4367;
   wire FE_PHN6423_n3140;
   wire FE_PHN6422_n2891;
   wire FE_PHN6421_n4146;
   wire FE_PHN6420_n2554;
   wire FE_PHN6419_n4363;
   wire FE_PHN6418_n3036;
   wire FE_PHN6417_n3241;
   wire FE_PHN6416_n2957;
   wire FE_PHN6415_n3135;
   wire FE_PHN6414_n4265;
   wire FE_PHN6413_n2910;
   wire FE_PHN6412_n2600;
   wire FE_PHN6411_n2974;
   wire FE_PHN6410_n4175;
   wire FE_PHN6409_n3123;
   wire FE_PHN6408_n2906;
   wire FE_PHN6407_n3999;
   wire FE_PHN6406_n3011;
   wire FE_PHN6405_n1023;
   wire FE_PHN6404_n4366;
   wire FE_PHN6403_n2960;
   wire FE_PHN6402_n3046;
   wire FE_PHN6401_n841;
   wire FE_PHN6400_n3265;
   wire FE_PHN6399_n1206;
   wire FE_PHN6398_n3139;
   wire FE_PHN6397_n3090;
   wire FE_PHN6396_n4261;
   wire FE_PHN6395_ram_17__14_;
   wire FE_PHN6394_n951;
   wire FE_PHN6393_n4170;
   wire FE_PHN6392_n4187;
   wire FE_PHN6391_n3091;
   wire FE_PHN6390_n3115;
   wire FE_PHN6389_n3085;
   wire FE_PHN6388_n2963;
   wire FE_PHN6387_n4267;
   wire FE_PHN6386_n4168;
   wire FE_PHN6385_n871;
   wire FE_PHN6384_n4138;
   wire FE_PHN6383_n4241;
   wire FE_PHN6382_n4266;
   wire FE_PHN6381_n863;
   wire FE_PHN6380_n2391;
   wire FE_PHN6379_n4201;
   wire FE_PHN6378_n3031;
   wire FE_PHN6377_n4254;
   wire FE_PHN6376_n976;
   wire FE_PHN6375_n991;
   wire FE_PHN6374_n3931;
   wire FE_PHN6373_n4316;
   wire FE_PHN6372_n3132;
   wire FE_PHN6371_n3083;
   wire FE_PHN6370_n4395;
   wire FE_PHN6369_n3137;
   wire FE_PHN6368_n3117;
   wire FE_PHN6367_n4227;
   wire FE_PHN6366_n4276;
   wire FE_PHN6365_n952;
   wire FE_PHN6364_n3920;
   wire FE_PHN6363_n4231;
   wire FE_PHN6362_n4382;
   wire FE_PHN6361_n3064;
   wire FE_PHN6360_n1911;
   wire FE_PHN6359_n2990;
   wire FE_PHN6358_n3038;
   wire FE_PHN6357_n4213;
   wire FE_PHN6356_n968;
   wire FE_PHN6355_n4236;
   wire FE_PHN6354_n4375;
   wire FE_PHN6353_n3947;
   wire FE_PHN6352_n3118;
   wire FE_PHN6351_n3111;
   wire FE_PHN6350_n877;
   wire FE_PHN6349_n3065;
   wire FE_PHN6348_n4270;
   wire FE_PHN6347_n2703;
   wire FE_PHN6346_n966;
   wire FE_PHN6345_n4290;
   wire FE_PHN6344_n922;
   wire FE_PHN6343_n1016;
   wire FE_PHN6342_n2926;
   wire FE_PHN6341_n3126;
   wire FE_PHN6340_n3939;
   wire FE_PHN6339_n3089;
   wire FE_PHN6338_n4356;
   wire FE_PHN6337_n3105;
   wire FE_PHN6336_n4420;
   wire FE_PHN6335_n1864;
   wire FE_PHN6334_ram_237__7_;
   wire FE_PHN6333_n4286;
   wire FE_PHN6332_n909;
   wire FE_PHN6331_n4412;
   wire FE_PHN6330_n3008;
   wire FE_PHN6329_n3917;
   wire FE_PHN6328_n4384;
   wire FE_PHN6327_n2966;
   wire FE_PHN6326_n4406;
   wire FE_PHN6325_n4414;
   wire FE_PHN6324_n4181;
   wire FE_PHN6323_n3058;
   wire FE_PHN6322_n3223;
   wire FE_PHN6321_n3127;
   wire FE_PHN6320_n3141;
   wire FE_PHN6319_ram_158__11_;
   wire FE_PHN6318_n4025;
   wire FE_PHN6317_n3950;
   wire FE_PHN6316_n843;
   wire FE_PHN6315_n4368;
   wire FE_PHN6314_n958;
   wire FE_PHN6313_n2898;
   wire FE_PHN6312_n4218;
   wire FE_PHN6311_n4171;
   wire FE_PHN6310_n850;
   wire FE_PHN6309_n4383;
   wire FE_PHN6308_n3099;
   wire FE_PHN6307_n1024;
   wire FE_PHN6306_n1002;
   wire FE_PHN6305_n3138;
   wire FE_PHN6304_n4094;
   wire FE_PHN6303_n4212;
   wire FE_PHN6302_n4283;
   wire FE_PHN6301_n3015;
   wire FE_PHN6300_n3918;
   wire FE_PHN6299_n1000;
   wire FE_PHN6298_n3114;
   wire FE_PHN6297_n4364;
   wire FE_PHN6296_n934;
   wire FE_PHN6295_n4103;
   wire FE_PHN6294_n4023;
   wire FE_PHN6293_n1029;
   wire FE_PHN6292_n4166;
   wire FE_PHN6291_n3026;
   wire FE_PHN6290_n3120;
   wire FE_PHN6289_n4185;
   wire FE_PHN6288_n895;
   wire FE_PHN6287_n847;
   wire FE_PHN6286_n4398;
   wire FE_PHN6285_n1062;
   wire FE_PHN6284_n4396;
   wire FE_PHN6283_n4373;
   wire FE_PHN6282_n2413;
   wire FE_PHN6281_n997;
   wire FE_PHN6280_n3946;
   wire FE_PHN6279_n986;
   wire FE_PHN6278_n886;
   wire FE_PHN6277_n4372;
   wire FE_PHN6276_n869;
   wire FE_PHN6275_n4245;
   wire FE_PHN6274_n960;
   wire FE_PHN6273_n3095;
   wire FE_PHN6272_n4269;
   wire FE_PHN6271_n978;
   wire FE_PHN6270_n4134;
   wire FE_PHN6269_ram_31__2_;
   wire FE_PHN6268_ram_145__1_;
   wire FE_PHN6267_n1916;
   wire FE_PHN6266_n3012;
   wire FE_PHN6265_n1921;
   wire FE_PHN6264_n3042;
   wire FE_PHN6263_n3032;
   wire FE_PHN6262_n854;
   wire FE_PHN6261_n3133;
   wire FE_PHN6260_n4097;
   wire FE_PHN6259_n3062;
   wire FE_PHN6258_n2986;
   wire FE_PHN6257_n3262;
   wire FE_PHN6256_n849;
   wire FE_PHN6255_n3035;
   wire FE_PHN6254_n1008;
   wire FE_PHN6253_n2982;
   wire FE_PHN6252_n2297;
   wire FE_PHN6251_n3922;
   wire FE_PHN6250_n3100;
   wire FE_PHN6249_n4003;
   wire FE_PHN6248_ram_221__1_;
   wire FE_PHN6247_n4339;
   wire FE_PHN6246_n993;
   wire FE_PHN6245_n947;
   wire FE_PHN6244_n3084;
   wire FE_PHN6243_n4233;
   wire FE_PHN6242_n2952;
   wire FE_PHN6241_n919;
   wire FE_PHN6240_n3080;
   wire FE_PHN6239_n3054;
   wire FE_PHN6238_n3094;
   wire FE_PHN6237_n897;
   wire FE_PHN6236_n3014;
   wire FE_PHN6235_n845;
   wire FE_PHN6234_n1005;
   wire FE_PHN6233_n3130;
   wire FE_PHN6232_n3125;
   wire FE_PHN6231_n1042;
   wire FE_PHN6230_n4167;
   wire FE_PHN6229_n3110;
   wire FE_PHN6228_n3092;
   wire FE_PHN6227_n3063;
   wire FE_PHN6226_n3078;
   wire FE_PHN6225_n3108;
   wire FE_PHN6224_n4289;
   wire FE_PHN6223_n4235;
   wire FE_PHN6222_n4199;
   wire FE_PHN6221_n2258;
   wire FE_PHN6220_n3104;
   wire FE_PHN6219_ram_20__10_;
   wire FE_PHN6218_n3102;
   wire FE_PHN6217_n3124;
   wire FE_PHN6216_n4238;
   wire FE_PHN6215_n4397;
   wire FE_PHN6214_n1018;
   wire FE_PHN6213_n2896;
   wire FE_PHN6212_ram_238__0_;
   wire FE_PHN6211_n3001;
   wire FE_PHN6210_n903;
   wire FE_PHN6209_n2886;
   wire FE_PHN6208_n4327;
   wire FE_PHN6207_n4388;
   wire FE_PHN6206_n4076;
   wire FE_PHN6205_n2158;
   wire FE_PHN6204_n838;
   wire FE_PHN6203_n1068;
   wire FE_PHN6202_n4179;
   wire FE_PHN6201_n2753;
   wire FE_PHN6200_n4026;
   wire FE_PHN6199_n4329;
   wire FE_PHN6198_n882;
   wire FE_PHN6197_n2959;
   wire FE_PHN6196_n3079;
   wire FE_PHN6195_n844;
   wire FE_PHN6194_n3940;
   wire FE_PHN6193_n2928;
   wire FE_PHN6192_n3952;
   wire FE_PHN6191_n4230;
   wire FE_PHN6190_n4333;
   wire FE_PHN6189_n3074;
   wire FE_PHN6188_n3936;
   wire FE_PHN6187_n3914;
   wire FE_PHN6186_n3985;
   wire FE_PHN6185_n918;
   wire FE_PHN6184_n2933;
   wire FE_PHN6183_n3122;
   wire FE_PHN6182_n3136;
   wire FE_PHN6181_n3974;
   wire FE_PHN6180_n3989;
   wire FE_PHN6179_n3003;
   wire FE_PHN6178_n982;
   wire FE_PHN6177_n2127;
   wire FE_PHN6176_n4416;
   wire FE_PHN6175_n1064;
   wire FE_PHN6174_n2993;
   wire FE_PHN6173_n3096;
   wire FE_PHN6172_n3951;
   wire FE_PHN6171_n2965;
   wire FE_PHN6170_n2396;
   wire FE_PHN6169_n4408;
   wire FE_PHN6168_n3954;
   wire FE_PHN6167_n4228;
   wire FE_PHN6166_n4417;
   wire FE_PHN6165_ram_214__13_;
   wire FE_PHN6164_n3006;
   wire FE_PHN6163_n4196;
   wire FE_PHN6162_n865;
   wire FE_PHN6161_n3013;
   wire FE_PHN6160_n4239;
   wire FE_PHN6159_n2973;
   wire FE_PHN6158_n1088;
   wire FE_PHN6157_n3942;
   wire FE_PHN6156_n1899;
   wire FE_PHN6155_n3019;
   wire FE_PHN6154_n3088;
   wire FE_PHN6153_n3961;
   wire FE_PHN6152_n3086;
   wire FE_PHN6151_n2991;
   wire FE_PHN6150_n2920;
   wire FE_PHN6149_n992;
   wire FE_PHN6148_n4281;
   wire FE_PHN6147_n2969;
   wire FE_PHN6146_n4271;
   wire FE_PHN6145_n969;
   wire FE_PHN6144_n874;
   wire FE_PHN6143_n2918;
   wire FE_PHN6142_n4415;
   wire FE_PHN6141_n3070;
   wire FE_PHN6140_n902;
   wire FE_PHN6139_n2141;
   wire FE_PHN6138_n3069;
   wire FE_PHN6137_n885;
   wire FE_PHN6136_n900;
   wire FE_PHN6135_n3210;
   wire FE_PHN6134_n4202;
   wire FE_PHN6133_n1026;
   wire FE_PHN6132_n3972;
   wire FE_PHN6131_n2984;
   wire FE_PHN6130_n2977;
   wire FE_PHN6129_n3107;
   wire FE_PHN6128_n3087;
   wire FE_PHN6127_n2979;
   wire FE_PHN6126_n2934;
   wire FE_PHN6125_n4394;
   wire FE_PHN6124_n3009;
   wire FE_PHN6123_n4380;
   wire FE_PHN6122_n2997;
   wire FE_PHN6121_n3050;
   wire FE_PHN6120_n2980;
   wire FE_PHN6119_n3921;
   wire FE_PHN6118_n4300;
   wire FE_PHN6117_n853;
   wire FE_PHN6116_n2946;
   wire FE_PHN6115_ram_229__12_;
   wire FE_PHN6114_n4169;
   wire FE_PHN6113_n3956;
   wire FE_PHN6112_n3024;
   wire FE_PHN6111_n3993;
   wire FE_PHN6110_n899;
   wire FE_PHN6109_n4262;
   wire FE_PHN6108_n3116;
   wire FE_PHN6107_n839;
   wire FE_PHN6106_n4284;
   wire FE_PHN6105_n4402;
   wire FE_PHN6104_n1074;
   wire FE_PHN6103_n2981;
   wire FE_PHN6102_ram_153__7_;
   wire FE_PHN6101_n2621;
   wire FE_PHN6100_n984;
   wire FE_PHN6099_n4111;
   wire FE_PHN6098_n1020;
   wire FE_PHN6097_n3959;
   wire FE_PHN6096_n2983;
   wire FE_PHN6095_n2996;
   wire FE_PHN6094_n3977;
   wire FE_PHN6093_n4007;
   wire FE_PHN6092_n3103;
   wire FE_PHN6091_n2944;
   wire FE_PHN6090_n4022;
   wire FE_PHN6089_n3975;
   wire FE_PHN6088_n2954;
   wire FE_PHN6087_n1009;
   wire FE_PHN6086_n2975;
   wire FE_PHN6085_n2888;
   wire FE_PHN6084_n4291;
   wire FE_PHN6083_n2916;
   wire FE_PHN6082_n1032;
   wire FE_PHN6081_n961;
   wire FE_PHN6080_n3044;
   wire FE_PHN6079_n4183;
   wire FE_PHN6078_n1077;
   wire FE_PHN6077_n3943;
   wire FE_PHN6076_n4386;
   wire FE_PHN6075_n3007;
   wire FE_PHN6074_n4251;
   wire FE_PHN6073_n3969;
   wire FE_PHN6072_n4222;
   wire FE_PHN6071_n4037;
   wire FE_PHN6070_n970;
   wire FE_PHN6069_n3998;
   wire FE_PHN6068_n3022;
   wire FE_PHN6067_n3255;
   wire FE_PHN6066_n3924;
   wire FE_PHN6065_n2953;
   wire FE_PHN6064_ram_145__7_;
   wire FE_PHN6063_n4204;
   wire FE_PHN6062_n3081;
   wire FE_PHN6061_n1072;
   wire FE_PHN6060_n1048;
   wire FE_PHN6059_n3112;
   wire FE_PHN6058_n2950;
   wire FE_PHN6057_n1896;
   wire FE_PHN6056_n4006;
   wire FE_PHN6055_n3996;
   wire FE_PHN6054_n3067;
   wire FE_PHN6053_n4260;
   wire FE_PHN6052_n941;
   wire FE_PHN6051_n3098;
   wire FE_PHN6050_n999;
   wire FE_PHN6049_n4279;
   wire FE_PHN6048_n856;
   wire FE_PHN6047_n3982;
   wire FE_PHN6046_n1025;
   wire FE_PHN6045_n887;
   wire FE_PHN6044_n1021;
   wire FE_PHN6043_n3910;
   wire FE_PHN6042_n4203;
   wire FE_PHN6041_n3134;
   wire FE_PHN6040_n2943;
   wire FE_PHN6039_n4332;
   wire FE_PHN6038_n4211;
   wire FE_PHN6037_n1066;
   wire FE_PHN6036_n3131;
   wire FE_PHN6035_n1014;
   wire FE_PHN6034_ram_145__10_;
   wire FE_PHN6033_n3060;
   wire FE_PHN6032_n998;
   wire FE_PHN6031_n890;
   wire FE_PHN6030_n989;
   wire FE_PHN6029_n1006;
   wire FE_PHN6028_n3053;
   wire FE_PHN6027_n889;
   wire FE_PHN6026_n4311;
   wire FE_PHN6025_n4418;
   wire FE_PHN6024_ram_145__0_;
   wire FE_PHN6023_n892;
   wire FE_PHN6022_n879;
   wire FE_PHN6021_ram_133__9_;
   wire FE_PHN6020_n3076;
   wire FE_PHN6019_n840;
   wire FE_PHN6018_n2976;
   wire FE_PHN6017_n3025;
   wire FE_PHN6016_n884;
   wire FE_PHN6015_n4405;
   wire FE_PHN6014_n3056;
   wire FE_PHN6013_n4419;
   wire FE_PHN6012_n2989;
   wire FE_PHN6011_n846;
   wire FE_PHN6010_n3929;
   wire FE_PHN6009_n4225;
   wire FE_PHN6008_n2994;
   wire FE_PHN6007_n4010;
   wire FE_PHN6006_n881;
   wire FE_PHN6005_n2930;
   wire FE_PHN6004_n4379;
   wire FE_PHN6003_n4360;
   wire FE_PHN6002_n1045;
   wire FE_PHN6001_n3093;
   wire FE_PHN6000_n893;
   wire FE_PHN5999_n848;
   wire FE_PHN5998_n3958;
   wire FE_PHN5997_n870;
   wire FE_PHN5996_n866;
   wire FE_PHN5995_n4009;
   wire FE_PHN5994_n1110;
   wire FE_PHN5993_n2992;
   wire FE_PHN5992_n2995;
   wire FE_PHN5991_n994;
   wire FE_PHN5990_n3976;
   wire FE_PHN5989_n3023;
   wire FE_PHN5988_n4188;
   wire FE_PHN5987_n3010;
   wire FE_PHN5986_ram_153__11_;
   wire FE_PHN5985_n2970;
   wire FE_PHN5984_n3987;
   wire FE_PHN5983_n913;
   wire FE_PHN5982_n1040;
   wire FE_PHN5981_n2961;
   wire FE_PHN5980_n3129;
   wire FE_PHN5979_n3984;
   wire FE_PHN5978_n3027;
   wire FE_PHN5977_n2978;
   wire FE_PHN5976_n3018;
   wire FE_PHN5975_n2374;
   wire FE_PHN5974_n4030;
   wire FE_PHN5973_n2430;
   wire FE_PHN5972_n876;
   wire FE_PHN5971_n4401;
   wire FE_PHN5970_n957;
   wire FE_PHN5969_n4172;
   wire FE_PHN5968_n2897;
   wire FE_PHN5967_n3916;
   wire FE_PHN5966_n3128;
   wire FE_PHN5965_n3978;
   wire FE_PHN5964_n4195;
   wire FE_PHN5963_n2998;
   wire FE_PHN5962_n943;
   wire FE_PHN5961_n4217;
   wire FE_PHN5960_n3075;
   wire FE_PHN5959_n4389;
   wire FE_PHN5958_n4355;
   wire FE_PHN5957_n929;
   wire FE_PHN5956_n4340;
   wire FE_PHN5955_n4219;
   wire FE_PHN5954_n1079;
   wire FE_PHN5953_n861;
   wire FE_PHN5952_n3020;
   wire FE_PHN5951_n3082;
   wire FE_PHN5950_n4295;
   wire FE_PHN5949_n4399;
   wire FE_PHN5948_n3963;
   wire FE_PHN5947_n1013;
   wire FE_PHN5946_n3029;
   wire FE_PHN5945_n4021;
   wire FE_PHN5944_n4263;
   wire FE_PHN5943_n3002;
   wire FE_PHN5942_n2987;
   wire FE_PHN5941_n3028;
   wire FE_PHN5940_n4029;
   wire FE_PHN5939_n3048;
   wire FE_PHN5938_n4243;
   wire FE_PHN5937_n4369;
   wire FE_PHN5936_n2735;
   wire FE_PHN5935_n4378;
   wire FE_PHN5934_n4033;
   wire FE_PHN5933_n911;
   wire FE_PHN5932_n4400;
   wire FE_PHN5931_n2962;
   wire FE_PHN5930_n3055;
   wire FE_PHN5929_n4240;
   wire FE_PHN5928_n4220;
   wire FE_PHN5927_n4421;
   wire FE_PHN5926_n975;
   wire FE_PHN5925_n1037;
   wire FE_PHN5924_n2722;
   wire FE_PHN5923_n3257;
   wire FE_PHN5922_n3258;
   wire FE_PHN5921_n3043;
   wire FE_PHN5920_n864;
   wire FE_PHN5919_n965;
   wire FE_PHN5918_n1090;
   wire FE_PHN5917_n4028;
   wire FE_PHN5916_n1030;
   wire FE_PHN5915_n3964;
   wire FE_PHN5914_n4324;
   wire FE_PHN5913_n4361;
   wire FE_PHN5912_n857;
   wire FE_PHN5911_n4215;
   wire FE_PHN5910_n3915;
   wire FE_PHN5909_n4164;
   wire FE_PHN5908_n4180;
   wire FE_PHN5907_n4299;
   wire FE_PHN5906_n910;
   wire FE_PHN5905_n3937;
   wire FE_PHN5904_n2964;
   wire FE_PHN5903_n2936;
   wire FE_PHN5902_n855;
   wire FE_PHN5901_n3207;
   wire FE_PHN5900_n1056;
   wire FE_PHN5899_n3926;
   wire FE_PHN5898_n4252;
   wire FE_PHN5897_n2754;
   wire FE_PHN5896_n4377;
   wire FE_PHN5895_n1051;
   wire FE_PHN5894_n2420;
   wire FE_PHN5893_n4226;
   wire FE_PHN5892_n4017;
   wire FE_PHN5891_n925;
   wire FE_PHN5890_n3948;
   wire FE_PHN5889_n3994;
   wire FE_PHN5888_n3049;
   wire FE_PHN5887_n4209;
   wire FE_PHN5886_n2958;
   wire FE_PHN5885_n4014;
   wire FE_PHN5884_n935;
   wire FE_PHN5883_n858;
   wire FE_PHN5882_n905;
   wire FE_PHN5881_n2564;
   wire FE_PHN5880_n2927;
   wire FE_PHN5879_n3052;
   wire FE_PHN5878_ram_144__8_;
   wire FE_PHN5877_n3992;
   wire FE_PHN5876_n4307;
   wire FE_PHN5875_n4385;
   wire FE_PHN5874_n2384;
   wire FE_PHN5873_n1920;
   wire FE_PHN5872_n1034;
   wire FE_PHN5871_n988;
   wire FE_PHN5870_n3927;
   wire FE_PHN5869_n851;
   wire FE_PHN5868_n4178;
   wire FE_PHN5867_n1106;
   wire FE_PHN5866_n945;
   wire FE_PHN5865_n894;
   wire FE_PHN5864_n852;
   wire FE_PHN5863_n1093;
   wire FE_PHN5862_n842;
   wire FE_PHN5861_n2385;
   wire FE_PHN5860_n4393;
   wire FE_PHN5859_n959;
   wire FE_PHN5858_n4277;
   wire FE_PHN5857_n4194;
   wire FE_PHN5856_n4046;
   wire FE_PHN5855_n4387;
   wire FE_PHN5854_n2955;
   wire FE_PHN5853_n1022;
   wire FE_PHN5852_n4350;
   wire FE_PHN5851_n1017;
   wire FE_PHN5850_n2178;
   wire FE_PHN5849_n2932;
   wire FE_PHN5848_n2956;
   wire FE_PHN5847_n3930;
   wire FE_PHN5846_n3071;
   wire FE_PHN5845_n2951;
   wire FE_PHN5844_n3988;
   wire FE_PHN5843_n2574;
   wire FE_PHN5842_n972;
   wire FE_PHN5841_n3072;
   wire FE_PHN5840_n2971;
   wire FE_PHN5839_n2405;
   wire FE_PHN5838_n2945;
   wire FE_PHN5837_n1087;
   wire FE_PHN5836_n1069;
   wire FE_PHN5835_n3073;
   wire FE_PHN5834_n2580;
   wire FE_PHN5833_n3040;
   wire FE_PHN5832_n4174;
   wire FE_PHN5831_n4334;
   wire FE_PHN5830_n4005;
   wire FE_PHN5829_n4323;
   wire FE_PHN5828_n2900;
   wire FE_PHN5827_n878;
   wire FE_PHN5826_n4001;
   wire FE_PHN5825_n4049;
   wire FE_PHN5824_n4278;
   wire FE_PHN5823_n4214;
   wire FE_PHN5822_n1870;
   wire FE_PHN5821_n4410;
   wire FE_PHN5820_n4232;
   wire FE_PHN5819_n2421;
   wire FE_PHN5818_n4359;
   wire FE_PHN5817_n4036;
   wire FE_PHN5816_n2383;
   wire FE_PHN5815_n4362;
   wire FE_PHN5814_n2437;
   wire FE_PHN5813_n4407;
   wire FE_PHN5812_n3919;
   wire FE_PHN5811_n1082;
   wire FE_PHN5810_n872;
   wire FE_PHN5809_n4371;
   wire FE_PHN5808_n4255;
   wire FE_PHN5807_n3219;
   wire FE_PHN5806_n948;
   wire FE_PHN5805_n4248;
   wire FE_PHN5804_n2400;
   wire FE_PHN5803_n1038;
   wire FE_PHN5802_n3263;
   wire FE_PHN5801_n2399;
   wire FE_PHN5800_n936;
   wire FE_PHN5799_n2389;
   wire FE_PHN5798_n2433;
   wire FE_PHN5797_n891;
   wire FE_PHN5796_n1078;
   wire FE_PHN5795_n1905;
   wire FE_PHN5794_n2599;
   wire FE_PHN5793_n4343;
   wire FE_PHN5792_n974;
   wire FE_PHN5791_n1902;
   wire FE_PHN5790_n2408;
   wire FE_PHN5789_n4000;
   wire FE_PHN5788_n2623;
   wire FE_PHN5787_n4229;
   wire FE_PHN5786_n946;
   wire FE_PHN5785_n2431;
   wire FE_PHN5784_n1873;
   wire FE_PHN5783_n2967;
   wire FE_PHN5782_n954;
   wire FE_PHN5781_n2415;
   wire FE_PHN5780_n3077;
   wire FE_PHN5779_n920;
   wire FE_PHN5778_n928;
   wire FE_PHN5777_n3068;
   wire FE_PHN5776_n3017;
   wire FE_PHN5775_n2577;
   wire FE_PHN5774_n3033;
   wire FE_PHN5773_n2406;
   wire FE_PHN5772_n3047;
   wire FE_PHN5771_n2414;
   wire FE_PHN5770_n2397;
   wire FE_PHN5769_n2422;
   wire FE_PHN5768_n2938;
   wire FE_PHN5767_n2619;
   wire FE_PHN5766_n2889;
   wire FE_PHN5765_n1913;
   wire FE_PHN5764_n2921;
   wire FE_PHN5763_n4135;
   wire FE_PHN5762_n1908;
   wire FE_PHN5761_n2697;
   wire FE_PHN5760_n1375;
   wire FE_PHN5759_n921;
   wire FE_PHN5758_n4151;
   wire FE_PHN5757_n1865;
   wire FE_PHN5756_n2908;
   wire FE_PHN5755_n2624;
   wire FE_PHN5754_n2386;
   wire FE_PHN5753_n4150;
   wire FE_PHN5752_n2390;
   wire FE_PHN5751_n2626;
   wire FE_PHN5750_n1012;
   wire FE_PHN5749_n2919;
   wire FE_PHN5748_n2587;
   wire FE_PHN5747_n2398;
   wire FE_PHN5746_n1003;
   wire FE_PHN5745_n973;
   wire FE_PHN5744_n2893;
   wire FE_PHN5743_n1007;
   wire FE_PHN5742_n2381;
   wire FE_PHN5741_n2907;
   wire FE_PHN5740_n981;
   wire FE_PHN5739_n1028;
   wire FE_PHN5738_n2941;
   wire FE_PHN5737_n2181;
   wire FE_PHN5736_n2172;
   wire FE_PHN5735_n3021;
   wire FE_PHN5734_n2925;
   wire FE_PHN5733_n983;
   wire FE_PHN5732_n4012;
   wire FE_PHN5731_n1142;
   wire FE_PHN5730_n2611;
   wire FE_PHN5729_n1094;
   wire FE_PHN5728_n2618;
   wire FE_PHN5727_n2747;
   wire FE_PHN5726_n985;
   wire FE_PHN5725_n977;
   wire FE_PHN5724_n2125;
   wire FE_PHN5723_n1019;
   wire FE_PHN5722_n2602;
   wire FE_PHN5721_n2594;
   wire FE_PHN5720_n2424;
   wire FE_PHN5719_n2376;
   wire FE_PHN5718_n2696;
   wire FE_PHN5717_n1031;
   wire FE_PHN5716_n996;
   wire FE_PHN5715_n2576;
   wire FE_PHN5714_n2423;
   wire FE_PHN5713_n3034;
   wire FE_PHN5712_n1001;
   wire FE_PHN5711_n2251;
   wire FE_PHN5710_n2148;
   wire FE_PHN5709_n3981;
   wire FE_PHN5708_n2695;
   wire FE_PHN5707_n2740;
   wire FE_PHN5706_n2380;
   wire FE_PHN5705_n953;
   wire FE_PHN5704_n2412;
   wire FE_PHN5703_n2156;
   wire FE_PHN5702_n2572;
   wire FE_PHN5701_n2615;
   wire FE_PHN5700_n2622;
   wire FE_PHN5699_n2138;
   wire FE_PHN5698_n3965;
   wire FE_PHN5697_n1158;
   wire FE_PHN5696_n980;
   wire FE_PHN5695_n4018;
   wire FE_PHN5694_n2257;
   wire FE_PHN5693_n1086;
   wire FE_PHN5692_n2566;
   wire FE_PHN5691_n1178;
   wire FE_PHN5690_n2124;
   wire FE_PHN5689_n2743;
   wire FE_PHN5688_n3150;
   wire FE_PHN5687_n2589;
   wire FE_PHN5686_n2749;
   wire FE_PHN5685_n2873;
   wire FE_PHN5684_n2612;
   wire FE_PHN5683_n1054;
   wire FE_PHN5682_n4158;
   wire FE_PHN5681_n2876;
   wire FE_PHN5680_n3004;
   wire FE_PHN5679_n2149;
   wire FE_PHN5678_n2609;
   wire FE_PHN5677_n967;
   wire FE_PHN5676_n1190;
   wire FE_PHN5675_n4062;
   wire FE_PHN5674_n1154;
   wire FE_PHN5673_n2857;
   wire FE_PHN5672_n2590;
   wire FE_PHN5671_n1015;
   wire FE_PHN5670_n3944;
   wire FE_PHN5669_n979;
   wire FE_PHN5668_n4114;
   wire FE_PHN5667_n2616;
   wire FE_PHN5666_n2177;
   wire FE_PHN5665_n2161;
   wire FE_PHN5664_n2122;
   wire FE_PHN5663_n2750;
   wire FE_PHN5662_n2176;
   wire FE_PHN5661_n2701;
   wire FE_PHN5660_n1286;
   wire FE_PHN5659_n2382;
   wire FE_PHN5658_n2123;
   wire FE_PHN5657_n2121;
   wire FE_PHN5656_n4107;
   wire FE_PHN5655_n2144;
   wire FE_PHN5654_n2375;
   wire FE_PHN5653_n2137;
   wire FE_PHN5652_n2171;
   wire FE_PHN5651_n2407;
   wire FE_PHN5650_n2428;
   wire FE_PHN5649_n2411;
   wire FE_PHN5648_n2429;
   wire FE_PHN5647_n2401;
   wire FE_PHN5646_n2923;
   wire FE_PHN5645_n2727;
   wire FE_PHN5644_n1027;
   wire FE_PHN5643_n2733;
   wire FE_PHN5642_n2732;
   wire FE_PHN5641_n3132;
   wire FE_PHN5640_n2605;
   wire FE_PHN5639_n3117;
   wire FE_PHN5638_n4270;
   wire FE_PHN5637_n2262;
   wire FE_PHN5636_n2554;
   wire FE_PHN5635_n4123;
   wire FE_PHN5634_n3913;
   wire FE_PHN5633_n4181;
   wire FE_PHN5632_n1206;
   wire FE_PHN5631_n2600;
   wire FE_PHN5630_n4175;
   wire FE_PHN5629_n1046;
   wire FE_PHN5628_n4170;
   wire FE_PHN5627_n4015;
   wire FE_PHN5626_n971;
   wire FE_PHN5625_n3016;
   wire FE_PHN5624_n3095;
   wire FE_PHN5623_n2391;
   wire FE_PHN5622_n3111;
   wire FE_PHN5621_n2413;
   wire FE_PHN5620_n3920;
   wire FE_PHN5619_n1062;
   wire FE_PHN5618_n2926;
   wire FE_PHN5617_n4268;
   wire FE_PHN5616_n3066;
   wire FE_PHN5615_n4290;
   wire FE_PHN5614_n3036;
   wire FE_PHN5613_n2910;
   wire FE_PHN5612_n3241;
   wire FE_PHN5611_n4094;
   wire FE_PHN5610_n3911;
   wire FE_PHN5609_n1068;
   wire FE_PHN5608_n2258;
   wire FE_PHN5607_n3031;
   wire FE_PHN5606_ram_154__5_;
   wire FE_PHN5605_n2127;
   wire FE_PHN5604_n2158;
   wire FE_PHN5603_n2396;
   wire FE_PHN5602_n3083;
   wire FE_PHN5601_n3085;
   wire FE_PHN5600_n3950;
   wire FE_PHN5599_n4231;
   wire FE_PHN5598_n4097;
   wire FE_PHN5597_n2141;
   wire FE_PHN5596_ram_20__10_;
   wire FE_PHN5595_n4138;
   wire FE_PHN5594_n3917;
   wire FE_PHN5593_n4398;
   wire FE_PHN5592_n2990;
   wire FE_PHN5591_n4076;
   wire FE_PHN5590_n4292;
   wire FE_PHN5589_n4267;
   wire FE_PHN5588_n3115;
   wire FE_PHN5587_n4417;
   wire FE_PHN5586_n4265;
   wire FE_PHN5585_n4261;
   wire FE_PHN5584_n4168;
   wire FE_PHN5583_n3005;
   wire FE_PHN5582_n3114;
   wire FE_PHN5581_n4397;
   wire FE_PHN5580_n4235;
   wire FE_PHN5579_n4413;
   wire FE_PHN5578_n3081;
   wire FE_PHN5577_n3952;
   wire FE_PHN5576_n3951;
   wire FE_PHN5575_n3120;
   wire FE_PHN5574_n4254;
   wire FE_PHN5573_n3091;
   wire FE_PHN5572_n3135;
   wire FE_PHN5571_n3946;
   wire FE_PHN5570_n871;
   wire FE_PHN5569_n2999;
   wire FE_PHN5568_n3133;
   wire FE_PHN5567_n3936;
   wire FE_PHN5566_n873;
   wire FE_PHN5565_n3038;
   wire FE_PHN5564_n4236;
   wire FE_PHN5563_n4187;
   wire FE_PHN5562_ram_237__7_;
   wire FE_PHN5561_n4382;
   wire FE_PHN5560_n3030;
   wire FE_PHN5559_n884;
   wire FE_PHN5558_n4227;
   wire FE_PHN5557_n3939;
   wire FE_PHN5556_n4366;
   wire FE_PHN5555_n909;
   wire FE_PHN5554_n4103;
   wire FE_PHN5553_n838;
   wire FE_PHN5552_ram_238__0_;
   wire FE_PHN5551_n2969;
   wire FE_PHN5550_n863;
   wire FE_PHN5549_n4213;
   wire FE_PHN5548_n3062;
   wire FE_PHN5547_n4384;
   wire FE_PHN5546_n4244;
   wire FE_PHN5545_n3127;
   wire FE_PHN5544_n3100;
   wire FE_PHN5543_n1899;
   wire FE_PHN5542_n2957;
   wire FE_PHN5541_n3129;
   wire FE_PHN5540_n895;
   wire FE_PHN5539_n3008;
   wire FE_PHN5538_n3019;
   wire FE_PHN5537_n934;
   wire FE_PHN5536_n4233;
   wire FE_PHN5535_n4245;
   wire FE_PHN5534_ram_145__1_;
   wire FE_PHN5533_n4003;
   wire FE_PHN5532_ram_158__11_;
   wire FE_PHN5531_n3940;
   wire FE_PHN5530_n4291;
   wire FE_PHN5529_n3109;
   wire FE_PHN5528_ram_229__3_;
   wire FE_PHN5527_n4269;
   wire FE_PHN5526_ram_229__12_;
   wire FE_PHN5525_n2963;
   wire FE_PHN5524_n4134;
   wire FE_PHN5523_n3119;
   wire FE_PHN5522_n3099;
   wire FE_PHN5521_n3956;
   wire FE_PHN5520_n3003;
   wire FE_PHN5519_n4262;
   wire FE_PHN5518_n4406;
   wire FE_PHN5517_n4230;
   wire FE_PHN5516_n2973;
   wire FE_PHN5515_n4395;
   wire FE_PHN5514_n918;
   wire FE_PHN5513_ram_221__1_;
   wire FE_PHN5512_n4367;
   wire FE_PHN5511_n3080;
   wire FE_PHN5510_n2965;
   wire FE_PHN5509_n4420;
   wire FE_PHN5508_n2886;
   wire FE_PHN5507_n2928;
   wire FE_PHN5506_n2896;
   wire FE_PHN5505_n2918;
   wire FE_PHN5504_n4295;
   wire FE_PHN5503_n3084;
   wire FE_PHN5502_n3001;
   wire FE_PHN5501_n1896;
   wire FE_PHN5500_n2974;
   wire FE_PHN5499_n3922;
   wire FE_PHN5498_n3046;
   wire FE_PHN5497_n3032;
   wire FE_PHN5496_n4171;
   wire FE_PHN5495_n4414;
   wire FE_PHN5494_n845;
   wire FE_PHN5493_n3058;
   wire FE_PHN5492_n4339;
   wire FE_PHN5491_n3035;
   wire FE_PHN5490_n1023;
   wire FE_PHN5489_n854;
   wire FE_PHN5488_n4276;
   wire FE_PHN5487_n3088;
   wire FE_PHN5486_n3954;
   wire FE_PHN5485_n2920;
   wire FE_PHN5484_n4239;
   wire FE_PHN5483_n843;
   wire FE_PHN5482_n3096;
   wire FE_PHN5481_n3123;
   wire FE_PHN5480_ram_17__14_;
   wire FE_PHN5479_n4238;
   wire FE_PHN5478_n4202;
   wire FE_PHN5477_n968;
   wire FE_PHN5476_ram_214__13_;
   wire FE_PHN5475_n3102;
   wire FE_PHN5474_n3914;
   wire FE_PHN5473_n3078;
   wire FE_PHN5472_n2944;
   wire FE_PHN5471_n1066;
   wire FE_PHN5470_n4195;
   wire FE_PHN5469_n874;
   wire FE_PHN5468_n4388;
   wire FE_PHN5467_n886;
   wire FE_PHN5466_n844;
   wire FE_PHN5465_n900;
   wire FE_PHN5464_n3044;
   wire FE_PHN5463_n4228;
   wire FE_PHN5462_n4412;
   wire FE_PHN5461_n4329;
   wire FE_PHN5460_n3110;
   wire FE_PHN5459_n2934;
   wire FE_PHN5458_n4201;
   wire FE_PHN5457_n2898;
   wire FE_PHN5456_n4219;
   wire FE_PHN5455_n3139;
   wire FE_PHN5454_n4169;
   wire FE_PHN5453_n4026;
   wire FE_PHN5452_n877;
   wire FE_PHN5451_n3116;
   wire FE_PHN5450_n3918;
   wire FE_PHN5449_n902;
   wire FE_PHN5448_n3094;
   wire FE_PHN5447_ram_145__7_;
   wire FE_PHN5446_n850;
   wire FE_PHN5445_n4183;
   wire FE_PHN5444_n1042;
   wire FE_PHN5443_n4240;
   wire FE_PHN5442_n2943;
   wire FE_PHN5441_n1005;
   wire FE_PHN5440_n4215;
   wire FE_PHN5439_n3141;
   wire FE_PHN5438_n839;
   wire FE_PHN5437_n847;
   wire FE_PHN5436_n3210;
   wire FE_PHN5435_n3126;
   wire FE_PHN5434_n1000;
   wire FE_PHN5433_n986;
   wire FE_PHN5432_n892;
   wire FE_PHN5431_n966;
   wire FE_PHN5430_n3972;
   wire FE_PHN5429_n869;
   wire FE_PHN5428_n3134;
   wire FE_PHN5427_n889;
   wire FE_PHN5426_n3011;
   wire FE_PHN5425_n3959;
   wire FE_PHN5424_n3112;
   wire FE_PHN5423_n3108;
   wire FE_PHN5422_n856;
   wire FE_PHN5421_n3976;
   wire FE_PHN5420_n4164;
   wire FE_PHN5419_n1021;
   wire FE_PHN5418_n4211;
   wire FE_PHN5417_n3013;
   wire FE_PHN5416_n2986;
   wire FE_PHN5415_n3916;
   wire FE_PHN5414_n991;
   wire FE_PHN5413_n3943;
   wire FE_PHN5412_n3124;
   wire FE_PHN5411_n4212;
   wire FE_PHN5410_ram_31__2_;
   wire FE_PHN5409_n3024;
   wire FE_PHN5408_n1020;
   wire FE_PHN5407_n993;
   wire FE_PHN5406_n3070;
   wire FE_PHN5405_n2888;
   wire FE_PHN5404_n3060;
   wire FE_PHN5403_n3258;
   wire FE_PHN5402_n3137;
   wire FE_PHN5401_n3040;
   wire FE_PHN5400_n882;
   wire FE_PHN5399_n3028;
   wire FE_PHN5398_n4392;
   wire FE_PHN5397_n4355;
   wire FE_PHN5396_n969;
   wire FE_PHN5395_n4225;
   wire FE_PHN5394_n4364;
   wire FE_PHN5393_n4188;
   wire FE_PHN5392_n3993;
   wire FE_PHN5391_n4209;
   wire FE_PHN5390_n4222;
   wire FE_PHN5389_n2995;
   wire FE_PHN5388_n3989;
   wire FE_PHN5387_n3118;
   wire FE_PHN5386_ram_133__9_;
   wire FE_PHN5385_n976;
   wire FE_PHN5384_n3130;
   wire FE_PHN5383_n4029;
   wire FE_PHN5382_n4179;
   wire FE_PHN5381_n911;
   wire FE_PHN5380_n3255;
   wire FE_PHN5379_n2916;
   wire FE_PHN5378_n3140;
   wire FE_PHN5377_n1014;
   wire FE_PHN5376_n3022;
   wire FE_PHN5375_n4396;
   wire FE_PHN5374_n3090;
   wire FE_PHN5373_n4251;
   wire FE_PHN5372_n4373;
   wire FE_PHN5371_n1024;
   wire FE_PHN5370_n3015;
   wire FE_PHN5369_n4226;
   wire FE_PHN5368_n3964;
   wire FE_PHN5367_n4178;
   wire FE_PHN5366_n4167;
   wire FE_PHN5365_n1016;
   wire FE_PHN5364_n4172;
   wire FE_PHN5363_n2984;
   wire FE_PHN5362_n4394;
   wire FE_PHN5361_n2420;
   wire FE_PHN5360_n4199;
   wire FE_PHN5359_n4023;
   wire FE_PHN5358_n903;
   wire FE_PHN5357_n2564;
   wire FE_PHN5356_n2959;
   wire FE_PHN5355_n866;
   wire FE_PHN5354_n3910;
   wire FE_PHN5353_n4030;
   wire FE_PHN5352_n3942;
   wire FE_PHN5351_n3014;
   wire FE_PHN5350_n861;
   wire FE_PHN5349_n4311;
   wire FE_PHN5348_n2580;
   wire FE_PHN5347_n2970;
   wire FE_PHN5346_n858;
   wire FE_PHN5345_n4368;
   wire FE_PHN5344_n4340;
   wire FE_PHN5343_n2997;
   wire FE_PHN5342_n849;
   wire FE_PHN5341_n997;
   wire FE_PHN5340_n2993;
   wire FE_PHN5339_n4402;
   wire FE_PHN5338_n3136;
   wire FE_PHN5337_n4046;
   wire FE_PHN5336_n4283;
   wire FE_PHN5335_n2754;
   wire FE_PHN5334_n4418;
   wire FE_PHN5333_n2992;
   wire FE_PHN5332_n4284;
   wire FE_PHN5331_n2946;
   wire FE_PHN5330_n959;
   wire FE_PHN5329_n3086;
   wire FE_PHN5328_n3098;
   wire FE_PHN5327_n3958;
   wire FE_PHN5326_n897;
   wire FE_PHN5325_n941;
   wire FE_PHN5324_n4252;
   wire FE_PHN5323_n3067;
   wire FE_PHN5322_n3131;
   wire FE_PHN5321_n2998;
   wire FE_PHN5320_n2950;
   wire FE_PHN5319_n3089;
   wire FE_PHN5318_n4281;
   wire FE_PHN5317_n3064;
   wire FE_PHN5316_n4408;
   wire FE_PHN5315_n885;
   wire FE_PHN5314_n3025;
   wire FE_PHN5313_n4185;
   wire FE_PHN5312_n3042;
   wire FE_PHN5311_n2753;
   wire FE_PHN5310_n4416;
   wire FE_PHN5309_n4166;
   wire FE_PHN5308_n4204;
   wire FE_PHN5307_n1013;
   wire FE_PHN5306_n1006;
   wire FE_PHN5305_n3125;
   wire FE_PHN5304_n4415;
   wire FE_PHN5303_n840;
   wire FE_PHN5302_n3963;
   wire FE_PHN5301_n3087;
   wire FE_PHN5300_n3105;
   wire FE_PHN5299_n4299;
   wire FE_PHN5298_n4203;
   wire FE_PHN5297_n2178;
   wire FE_PHN5296_n2297;
   wire FE_PHN5295_n3924;
   wire FE_PHN5294_n3985;
   wire FE_PHN5293_n876;
   wire FE_PHN5292_n4360;
   wire FE_PHN5291_n4007;
   wire FE_PHN5290_n2405;
   wire FE_PHN5289_n3023;
   wire FE_PHN5288_n4350;
   wire FE_PHN5287_n913;
   wire FE_PHN5286_n3103;
   wire FE_PHN5285_n4196;
   wire FE_PHN5284_n3257;
   wire FE_PHN5283_n975;
   wire FE_PHN5282_n2936;
   wire FE_PHN5281_n943;
   wire FE_PHN5280_n957;
   wire FE_PHN5279_n3138;
   wire FE_PHN5278_n2954;
   wire FE_PHN5277_n1079;
   wire FE_PHN5276_n1106;
   wire FE_PHN5275_n2980;
   wire FE_PHN5274_n4025;
   wire FE_PHN5273_ram_153__11_;
   wire FE_PHN5272_n1018;
   wire FE_PHN5271_n881;
   wire FE_PHN5270_n2996;
   wire FE_PHN5269_n3996;
   wire FE_PHN5268_n905;
   wire FE_PHN5267_n4419;
   wire FE_PHN5266_n3065;
   wire FE_PHN5265_n4217;
   wire FE_PHN5264_n3006;
   wire FE_PHN5263_n4049;
   wire FE_PHN5262_n1920;
   wire FE_PHN5261_n3207;
   wire FE_PHN5260_n4220;
   wire FE_PHN5259_n4383;
   wire FE_PHN5258_n4277;
   wire FE_PHN5257_n4278;
   wire FE_PHN5256_n2927;
   wire FE_PHN5255_n972;
   wire FE_PHN5254_n2384;
   wire FE_PHN5253_n2897;
   wire FE_PHN5252_n1037;
   wire FE_PHN5251_n935;
   wire FE_PHN5250_n3069;
   wire FE_PHN5249_n994;
   wire FE_PHN5248_n965;
   wire FE_PHN5247_n894;
   wire FE_PHN5246_n2574;
   wire FE_PHN5245_n2987;
   wire FE_PHN5244_n3082;
   wire FE_PHN5243_n3969;
   wire FE_PHN5242_n3002;
   wire FE_PHN5241_n1870;
   wire FE_PHN5240_n2722;
   wire FE_PHN5239_n1002;
   wire FE_PHN5238_n4232;
   wire FE_PHN5237_n3029;
   wire FE_PHN5236_n841;
   wire FE_PHN5235_n4378;
   wire FE_PHN5234_n2385;
   wire FE_PHN5233_n3075;
   wire FE_PHN5232_n4316;
   wire FE_PHN5231_n3026;
   wire FE_PHN5230_n4174;
   wire FE_PHN5229_n2930;
   wire FE_PHN5228_n4206;
   wire FE_PHN5227_n4342;
   wire FE_PHN5226_n3998;
   wire FE_PHN5225_n2964;
   wire FE_PHN5224_n4400;
   wire FE_PHN5223_n929;
   wire FE_PHN5222_n4255;
   wire FE_PHN5221_ram_153__7_;
   wire FE_PHN5220_n3054;
   wire FE_PHN5219_n4380;
   wire FE_PHN5218_n3074;
   wire FE_PHN5217_n3219;
   wire FE_PHN5216_n4037;
   wire FE_PHN5215_n4286;
   wire FE_PHN5214_n3987;
   wire FE_PHN5213_n864;
   wire FE_PHN5212_n3048;
   wire FE_PHN5211_n4377;
   wire FE_PHN5210_n3020;
   wire FE_PHN5209_n948;
   wire FE_PHN5208_n988;
   wire FE_PHN5207_n2891;
   wire FE_PHN5206_n3093;
   wire FE_PHN5205_n4393;
   wire FE_PHN5204_n890;
   wire FE_PHN5203_ram_145__0_;
   wire FE_PHN5202_n982;
   wire FE_PHN5201_n3992;
   wire FE_PHN5200_n2975;
   wire FE_PHN5199_n4021;
   wire FE_PHN5198_n3055;
   wire FE_PHN5197_n2991;
   wire FE_PHN5196_n910;
   wire FE_PHN5195_n2735;
   wire FE_PHN5194_n2989;
   wire FE_PHN5193_n3104;
   wire FE_PHN5192_n887;
   wire FE_PHN5191_n1029;
   wire FE_PHN5190_n3012;
   wire FE_PHN5189_n3122;
   wire FE_PHN5188_n878;
   wire FE_PHN5187_n1017;
   wire FE_PHN5186_n936;
   wire FE_PHN5185_n3050;
   wire FE_PHN5184_n3007;
   wire FE_PHN5183_n3063;
   wire FE_PHN5182_n3919;
   wire FE_PHN5181_n3921;
   wire FE_PHN5180_n4411;
   wire FE_PHN5179_n3052;
   wire FE_PHN5178_n4363;
   wire FE_PHN5177_n4369;
   wire FE_PHN5176_n4285;
   wire FE_PHN5175_n2960;
   wire FE_PHN5174_n4014;
   wire FE_PHN5173_n846;
   wire FE_PHN5172_n1110;
   wire FE_PHN5171_n3072;
   wire FE_PHN5170_n999;
   wire FE_PHN5169_n4361;
   wire FE_PHN5168_n4333;
   wire FE_PHN5167_n4334;
   wire FE_PHN5166_n848;
   wire FE_PHN5165_n893;
   wire FE_PHN5164_n4229;
   wire FE_PHN5163_n3975;
   wire FE_PHN5162_n3053;
   wire FE_PHN5161_n3027;
   wire FE_PHN5160_n2983;
   wire FE_PHN5159_n4180;
   wire FE_PHN5158_n3974;
   wire FE_PHN5157_n4028;
   wire FE_PHN5156_n3977;
   wire FE_PHN5155_n3984;
   wire FE_PHN5154_n4241;
   wire FE_PHN5153_n2933;
   wire FE_PHN5152_n2932;
   wire FE_PHN5151_n865;
   wire FE_PHN5150_n3018;
   wire FE_PHN5149_n1077;
   wire FE_PHN5148_n925;
   wire FE_PHN5147_n870;
   wire FE_PHN5146_n4260;
   wire FE_PHN5145_n3076;
   wire FE_PHN5144_n4300;
   wire FE_PHN5143_n1038;
   wire FE_PHN5142_n4194;
   wire FE_PHN5141_n3263;
   wire FE_PHN5140_n3079;
   wire FE_PHN5139_n4327;
   wire FE_PHN5138_n1030;
   wire FE_PHN5137_n1072;
   wire FE_PHN5136_n2982;
   wire FE_PHN5135_n842;
   wire FE_PHN5134_n978;
   wire FE_PHN5133_n2951;
   wire FE_PHN5132_n3982;
   wire FE_PHN5131_n852;
   wire FE_PHN5130_n4243;
   wire FE_PHN5129_n3915;
   wire FE_PHN5128_n4214;
   wire FE_PHN5127_n4401;
   wire FE_PHN5126_n3948;
   wire FE_PHN5125_n1082;
   wire FE_PHN5124_n989;
   wire FE_PHN5123_n4279;
   wire FE_PHN5122_n879;
   wire FE_PHN5121_n4218;
   wire FE_PHN5120_n2971;
   wire FE_PHN5119_n4266;
   wire FE_PHN5118_n4338;
   wire FE_PHN5117_n3961;
   wire FE_PHN5116_n3929;
   wire FE_PHN5115_n3009;
   wire FE_PHN5114_n1069;
   wire FE_PHN5113_n1911;
   wire FE_PHN5112_n2988;
   wire FE_PHN5111_n1864;
   wire FE_PHN5110_n2621;
   wire FE_PHN5109_n2400;
   wire FE_PHN5108_n853;
   wire FE_PHN5107_n3926;
   wire FE_PHN5106_n945;
   wire FE_PHN5105_n3262;
   wire FE_PHN5104_n3092;
   wire FE_PHN5103_n3043;
   wire FE_PHN5102_n4248;
   wire FE_PHN5101_n2599;
   wire FE_PHN5100_n2945;
   wire FE_PHN5099_n1074;
   wire FE_PHN5098_n1902;
   wire FE_PHN5097_n3937;
   wire FE_PHN5096_n2976;
   wire FE_PHN5095_n946;
   wire FE_PHN5094_n1009;
   wire FE_PHN5093_n1064;
   wire FE_PHN5092_n992;
   wire FE_PHN5091_n3107;
   wire FE_PHN5090_n4386;
   wire FE_PHN5089_n1040;
   wire FE_PHN5088_n922;
   wire FE_PHN5087_n974;
   wire FE_PHN5086_n4405;
   wire FE_PHN5085_n2623;
   wire FE_PHN5084_n3049;
   wire FE_PHN5083_n3217;
   wire FE_PHN5082_n4263;
   wire FE_PHN5081_n954;
   wire FE_PHN5080_n3056;
   wire FE_PHN5079_n1886;
   wire FE_PHN5078_n1034;
   wire FE_PHN5077_n1026;
   wire FE_PHN5076_n891;
   wire FE_PHN5075_n4006;
   wire FE_PHN5074_ram_145__10_;
   wire FE_PHN5073_n1873;
   wire FE_PHN5072_n3071;
   wire FE_PHN5071_n3988;
   wire FE_PHN5070_n4289;
   wire FE_PHN5069_n1022;
   wire FE_PHN5068_n1051;
   wire FE_PHN5067_n2956;
   wire FE_PHN5066_n855;
   wire FE_PHN5065_n4010;
   wire FE_PHN5064_n2421;
   wire FE_PHN5063_n2383;
   wire FE_PHN5062_n2900;
   wire FE_PHN5061_n4385;
   wire FE_PHN5060_n4111;
   wire FE_PHN5059_n2430;
   wire FE_PHN5058_n4407;
   wire FE_PHN5057_n947;
   wire FE_PHN5056_n1905;
   wire FE_PHN5055_n1904;
   wire FE_PHN5054_n919;
   wire FE_PHN5053_n952;
   wire FE_PHN5052_n2955;
   wire FE_PHN5051_n4271;
   wire FE_PHN5050_n4410;
   wire FE_PHN5049_n4356;
   wire FE_PHN5048_n4359;
   wire FE_PHN5047_n2958;
   wire FE_PHN5046_ram_144__8_;
   wire FE_PHN5045_n1088;
   wire FE_PHN5044_n2437;
   wire FE_PHN5043_n857;
   wire FE_PHN5042_n4421;
   wire FE_PHN5041_n951;
   wire FE_PHN5040_n920;
   wire FE_PHN5039_n3930;
   wire FE_PHN5038_n1025;
   wire FE_PHN5037_n2433;
   wire FE_PHN5036_n3077;
   wire FE_PHN5035_n2399;
   wire FE_PHN5034_n872;
   wire FE_PHN5033_n904;
   wire FE_PHN5032_n4324;
   wire FE_PHN5031_n1056;
   wire FE_PHN5030_n4372;
   wire FE_PHN5029_n4036;
   wire FE_PHN5028_n1916;
   wire FE_PHN5027_n3978;
   wire FE_PHN5026_n4001;
   wire FE_PHN5025_n4017;
   wire FE_PHN5024_n3010;
   wire FE_PHN5023_n2431;
   wire FE_PHN5022_n851;
   wire FE_PHN5021_n4362;
   wire FE_PHN5020_n998;
   wire FE_PHN5019_n2703;
   wire FE_PHN5018_n1008;
   wire FE_PHN5017_n3128;
   wire FE_PHN5016_n2374;
   wire FE_PHN5015_n2389;
   wire FE_PHN5014_n4399;
   wire FE_PHN5013_n2952;
   wire FE_PHN5012_n3223;
   wire FE_PHN5011_n4375;
   wire FE_PHN5010_n4387;
   wire FE_PHN5009_n3927;
   wire FE_PHN5008_n4307;
   wire FE_PHN5007_n4033;
   wire FE_PHN5006_n1032;
   wire FE_PHN5005_n2967;
   wire FE_PHN5004_n1045;
   wire FE_PHN5003_n4146;
   wire FE_PHN5002_n4332;
   wire FE_PHN5001_n4379;
   wire FE_PHN5000_n984;
   wire FE_PHN4999_n2977;
   wire FE_PHN4998_n2994;
   wire FE_PHN4997_n3994;
   wire FE_PHN4996_n4005;
   wire FE_PHN4995_n4371;
   wire FE_PHN4994_n2981;
   wire FE_PHN4993_n4000;
   wire FE_PHN4992_n4343;
   wire FE_PHN4991_n3947;
   wire FE_PHN4990_n2953;
   wire FE_PHN4989_n3073;
   wire FE_PHN4988_n1087;
   wire FE_PHN4987_n2415;
   wire FE_PHN4986_n2978;
   wire FE_PHN4985_n4022;
   wire FE_PHN4984_n2966;
   wire FE_PHN4983_n2979;
   wire FE_PHN4982_n958;
   wire FE_PHN4981_n4389;
   wire FE_PHN4980_n2408;
   wire FE_PHN4979_n961;
   wire FE_PHN4978_n928;
   wire FE_PHN4977_n1093;
   wire FE_PHN4976_n960;
   wire FE_PHN4975_n2906;
   wire FE_PHN4974_n1921;
   wire FE_PHN4973_n3931;
   wire FE_PHN4972_n2961;
   wire FE_PHN4971_ram_98__3_;
   wire FE_PHN4970_n2962;
   wire FE_PHN4969_n1090;
   wire FE_PHN4968_n3265;
   wire FE_PHN4967_n3999;
   wire FE_PHN4966_n970;
   wire FE_PHN4965_n1048;
   wire FE_PHN4964_n4009;
   wire FE_PHN4963_n899;
   wire FE_PHN4962_n1078;
   wire FE_PHN4961_n4323;
   wire FE_PHN4960_n3150;
   wire FE_PHN4959_n1913;
   wire FE_PHN4958_n4002;
   wire FE_PHN4957_n1019;
   wire FE_PHN4956_n2155;
   wire FE_PHN4955_n2154;
   wire FE_PHN4954_n2257;
   wire FE_PHN4953_n2577;
   wire FE_PHN4952_n2740;
   wire FE_PHN4951_n1086;
   wire FE_PHN4950_n2126;
   wire FE_PHN4949_n1865;
   wire FE_PHN4948_n2172;
   wire FE_PHN4947_n2406;
   wire FE_PHN4946_n921;
   wire FE_PHN4945_n2251;
   wire FE_PHN4944_n3017;
   wire FE_PHN4943_n1012;
   wire FE_PHN4942_n4102;
   wire FE_PHN4941_n2747;
   wire FE_PHN4940_n2615;
   wire FE_PHN4939_n1178;
   wire FE_PHN4938_n2133;
   wire FE_PHN4937_n3021;
   wire FE_PHN4936_n2414;
   wire FE_PHN4935_n973;
   wire FE_PHN4934_n1190;
   wire FE_PHN4933_n1908;
   wire FE_PHN4932_n2181;
   wire FE_PHN4931_n2622;
   wire FE_PHN4930_n2610;
   wire FE_PHN4929_n1028;
   wire FE_PHN4928_n967;
   wire FE_PHN4927_n2625;
   wire FE_PHN4926_n2177;
   wire FE_PHN4925_n1286;
   wire FE_PHN4924_n2743;
   wire FE_PHN4923_n2696;
   wire FE_PHN4922_n2180;
   wire FE_PHN4921_n2175;
   wire FE_PHN4920_n977;
   wire FE_PHN4919_n1863;
   wire FE_PHN4918_n2750;
   wire FE_PHN4917_n2397;
   wire FE_PHN4916_n2876;
   wire FE_PHN4915_n2566;
   wire FE_PHN4914_n2125;
   wire FE_PHN4913_n2873;
   wire FE_PHN4912_n2611;
   wire FE_PHN4911_n2857;
   wire FE_PHN4910_n2590;
   wire FE_PHN4909_n2119;
   wire FE_PHN4908_n2378;
   wire FE_PHN4907_n1003;
   wire FE_PHN4906_n2624;
   wire FE_PHN4905_n2381;
   wire FE_PHN4904_n981;
   wire FE_PHN4903_n4147;
   wire FE_PHN4902_n1031;
   wire FE_PHN4901_n2619;
   wire FE_PHN4900_n2123;
   wire FE_PHN4899_n2921;
   wire FE_PHN4898_n979;
   wire FE_PHN4897_n2919;
   wire FE_PHN4896_n2749;
   wire FE_PHN4895_n2434;
   wire FE_PHN4894_n996;
   wire FE_PHN4893_n1054;
   wire FE_PHN4892_n2594;
   wire FE_PHN4891_n1007;
   wire FE_PHN4890_n2603;
   wire FE_PHN4889_n2614;
   wire FE_PHN4888_n2890;
   wire FE_PHN4887_n2589;
   wire FE_PHN4886_n2159;
   wire FE_PHN4885_n2572;
   wire FE_PHN4884_n2161;
   wire FE_PHN4883_n2576;
   wire FE_PHN4882_n1001;
   wire FE_PHN4881_n2423;
   wire FE_PHN4880_n2570;
   wire FE_PHN4879_n2697;
   wire FE_PHN4878_n4107;
   wire FE_PHN4877_n4013;
   wire FE_PHN4876_n1015;
   wire FE_PHN4875_n3047;
   wire FE_PHN4874_n2169;
   wire FE_PHN4873_n3230;
   wire FE_PHN4872_n1375;
   wire FE_PHN4871_n1142;
   wire FE_PHN4870_n2592;
   wire FE_PHN4869_n2422;
   wire FE_PHN4868_n2892;
   wire FE_PHN4867_n985;
   wire FE_PHN4866_n2118;
   wire FE_PHN4865_n2695;
   wire FE_PHN4864_n2889;
   wire FE_PHN4863_n1154;
   wire FE_PHN4862_n2604;
   wire FE_PHN4861_n4139;
   wire FE_PHN4860_n2166;
   wire FE_PHN4859_n2628;
   wire FE_PHN4858_n2616;
   wire FE_PHN4857_n4114;
   wire FE_PHN4856_n2701;
   wire FE_PHN4855_n2609;
   wire FE_PHN4854_n2376;
   wire FE_PHN4853_n2402;
   wire FE_PHN4852_n2612;
   wire FE_PHN4851_n2120;
   wire FE_PHN4850_n2379;
   wire FE_PHN4849_n2626;
   wire FE_PHN4848_n2386;
   wire FE_PHN4847_n2582;
   wire FE_PHN4846_n4155;
   wire FE_PHN4845_n2132;
   wire FE_PHN4844_n1094;
   wire FE_PHN4843_n2578;
   wire FE_PHN4842_n2144;
   wire FE_PHN4841_n2893;
   wire FE_PHN4840_n2165;
   wire FE_PHN4839_n2426;
   wire FE_PHN4838_n953;
   wire FE_PHN4837_n2375;
   wire FE_PHN4836_n1158;
   wire FE_PHN4835_n4135;
   wire FE_PHN4834_n980;
   wire FE_PHN4833_n2424;
   wire FE_PHN4832_n4137;
   wire FE_PHN4831_n3981;
   wire FE_PHN4830_n2382;
   wire FE_PHN4829_n2427;
   wire FE_PHN4828_n2124;
   wire FE_PHN4827_n2377;
   wire FE_PHN4826_n2122;
   wire FE_PHN4825_n2138;
   wire FE_PHN4824_n2152;
   wire FE_PHN4823_n2137;
   wire FE_PHN4822_n2121;
   wire FE_PHN4821_n2156;
   wire FE_PHN4820_n2587;
   wire FE_PHN4819_n2571;
   wire FE_PHN4818_n4150;
   wire FE_PHN4817_n3033;
   wire FE_PHN4816_n2135;
   wire FE_PHN4815_n2618;
   wire FE_PHN4814_n2390;
   wire FE_PHN4813_n2171;
   wire FE_PHN4812_n2429;
   wire FE_PHN4811_n2398;
   wire FE_PHN4810_n2938;
   wire FE_PHN4809_n2170;
   wire FE_PHN4808_n2908;
   wire FE_PHN4807_n2407;
   wire FE_PHN4806_n2148;
   wire FE_PHN4805_n4151;
   wire FE_PHN4804_n2887;
   wire FE_PHN4803_n2410;
   wire FE_PHN4802_n2393;
   wire FE_PHN4801_n2417;
   wire FE_PHN4800_n2411;
   wire FE_PHN4799_n2907;
   wire FE_PHN4798_n2401;
   wire FE_PHN4797_n2380;
   wire FE_PHN4796_n2176;
   wire FE_PHN4795_n2167;
   wire FE_PHN4794_n983;
   wire FE_PHN4793_n2602;
   wire FE_PHN4792_n2394;
   wire FE_PHN4791_n2151;
   wire FE_PHN4790_n2425;
   wire FE_PHN4789_n2164;
   wire FE_PHN4788_n2149;
   wire FE_PHN4787_n4011;
   wire FE_PHN4786_n2941;
   wire FE_PHN4785_n2179;
   wire FE_PHN4784_n4012;
   wire FE_PHN4783_n2925;
   wire FE_PHN4782_n4163;
   wire FE_PHN4781_n2412;
   wire FE_PHN4780_n4153;
   wire FE_PHN4779_n2130;
   wire FE_PHN4778_n2395;
   wire FE_PHN4777_n4121;
   wire FE_PHN4776_n4018;
   wire FE_PHN4775_n2168;
   wire FE_PHN4774_n2428;
   wire FE_PHN4773_n1027;
   wire FE_PHN4772_n2413;
   wire FE_PHN4771_n1062;
   wire FE_PHN4770_n4123;
   wire FE_PHN4769_n2262;
   wire FE_PHN4768_n2127;
   wire FE_PHN4767_n1068;
   wire FE_PHN4766_n2926;
   wire FE_PHN4765_n2258;
   wire FE_PHN4764_n971;
   wire FE_PHN4763_n2158;
   wire FE_PHN4762_n2923;
   wire FE_PHN4761_n2396;
   wire FE_PHN4760_n2141;
   wire FE_PHN4759_n2733;
   wire FE_PHN4758_n2605;
   wire FE_PHN4757_n2732;
   wire FE_PHN4756_n2727;
   wire FE_PHN4755_n3241;
   wire FE_PHN4754_n1206;
   wire FE_PHN4753_n4175;
   wire FE_PHN4752_n2600;
   wire FE_PHN4751_n4170;
   wire FE_PHN4750_n1046;
   wire FE_PHN4749_n2391;
   wire FE_PHN4748_n3920;
   wire FE_PHN4747_n2910;
   wire FE_PHN4746_n4015;
   wire FE_PHN4745_n4094;
   wire FE_PHN4744_n4097;
   wire FE_PHN4743_n3950;
   wire FE_PHN4742_n2990;
   wire FE_PHN4741_n3917;
   wire FE_PHN4740_n4265;
   wire FE_PHN4739_n4076;
   wire FE_PHN4738_n3951;
   wire FE_PHN4737_n3936;
   wire FE_PHN4736_n4236;
   wire FE_PHN4735_n3952;
   wire FE_PHN4734_n873;
   wire FE_PHN4733_n4366;
   wire FE_PHN4732_n4395;
   wire FE_PHN4731_n3135;
   wire FE_PHN4730_n4267;
   wire FE_PHN4729_n4420;
   wire FE_PHN4728_n2974;
   wire FE_PHN4727_n4087;
   wire FE_PHN4726_n4207;
   wire FE_PHN4725_n3008;
   wire FE_PHN4724_n3940;
   wire FE_PHN4723_n3062;
   wire FE_PHN4722_n838;
   wire FE_PHN4721_n4235;
   wire FE_PHN4720_n2957;
   wire FE_PHN4719_n4262;
   wire FE_PHN4718_n4233;
   wire FE_PHN4717_n3038;
   wire FE_PHN4716_n4171;
   wire FE_PHN4715_n3956;
   wire FE_PHN4714_n4202;
   wire FE_PHN4713_n4414;
   wire FE_PHN4712_n2928;
   wire FE_PHN4711_n863;
   wire FE_PHN4710_n2918;
   wire FE_PHN4709_n2886;
   wire FE_PHN4708_n3210;
   wire FE_PHN4707_n895;
   wire FE_PHN4706_n4329;
   wire FE_PHN4705_n1066;
   wire FE_PHN4704_n4215;
   wire FE_PHN4703_n4240;
   wire FE_PHN4702_n2943;
   wire FE_PHN4701_n2920;
   wire FE_PHN4700_n4209;
   wire FE_PHN4699_n892;
   wire FE_PHN4698_n839;
   wire FE_PHN4697_n854;
   wire FE_PHN4696_n843;
   wire FE_PHN4695_n4402;
   wire FE_PHN4694_n2564;
   wire FE_PHN4693_n2888;
   wire FE_PHN4692_n3126;
   wire FE_PHN4691_n3916;
   wire FE_PHN4690_n4276;
   wire FE_PHN4689_n4164;
   wire FE_PHN4688_n880;
   wire FE_PHN4687_n896;
   wire FE_PHN4686_n3258;
   wire FE_PHN4685_n4178;
   wire FE_PHN4684_n4226;
   wire FE_PHN4683_n4311;
   wire FE_PHN4682_n4222;
   wire FE_PHN4681_n911;
   wire FE_PHN4680_n4210;
   wire FE_PHN4679_n886;
   wire FE_PHN4678_n3109;
   wire FE_PHN4677_n4046;
   wire FE_PHN4676_n966;
   wire FE_PHN4675_n2970;
   wire FE_PHN4674_n3980;
   wire FE_PHN4673_n874;
   wire FE_PHN4672_n2297;
   wire FE_PHN4671_n2580;
   wire FE_PHN4670_n3932;
   wire FE_PHN4669_n3924;
   wire FE_PHN4668_n4029;
   wire FE_PHN4667_n903;
   wire FE_PHN4666_n2916;
   wire FE_PHN4665_n4412;
   wire FE_PHN4664_n1920;
   wire FE_PHN4663_n962;
   wire FE_PHN4662_n3976;
   wire FE_PHN4661_n4299;
   wire FE_PHN4660_n4364;
   wire FE_PHN4659_n3086;
   wire FE_PHN4658_n3131;
   wire FE_PHN4657_n3945;
   wire FE_PHN4656_n3044;
   wire FE_PHN4655_n2420;
   wire FE_PHN4654_n2984;
   wire FE_PHN4653_n3964;
   wire FE_PHN4652_n3255;
   wire FE_PHN4651_n2936;
   wire FE_PHN4650_n4392;
   wire FE_PHN4649_n4281;
   wire FE_PHN4648_n2963;
   wire FE_PHN4647_n850;
   wire FE_PHN4646_n3028;
   wire FE_PHN4645_n2965;
   wire FE_PHN4644_n2950;
   wire FE_PHN4643_n4227;
   wire FE_PHN4642_n4284;
   wire FE_PHN4641_n3098;
   wire FE_PHN4640_n4368;
   wire FE_PHN4639_n3020;
   wire FE_PHN4638_n4396;
   wire FE_PHN4637_n4187;
   wire FE_PHN4636_n1106;
   wire FE_PHN4635_n4268;
   wire FE_PHN4634_n2944;
   wire FE_PHN4633_n4212;
   wire FE_PHN4632_n3130;
   wire FE_PHN4631_n4252;
   wire FE_PHN4630_n2987;
   wire FE_PHN4629_n3040;
   wire FE_PHN4628_n898;
   wire FE_PHN4627_n3136;
   wire FE_PHN4626_n1870;
   wire FE_PHN4625_n1042;
   wire FE_PHN4624_n1014;
   wire FE_PHN4623_n4049;
   wire FE_PHN4622_n969;
   wire FE_PHN4621_n1023;
   wire FE_PHN4620_n4278;
   wire FE_PHN4619_n4241;
   wire FE_PHN4618_n4172;
   wire FE_PHN4617_n2927;
   wire FE_PHN4616_n4416;
   wire FE_PHN4615_n4016;
   wire FE_PHN4614_n1922;
   wire FE_PHN4613_n3958;
   wire FE_PHN4612_n2983;
   wire FE_PHN4611_n935;
   wire FE_PHN4610_n4179;
   wire FE_PHN4609_n1874;
   wire FE_PHN4608_n2986;
   wire FE_PHN4607_n993;
   wire FE_PHN4606_n1021;
   wire FE_PHN4605_n841;
   wire FE_PHN4604_n4219;
   wire FE_PHN4603_n2722;
   wire FE_PHN4602_n2384;
   wire FE_PHN4601_n877;
   wire FE_PHN4600_n2405;
   wire FE_PHN4599_n3058;
   wire FE_PHN4598_n3015;
   wire FE_PHN4597_n4232;
   wire FE_PHN4596_n2891;
   wire FE_PHN4595_n1020;
   wire FE_PHN4594_n3962;
   wire FE_PHN4593_n910;
   wire FE_PHN4592_n878;
   wire FE_PHN4591_n3139;
   wire FE_PHN4590_n889;
   wire FE_PHN4589_n4231;
   wire FE_PHN4588_n847;
   wire FE_PHN4587_n858;
   wire FE_PHN4586_n1110;
   wire FE_PHN4585_n975;
   wire FE_PHN4584_n3082;
   wire FE_PHN4583_n4021;
   wire FE_PHN4582_n2574;
   wire FE_PHN4581_n948;
   wire FE_PHN4580_n3257;
   wire FE_PHN4579_n2989;
   wire FE_PHN4578_n3052;
   wire FE_PHN4577_n991;
   wire FE_PHN4576_n4316;
   wire FE_PHN4575_n882;
   wire FE_PHN4574_n4228;
   wire FE_PHN4573_n4181;
   wire FE_PHN4572_n4259;
   wire FE_PHN4571_n2388;
   wire FE_PHN4570_n4169;
   wire FE_PHN4569_n4211;
   wire FE_PHN4568_n4277;
   wire FE_PHN4567_n4401;
   wire FE_PHN4566_n1018;
   wire FE_PHN4565_n986;
   wire FE_PHN4564_n2554;
   wire FE_PHN4563_n2992;
   wire FE_PHN4562_n4203;
   wire FE_PHN4561_n4243;
   wire FE_PHN4560_n913;
   wire FE_PHN4559_n3219;
   wire FE_PHN4558_n4183;
   wire FE_PHN4557_n905;
   wire FE_PHN4556_n1143;
   wire FE_PHN4555_n3918;
   wire FE_PHN4554_n4382;
   wire FE_PHN4553_n869;
   wire FE_PHN4552_n4418;
   wire FE_PHN4551_n3066;
   wire FE_PHN4550_n3024;
   wire FE_PHN4549_n1013;
   wire FE_PHN4548_n4026;
   wire FE_PHN4547_n4148;
   wire FE_PHN4546_n3989;
   wire FE_PHN4545_n968;
   wire FE_PHN4544_n2995;
   wire FE_PHN4543_n4168;
   wire FE_PHN4542_n972;
   wire FE_PHN4541_n3119;
   wire FE_PHN4540_n4255;
   wire FE_PHN4539_n2971;
   wire FE_PHN4538_n1872;
   wire FE_PHN4537_n1037;
   wire FE_PHN4536_n4415;
   wire FE_PHN4535_n3207;
   wire FE_PHN4534_n2933;
   wire FE_PHN4533_n1082;
   wire FE_PHN4532_n3088;
   wire FE_PHN4531_n3091;
   wire FE_PHN4530_n4037;
   wire FE_PHN4529_n2898;
   wire FE_PHN4528_n2896;
   wire FE_PHN4527_ram_158__11_;
   wire FE_PHN4526_n4116;
   wire FE_PHN4525_n3140;
   wire FE_PHN4524_n3018;
   wire FE_PHN4523_n2954;
   wire FE_PHN4522_n3942;
   wire FE_PHN4521_n3029;
   wire FE_PHN4520_n844;
   wire FE_PHN4519_n3212;
   wire FE_PHN4518_n4403;
   wire FE_PHN4517_n999;
   wire FE_PHN4516_n4294;
   wire FE_PHN4515_n4030;
   wire FE_PHN4514_n3970;
   wire FE_PHN4513_n2753;
   wire FE_PHN4512_n3069;
   wire FE_PHN4511_ram_133__9_;
   wire FE_PHN4510_n4394;
   wire FE_PHN4509_n3065;
   wire FE_PHN4508_n917;
   wire FE_PHN4507_n3137;
   wire FE_PHN4506_n2385;
   wire FE_PHN4505_n2996;
   wire FE_PHN4504_n870;
   wire FE_PHN4503_n4229;
   wire FE_PHN4502_n3913;
   wire FE_PHN4501_n3971;
   wire FE_PHN4500_n4400;
   wire FE_PHN4499_n4373;
   wire FE_PHN4498_n4355;
   wire FE_PHN4497_n2951;
   wire FE_PHN4496_n4285;
   wire FE_PHN4495_n4201;
   wire FE_PHN4494_n1017;
   wire FE_PHN4493_n3072;
   wire FE_PHN4492_n4308;
   wire FE_PHN4491_n849;
   wire FE_PHN4490_n900;
   wire FE_PHN4489_n4174;
   wire FE_PHN4488_n888;
   wire FE_PHN4487_n4350;
   wire FE_PHN4486_n2623;
   wire FE_PHN4485_n4199;
   wire FE_PHN4484_n4391;
   wire FE_PHN4483_n2946;
   wire FE_PHN4482_n3013;
   wire FE_PHN4481_n4393;
   wire FE_PHN4480_n879;
   wire FE_PHN4479_n4360;
   wire FE_PHN4478_n3076;
   wire FE_PHN4477_n4188;
   wire FE_PHN4476_n1918;
   wire FE_PHN4475_n3036;
   wire FE_PHN4474_n944;
   wire FE_PHN4473_n4334;
   wire FE_PHN4472_n4261;
   wire FE_PHN4471_n2131;
   wire FE_PHN4470_n941;
   wire FE_PHN4469_n3016;
   wire FE_PHN4468_n936;
   wire FE_PHN4467_n897;
   wire FE_PHN4466_n2998;
   wire FE_PHN4465_n3141;
   wire FE_PHN4464_n4273;
   wire FE_PHN4463_n4419;
   wire FE_PHN4462_n4300;
   wire FE_PHN4461_n3963;
   wire FE_PHN4460_n3064;
   wire FE_PHN4459_ram_20__10_;
   wire FE_PHN4458_n938;
   wire FE_PHN4457_n881;
   wire FE_PHN4456_n4270;
   wire FE_PHN4455_n1000;
   wire FE_PHN4454_n965;
   wire FE_PHN4453_n4404;
   wire FE_PHN4452_n997;
   wire FE_PHN4451_n4213;
   wire FE_PHN4450_n894;
   wire FE_PHN4449_n4032;
   wire FE_PHN4448_n2930;
   wire FE_PHN4447_n2735;
   wire FE_PHN4446_n3262;
   wire FE_PHN4445_n1034;
   wire FE_PHN4444_n861;
   wire FE_PHN4443_n988;
   wire FE_PHN4442_n2906;
   wire FE_PHN4441_ram_214__13_;
   wire FE_PHN4440_n909;
   wire FE_PHN4439_n3120;
   wire FE_PHN4438_n2598;
   wire FE_PHN4437_n4218;
   wire FE_PHN4436_n2897;
   wire FE_PHN4435_n957;
   wire FE_PHN4434_n3985;
   wire FE_PHN4433_n4166;
   wire FE_PHN4432_n3919;
   wire FE_PHN4431_n4185;
   wire FE_PHN4430_n3910;
   wire FE_PHN4429_n4180;
   wire FE_PHN4428_n1030;
   wire FE_PHN4427_n4194;
   wire FE_PHN4426_n2599;
   wire FE_PHN4425_n3969;
   wire FE_PHN4424_n2975;
   wire FE_PHN4423_n4378;
   wire FE_PHN4422_n2430;
   wire FE_PHN4421_n3075;
   wire FE_PHN4420_n3011;
   wire FE_PHN4419_n3002;
   wire FE_PHN4418_n2403;
   wire FE_PHN4417_n4206;
   wire FE_PHN4416_n4017;
   wire FE_PHN4415_n4342;
   wire FE_PHN4414_ram_31__2_;
   wire FE_PHN4413_n3996;
   wire FE_PHN4412_n4035;
   wire FE_PHN4411_n1016;
   wire FE_PHN4410_n4370;
   wire FE_PHN4409_n2997;
   wire FE_PHN4408_n2959;
   wire FE_PHN4407_n4266;
   wire FE_PHN4406_ram_153__11_;
   wire FE_PHN4405_n2993;
   wire FE_PHN4404_n3006;
   wire FE_PHN4403_n4338;
   wire FE_PHN4402_n4242;
   wire FE_PHN4401_n2922;
   wire FE_PHN4400_n1906;
   wire FE_PHN4399_n976;
   wire FE_PHN4398_n4134;
   wire FE_PHN4397_n1074;
   wire FE_PHN4396_n3055;
   wire FE_PHN4395_n2960;
   wire FE_PHN4394_n1002;
   wire FE_PHN4393_n885;
   wire FE_PHN4392_n1051;
   wire FE_PHN4391_n4027;
   wire FE_PHN4390_n4283;
   wire FE_PHN4389_n2934;
   wire FE_PHN4388_n3063;
   wire FE_PHN4387_n4271;
   wire FE_PHN4386_n4397;
   wire FE_PHN4385_n3074;
   wire FE_PHN4384_n3994;
   wire FE_PHN4383_n3974;
   wire FE_PHN4382_n3050;
   wire FE_PHN4381_n3025;
   wire FE_PHN4380_n964;
   wire FE_PHN4379_n3080;
   wire FE_PHN4378_n3992;
   wire FE_PHN4377_n4358;
   wire FE_PHN4376_n2945;
   wire FE_PHN4375_n3927;
   wire FE_PHN4374_n890;
   wire FE_PHN4373_n1022;
   wire FE_PHN4372_n3014;
   wire FE_PHN4371_n1024;
   wire FE_PHN4370_n1880;
   wire FE_PHN4369_n3263;
   wire FE_PHN4368_n1009;
   wire FE_PHN4367_n3921;
   wire FE_PHN4366_n4411;
   wire FE_PHN4365_n3961;
   wire FE_PHN4364_n4217;
   wire FE_PHN4363_n1916;
   wire FE_PHN4362_n4407;
   wire FE_PHN4361_n906;
   wire FE_PHN4360_n3122;
   wire FE_PHN4359_n2935;
   wire FE_PHN4358_ram_154__5_;
   wire FE_PHN4357_n3049;
   wire FE_PHN4356_n1899;
   wire FE_PHN4355_n974;
   wire FE_PHN4354_n949;
   wire FE_PHN4353_n2621;
   wire FE_PHN4352_n4333;
   wire FE_PHN4351_n3093;
   wire FE_PHN4350_n998;
   wire FE_PHN4349_n3079;
   wire FE_PHN4348_n3129;
   wire FE_PHN4347_n2421;
   wire FE_PHN4346_n1029;
   wire FE_PHN4345_n2399;
   wire FE_PHN4344_n4025;
   wire FE_PHN4343_n2419;
   wire FE_PHN4342_n1079;
   wire FE_PHN4341_n3975;
   wire FE_PHN4340_n933;
   wire FE_PHN4339_n891;
   wire FE_PHN4338_n904;
   wire FE_PHN4337_n4036;
   wire FE_PHN4336_n1006;
   wire FE_PHN4335_n3067;
   wire FE_PHN4334_n4369;
   wire FE_PHN4333_n851;
   wire FE_PHN4332_n3090;
   wire FE_PHN4331_n853;
   wire FE_PHN4330_n845;
   wire FE_PHN4329_n902;
   wire FE_PHN4328_n4374;
   wire FE_PHN4327_n3955;
   wire FE_PHN4326_n982;
   wire FE_PHN4325_n4248;
   wire FE_PHN4324_n840;
   wire FE_PHN4323_n3054;
   wire FE_PHN4322_n3988;
   wire FE_PHN4321_n2432;
   wire FE_PHN4320_n3984;
   wire FE_PHN4319_n2163;
   wire FE_PHN4318_n3085;
   wire FE_PHN4317_n2437;
   wire FE_PHN4316_n4386;
   wire FE_PHN4315_n994;
   wire FE_PHN4314_n2904;
   wire FE_PHN4313_n1026;
   wire FE_PHN4312_n2988;
   wire FE_PHN4311_n929;
   wire FE_PHN4310_n3977;
   wire FE_PHN4309_n954;
   wire FE_PHN4308_n4332;
   wire FE_PHN4307_n2754;
   wire FE_PHN4306_n3005;
   wire FE_PHN4305_n1038;
   wire FE_PHN4304_n2383;
   wire FE_PHN4303_n3060;
   wire FE_PHN4302_n2964;
   wire FE_PHN4301_n4244;
   wire FE_PHN4300_n4291;
   wire FE_PHN4299_n3046;
   wire FE_PHN4298_n3946;
   wire FE_PHN4297_n2967;
   wire FE_PHN4296_n4034;
   wire FE_PHN4295_n4103;
   wire FE_PHN4294_n3030;
   wire FE_PHN4293_n4286;
   wire FE_PHN4292_n3983;
   wire FE_PHN4291_n951;
   wire FE_PHN4290_n1902;
   wire FE_PHN4289_n1069;
   wire FE_PHN4288_n1896;
   wire FE_PHN4287_n3087;
   wire FE_PHN4286_n1025;
   wire FE_PHN4285_n992;
   wire FE_PHN4284_n2968;
   wire FE_PHN4283_n934;
   wire FE_PHN4282_n1064;
   wire FE_PHN4281_n3929;
   wire FE_PHN4280_n2433;
   wire FE_PHN4279_n4408;
   wire FE_PHN4278_n4361;
   wire FE_PHN4277_n4362;
   wire FE_PHN4276_n3071;
   wire FE_PHN4275_n4260;
   wire FE_PHN4274_n2703;
   wire FE_PHN4273_n4398;
   wire FE_PHN4272_n4220;
   wire FE_PHN4271_n1032;
   wire FE_PHN4270_n3132;
   wire FE_PHN4269_n2900;
   wire FE_PHN4268_n3117;
   wire FE_PHN4267_n846;
   wire FE_PHN4266_n887;
   wire FE_PHN4265_n2953;
   wire FE_PHN4264_n4307;
   wire FE_PHN4263_n4167;
   wire FE_PHN4262_n4023;
   wire FE_PHN4261_n852;
   wire FE_PHN4260_n3042;
   wire FE_PHN4259_n2985;
   wire FE_PHN4258_n3031;
   wire FE_PHN4257_ram_153__7_;
   wire FE_PHN4256_n4274;
   wire FE_PHN4255_n4010;
   wire FE_PHN4254_n3114;
   wire FE_PHN4253_n3966;
   wire FE_PHN4252_n3083;
   wire FE_PHN4251_n1873;
   wire FE_PHN4250_n1919;
   wire FE_PHN4249_n872;
   wire FE_PHN4248_n864;
   wire FE_PHN4247_n2932;
   wire FE_PHN4246_n1886;
   wire FE_PHN4245_n2969;
   wire FE_PHN4244_n3095;
   wire FE_PHN4243_n3223;
   wire FE_PHN4242_n947;
   wire FE_PHN4241_n978;
   wire FE_PHN4240_n3911;
   wire FE_PHN4239_n1911;
   wire FE_PHN4238_n2980;
   wire FE_PHN4237_n4290;
   wire FE_PHN4236_n1904;
   wire FE_PHN4235_n959;
   wire FE_PHN4234_n871;
   wire FE_PHN4233_n950;
   wire FE_PHN4232_n920;
   wire FE_PHN4231_n3110;
   wire FE_PHN4230_n1072;
   wire FE_PHN4229_n4327;
   wire FE_PHN4228_n945;
   wire FE_PHN4227_n3073;
   wire FE_PHN4226_n4363;
   wire FE_PHN4225_n989;
   wire FE_PHN4224_ram_238__0_;
   wire FE_PHN4223_n3123;
   wire FE_PHN4222_n4110;
   wire FE_PHN4221_n848;
   wire FE_PHN4220_n4289;
   wire FE_PHN4219_n3987;
   wire FE_PHN4218_n1864;
   wire FE_PHN4217_n842;
   wire FE_PHN4216_n1087;
   wire FE_PHN4215_n2958;
   wire FE_PHN4214_n3007;
   wire FE_PHN4213_n4379;
   wire FE_PHN4212_n1077;
   wire FE_PHN4211_n2952;
   wire FE_PHN4210_n3138;
   wire FE_PHN4209_n2408;
   wire FE_PHN4208_n927;
   wire FE_PHN4207_n4000;
   wire FE_PHN4206_n3089;
   wire FE_PHN4205_n2415;
   wire FE_PHN4204_n3043;
   wire FE_PHN4203_n4375;
   wire FE_PHN4202_n3070;
   wire FE_PHN4201_n4417;
   wire FE_PHN4200_n2982;
   wire FE_PHN4199_n4292;
   wire FE_PHN4198_n952;
   wire FE_PHN4197_n3972;
   wire FE_PHN4196_n3077;
   wire FE_PHN4195_n3012;
   wire FE_PHN4194_n893;
   wire FE_PHN4193_n1905;
   wire FE_PHN4192_n922;
   wire FE_PHN4191_n4001;
   wire FE_PHN4190_n4383;
   wire FE_PHN4189_n3111;
   wire FE_PHN4188_n4331;
   wire FE_PHN4187_n3027;
   wire FE_PHN4186_n1921;
   wire FE_PHN4185_ram_144__8_;
   wire FE_PHN4184_n3133;
   wire FE_PHN4183_n961;
   wire FE_PHN4182_n1040;
   wire FE_PHN4181_n4033;
   wire FE_PHN4180_n3959;
   wire FE_PHN4179_n3217;
   wire FE_PHN4178_n4410;
   wire FE_PHN4177_n3078;
   wire FE_PHN4176_n4007;
   wire FE_PHN4175_n2999;
   wire FE_PHN4174_n3000;
   wire FE_PHN4173_n3026;
   wire FE_PHN4172_ram_237__7_;
   wire FE_PHN4171_n4269;
   wire FE_PHN4170_n3103;
   wire FE_PHN4169_n3978;
   wire FE_PHN4168_n943;
   wire FE_PHN4167_n3023;
   wire FE_PHN4166_n4111;
   wire FE_PHN4165_n884;
   wire FE_PHN4164_n946;
   wire FE_PHN4163_n4225;
   wire FE_PHN4162_n3056;
   wire FE_PHN4161_ram_145__0_;
   wire FE_PHN4160_n4028;
   wire FE_PHN4159_n4413;
   wire FE_PHN4158_n3003;
   wire FE_PHN4157_n4022;
   wire FE_PHN4156_n4254;
   wire FE_PHN4155_ram_229__3_;
   wire FE_PHN4154_n901;
   wire FE_PHN4153_n4239;
   wire FE_PHN4152_n1088;
   wire FE_PHN4151_n3053;
   wire FE_PHN4150_n930;
   wire FE_PHN4149_n4031;
   wire FE_PHN4148_n1078;
   wire FE_PHN4147_n928;
   wire FE_PHN4146_n3979;
   wire FE_PHN4145_n4214;
   wire FE_PHN4144_n919;
   wire FE_PHN4143_n3943;
   wire FE_PHN4142_n4380;
   wire FE_PHN4141_n3115;
   wire FE_PHN4140_n4014;
   wire FE_PHN4139_n4009;
   wire FE_PHN4138_n2389;
   wire FE_PHN4137_n3982;
   wire FE_PHN4136_n4245;
   wire FE_PHN4135_n3265;
   wire FE_PHN4134_ram_145__1_;
   wire FE_PHN4133_n4008;
   wire FE_PHN4132_n4279;
   wire FE_PHN4131_n1008;
   wire FE_PHN4130_n1056;
   wire FE_PHN4129_ram_229__12_;
   wire FE_PHN4128_n865;
   wire FE_PHN4127_n3019;
   wire FE_PHN4126_n3009;
   wire FE_PHN4125_n4421;
   wire FE_PHN4124_n866;
   wire FE_PHN4123_ram_145__7_;
   wire FE_PHN4122_n4196;
   wire FE_PHN4121_n857;
   wire FE_PHN4120_n3081;
   wire FE_PHN4119_n4295;
   wire FE_PHN4118_n925;
   wire FE_PHN4117_n2374;
   wire FE_PHN4116_n4238;
   wire FE_PHN4115_n4146;
   wire FE_PHN4114_n4340;
   wire FE_PHN4113_n3915;
   wire FE_PHN4112_n2400;
   wire FE_PHN4111_n4387;
   wire FE_PHN4110_n3134;
   wire FE_PHN4109_n4138;
   wire FE_PHN4108_n3099;
   wire FE_PHN4107_n2994;
   wire FE_PHN4106_n3010;
   wire FE_PHN4105_ram_221__1_;
   wire FE_PHN4104_n958;
   wire FE_PHN4103_n876;
   wire FE_PHN4102_n2961;
   wire FE_PHN4101_n3102;
   wire FE_PHN4100_n4006;
   wire FE_PHN4099_n4371;
   wire FE_PHN4098_n3084;
   wire FE_PHN4097_n2991;
   wire FE_PHN4096_n3124;
   wire FE_PHN4095_n4356;
   wire FE_PHN4094_n4263;
   wire FE_PHN4093_n4389;
   wire FE_PHN4092_ram_17__14_;
   wire FE_PHN4091_n4367;
   wire FE_PHN4090_n2955;
   wire FE_PHN4089_n3948;
   wire FE_PHN4088_n3127;
   wire FE_PHN4087_ram_98__3_;
   wire FE_PHN4086_n4142;
   wire FE_PHN4085_n3048;
   wire FE_PHN4084_n2956;
   wire FE_PHN4083_n855;
   wire FE_PHN4082_n914;
   wire FE_PHN4081_n2973;
   wire FE_PHN4080_n3105;
   wire FE_PHN4079_n3092;
   wire FE_PHN4078_n3104;
   wire FE_PHN4077_n3107;
   wire FE_PHN4076_n4406;
   wire FE_PHN4075_n2962;
   wire FE_PHN4074_n4359;
   wire FE_PHN4073_n1005;
   wire FE_PHN4072_n3939;
   wire FE_PHN4071_n4003;
   wire FE_PHN4070_n4323;
   wire FE_PHN4069_n3260;
   wire FE_PHN4068_n3108;
   wire FE_PHN4067_n1045;
   wire FE_PHN4066_n4339;
   wire FE_PHN4065_n3128;
   wire FE_PHN4064_n4005;
   wire FE_PHN4063_n2979;
   wire FE_PHN4062_n2431;
   wire FE_PHN4061_n3118;
   wire FE_PHN4060_n4251;
   wire FE_PHN4059_n3001;
   wire FE_PHN4058_n2178;
   wire FE_PHN4057_n2977;
   wire FE_PHN4056_n4388;
   wire FE_PHN4055_n4405;
   wire FE_PHN4054_n984;
   wire FE_PHN4053_n1093;
   wire FE_PHN4052_n3116;
   wire FE_PHN4051_n1048;
   wire FE_PHN4050_n2981;
   wire FE_PHN4049_n3022;
   wire FE_PHN4048_n4372;
   wire FE_PHN4047_n2978;
   wire FE_PHN4046_n960;
   wire FE_PHN4045_n3112;
   wire FE_PHN4044_n3999;
   wire FE_PHN4043_n3930;
   wire FE_PHN4042_n3035;
   wire FE_PHN4041_n3100;
   wire FE_PHN4040_n4385;
   wire FE_PHN4039_n4384;
   wire FE_PHN4038_n856;
   wire FE_PHN4037_n1090;
   wire FE_PHN4036_n3914;
   wire FE_PHN4035_n4230;
   wire FE_PHN4034_n3937;
   wire FE_PHN4033_n918;
   wire FE_PHN4032_n4204;
   wire FE_PHN4031_n3947;
   wire FE_PHN4030_n2976;
   wire FE_PHN4029_n3032;
   wire FE_PHN4028_n3922;
   wire FE_PHN4027_n970;
   wire FE_PHN4026_ram_145__10_;
   wire FE_PHN4025_n3931;
   wire FE_PHN4024_n4324;
   wire FE_PHN4023_n4343;
   wire FE_PHN4022_n899;
   wire FE_PHN4021_n4399;
   wire FE_PHN4020_n3096;
   wire FE_PHN4019_n2966;
   wire FE_PHN4018_n3094;
   wire FE_PHN4017_n3926;
   wire FE_PHN4016_n3954;
   wire FE_PHN4015_n3993;
   wire FE_PHN4014_n4377;
   wire FE_PHN4013_n3998;
   wire FE_PHN4012_n4195;
   wire FE_PHN4011_n3125;
   wire FE_PHN4009_n2297;
   wire FE_PHN4008_n889;
   wire FE_PHN4007_n4416;
   wire FE_PHN4006_n961;
   wire FE_PHN4005_n898;
   wire FE_PHN4004_n3034;
   wire FE_PHN4003_n4032;
   wire FE_PHN4002_n1143;
   wire FE_PHN4001_n3004;
   wire FE_PHN4000_n4370;
   wire FE_PHN3999_n1042;
   wire FE_PHN3998_n896;
   wire FE_PHN3997_n892;
   wire FE_PHN3996_n2944;
   wire FE_PHN3995_n3135;
   wire FE_PHN3994_n4407;
   wire FE_PHN3993_n2954;
   wire FE_PHN3992_n2388;
   wire FE_PHN3991_n3130;
   wire FE_PHN3990_n870;
   wire FE_PHN3989_n976;
   wire FE_PHN3988_n4202;
   wire FE_PHN3987_n2963;
   wire FE_PHN3986_n3977;
   wire FE_PHN3985_n3257;
   wire FE_PHN3984_n1000;
   wire FE_PHN3983_n2722;
   wire FE_PHN3982_n3920;
   wire FE_PHN3981_n4403;
   wire FE_PHN3980_n2952;
   wire FE_PHN3979_n2933;
   wire FE_PHN3978_n2959;
   wire FE_PHN3977_n846;
   wire FE_PHN3976_n944;
   wire FE_PHN3975_n4289;
   wire FE_PHN3974_n1911;
   wire FE_PHN3973_n3114;
   wire FE_PHN3972_n2258;
   wire FE_PHN3971_n891;
   wire FE_PHN3970_n4361;
   wire FE_PHN3969_n2623;
   wire FE_PHN3968_n3255;
   wire FE_PHN3967_n3066;
   wire FE_PHN3966_n3962;
   wire FE_PHN3965_n4248;
   wire FE_PHN3964_n4401;
   wire FE_PHN3963_n3943;
   wire FE_PHN3962_n2621;
   wire FE_PHN3961_n4276;
   wire FE_PHN3960_n885;
   wire FE_PHN3959_n3076;
   wire FE_PHN3958_n3122;
   wire FE_PHN3957_n969;
   wire FE_PHN3956_n966;
   wire FE_PHN3955_n2605;
   wire FE_PHN3954_n3080;
   wire FE_PHN3953_n4268;
   wire FE_PHN3952_n4036;
   wire FE_PHN3951_n2946;
   wire FE_PHN3950_n4097;
   wire FE_PHN3949_n2564;
   wire FE_PHN3948_n4168;
   wire FE_PHN3947_n4273;
   wire FE_PHN3946_n3141;
   wire FE_PHN3945_n4420;
   wire FE_PHN3944_n3960;
   wire FE_PHN3943_n4387;
   wire FE_PHN3942_n3139;
   wire FE_PHN3941_n3953;
   wire FE_PHN3940_n968;
   wire FE_PHN3939_n2385;
   wire FE_PHN3938_n1110;
   wire FE_PHN3937_n4225;
   wire FE_PHN3936_n4333;
   wire FE_PHN3935_n1034;
   wire FE_PHN3934_n4185;
   wire FE_PHN3933_n4241;
   wire FE_PHN3932_n3050;
   wire FE_PHN3931_n876;
   wire FE_PHN3930_n4210;
   wire FE_PHN3929_n2945;
   wire FE_PHN3928_n3975;
   wire FE_PHN3927_n4046;
   wire FE_PHN3926_n886;
   wire FE_PHN3925_n4259;
   wire FE_PHN3924_ram_20__10_;
   wire FE_PHN3923_n4368;
   wire FE_PHN3922_n988;
   wire FE_PHN3921_n2419;
   wire FE_PHN3920_n2580;
   wire FE_PHN3919_n936;
   wire FE_PHN3918_n4187;
   wire FE_PHN3917_n2554;
   wire FE_PHN3916_n3219;
   wire FE_PHN3915_n4215;
   wire FE_PHN3914_n4410;
   wire FE_PHN3913_n4094;
   wire FE_PHN3912_n4373;
   wire FE_PHN3911_n3085;
   wire FE_PHN3910_n4242;
   wire FE_PHN3909_n951;
   wire FE_PHN3908_n3207;
   wire FE_PHN3907_n986;
   wire FE_PHN3906_n3067;
   wire FE_PHN3905_n3217;
   wire FE_PHN3904_n2965;
   wire FE_PHN3903_n851;
   wire FE_PHN3902_n4217;
   wire FE_PHN3901_n3011;
   wire FE_PHN3900_n2735;
   wire FE_PHN3899_n954;
   wire FE_PHN3898_n4183;
   wire FE_PHN3897_n3036;
   wire FE_PHN3896_n4338;
   wire FE_PHN3895_n2993;
   wire FE_PHN3894_n900;
   wire FE_PHN3893_n1918;
   wire FE_PHN3892_n945;
   wire FE_PHN3891_n3025;
   wire FE_PHN3890_n850;
   wire FE_PHN3889_n3079;
   wire FE_PHN3888_n3082;
   wire FE_PHN3887_n2383;
   wire FE_PHN3886_n3016;
   wire FE_PHN3885_n1024;
   wire FE_PHN3884_n895;
   wire FE_PHN3883_n2163;
   wire FE_PHN3882_n1023;
   wire FE_PHN3881_n3129;
   wire FE_PHN3880_n2995;
   wire FE_PHN3879_n3020;
   wire FE_PHN3878_n2900;
   wire FE_PHN3877_n999;
   wire FE_PHN3876_n920;
   wire FE_PHN3875_n1006;
   wire FE_PHN3874_n2408;
   wire FE_PHN3873_n3058;
   wire FE_PHN3872_n873;
   wire FE_PHN3871_n3951;
   wire FE_PHN3870_n904;
   wire FE_PHN3869_n1921;
   wire FE_PHN3868_n3075;
   wire FE_PHN3867_n2970;
   wire FE_PHN3866_n3074;
   wire FE_PHN3865_n902;
   wire FE_PHN3864_n1899;
   wire FE_PHN3863_n844;
   wire FE_PHN3862_ram_31__2_;
   wire FE_PHN3861_n905;
   wire FE_PHN3860_n3946;
   wire FE_PHN3859_n2967;
   wire FE_PHN3858_n2896;
   wire FE_PHN3857_n840;
   wire FE_PHN3856_n2753;
   wire FE_PHN3855_n4229;
   wire FE_PHN3854_ram_238__0_;
   wire FE_PHN3853_n1874;
   wire FE_PHN3852_n2916;
   wire FE_PHN3851_n3119;
   wire FE_PHN3850_n3109;
   wire FE_PHN3849_n3054;
   wire FE_PHN3848_n4397;
   wire FE_PHN3847_n934;
   wire FE_PHN3846_n913;
   wire FE_PHN3845_n952;
   wire FE_PHN3844_n4227;
   wire FE_PHN3843_n2986;
   wire FE_PHN3842_n1079;
   wire FE_PHN3841_n3060;
   wire FE_PHN3840_n1922;
   wire FE_PHN3839_n2384;
   wire FE_PHN3838_n3090;
   wire FE_PHN3837_n3029;
   wire FE_PHN3836_n906;
   wire FE_PHN3835_n3262;
   wire FE_PHN3834_n4209;
   wire FE_PHN3833_n1880;
   wire FE_PHN3832_n949;
   wire FE_PHN3831_n1906;
   wire FE_PHN3830_n3015;
   wire FE_PHN3829_n1021;
   wire FE_PHN3828_n4400;
   wire FE_PHN3827_n959;
   wire FE_PHN3826_n2943;
   wire FE_PHN3825_n4283;
   wire FE_PHN3824_n4265;
   wire FE_PHN3823_n4134;
   wire FE_PHN3822_n4366;
   wire FE_PHN3821_n2574;
   wire FE_PHN3820_n1030;
   wire FE_PHN3819_n3994;
   wire FE_PHN3818_n4111;
   wire FE_PHN3817_n1916;
   wire FE_PHN3816_n1037;
   wire FE_PHN3815_n3963;
   wire FE_PHN3814_n1896;
   wire FE_PHN3813_n888;
   wire FE_PHN3812_n3210;
   wire FE_PHN3811_n841;
   wire FE_PHN3810_n2962;
   wire FE_PHN3809_n2437;
   wire FE_PHN3808_n4291;
   wire FE_PHN3807_n3062;
   wire FE_PHN3806_n845;
   wire FE_PHN3805_n2990;
   wire FE_PHN3804_n4037;
   wire FE_PHN3803_n962;
   wire FE_PHN3802_n1038;
   wire FE_PHN3801_n3916;
   wire FE_PHN3800_n4231;
   wire FE_PHN3799_n3942;
   wire FE_PHN3798_n3968;
   wire FE_PHN3797_n4362;
   wire FE_PHN3796_n1077;
   wire FE_PHN3795_n3940;
   wire FE_PHN3794_n4277;
   wire FE_PHN3793_n3046;
   wire FE_PHN3792_n1919;
   wire FE_PHN3791_n1002;
   wire FE_PHN3790_n910;
   wire FE_PHN3789_n965;
   wire FE_PHN3788_n3956;
   wire FE_PHN3787_n3019;
   wire FE_PHN3786_n4158;
   wire FE_PHN3785_n2898;
   wire FE_PHN3784_n853;
   wire FE_PHN3783_n943;
   wire FE_PHN3782_n2415;
   wire FE_PHN3781_n4076;
   wire FE_PHN3780_n3955;
   wire FE_PHN3779_n3026;
   wire FE_PHN3778_n2957;
   wire FE_PHN3777_n2732;
   wire FE_PHN3776_n843;
   wire FE_PHN3775_n3965;
   wire FE_PHN3774_n3932;
   wire FE_PHN3773_n4207;
   wire FE_PHN3772_n3110;
   wire FE_PHN3771_n880;
   wire FE_PHN3770_n4409;
   wire FE_PHN3769_n2598;
   wire FE_PHN3768_n3077;
   wire FE_PHN3767_n947;
   wire FE_PHN3766_n2897;
   wire FE_PHN3765_n2975;
   wire FE_PHN3764_n1902;
   wire FE_PHN3763_n1873;
   wire FE_PHN3762_n2958;
   wire FE_PHN3761_n3126;
   wire FE_PHN3760_n1864;
   wire FE_PHN3759_n3028;
   wire FE_PHN3758_n3042;
   wire FE_PHN3757_n919;
   wire FE_PHN3756_n2969;
   wire FE_PHN3755_n4172;
   wire FE_PHN3754_n2922;
   wire FE_PHN3753_n4218;
   wire FE_PHN3752_n1905;
   wire FE_PHN3751_n3989;
   wire FE_PHN3750_n4035;
   wire FE_PHN3749_n3005;
   wire FE_PHN3748_n4062;
   wire FE_PHN3747_n4222;
   wire FE_PHN3746_n3040;
   wire FE_PHN3745_n1020;
   wire FE_PHN3744_n928;
   wire FE_PHN3743_n3069;
   wire FE_PHN3742_n4027;
   wire FE_PHN3741_n3980;
   wire FE_PHN3740_n3012;
   wire FE_PHN3739_n3084;
   wire FE_PHN3738_n3000;
   wire FE_PHN3737_n2991;
   wire FE_PHN3736_n2997;
   wire FE_PHN3735_n4255;
   wire FE_PHN3734_n978;
   wire FE_PHN3733_n2982;
   wire FE_PHN3732_n872;
   wire FE_PHN3731_n4236;
   wire FE_PHN3730_n3007;
   wire FE_PHN3729_n2961;
   wire FE_PHN3728_n4395;
   wire FE_PHN3727_n1029;
   wire FE_PHN3726_n903;
   wire FE_PHN3725_n1072;
   wire FE_PHN3724_n3926;
   wire FE_PHN3723_n972;
   wire FE_PHN3722_ram_154__5_;
   wire FE_PHN3721_n4049;
   wire FE_PHN3720_n3966;
   wire FE_PHN3719_n3083;
   wire FE_PHN3718_n2928;
   wire FE_PHN3717_n1920;
   wire FE_PHN3716_n1904;
   wire FE_PHN3715_n1106;
   wire FE_PHN3714_n4175;
   wire FE_PHN3713_n4103;
   wire FE_PHN3712_n3136;
   wire FE_PHN3711_n991;
   wire FE_PHN3710_n3921;
   wire FE_PHN3709_n925;
   wire FE_PHN3708_n941;
   wire FE_PHN3707_n2955;
   wire FE_PHN3706_n2983;
   wire FE_PHN3705_n4232;
   wire FE_PHN3704_n3964;
   wire FE_PHN3703_n3070;
   wire FE_PHN3702_n2733;
   wire FE_PHN3701_n2405;
   wire FE_PHN3700_n2599;
   wire FE_PHN3699_n4261;
   wire FE_PHN3698_n4170;
   wire FE_PHN3697_n2968;
   wire FE_PHN3696_n887;
   wire FE_PHN3695_n1088;
   wire FE_PHN3694_n3241;
   wire FE_PHN3693_n3984;
   wire FE_PHN3692_n2430;
   wire FE_PHN3691_ram_214__13_;
   wire FE_PHN3690_ram_153__11_;
   wire FE_PHN3689_n4148;
   wire FE_PHN3688_n3265;
   wire FE_PHN3687_n4269;
   wire FE_PHN3686_n1051;
   wire FE_PHN3685_n1068;
   wire FE_PHN3684_n871;
   wire FE_PHN3683_n4308;
   wire FE_PHN3682_n957;
   wire FE_PHN3681_n3918;
   wire FE_PHN3680_n4016;
   wire FE_PHN3679_n3072;
   wire FE_PHN3678_n4181;
   wire FE_PHN3677_n2960;
   wire FE_PHN3676_n1082;
   wire FE_PHN3675_n4204;
   wire FE_PHN3674_n4290;
   wire FE_PHN3673_n1069;
   wire FE_PHN3672_n1027;
   wire FE_PHN3671_n3006;
   wire FE_PHN3670_n950;
   wire FE_PHN3669_n3013;
   wire FE_PHN3668_n852;
   wire FE_PHN3667_n4365;
   wire FE_PHN3666_n2998;
   wire FE_PHN3665_n4178;
   wire FE_PHN3664_n842;
   wire FE_PHN3663_n2953;
   wire FE_PHN3662_n3978;
   wire FE_PHN3661_n4007;
   wire FE_PHN3660_n839;
   wire FE_PHN3659_n1040;
   wire FE_PHN3658_n1087;
   wire FE_PHN3657_n4240;
   wire FE_PHN3656_n3088;
   wire FE_PHN3655_n4025;
   wire FE_PHN3654_n863;
   wire FE_PHN3653_n2989;
   wire FE_PHN3652_n4271;
   wire FE_PHN3651_n2971;
   wire FE_PHN3650_n4000;
   wire FE_PHN3649_n3128;
   wire FE_PHN3648_n3056;
   wire FE_PHN3647_n992;
   wire FE_PHN3646_n2985;
   wire FE_PHN3645_n4329;
   wire FE_PHN3644_n4213;
   wire FE_PHN3643_n4415;
   wire FE_PHN3642_n3086;
   wire FE_PHN3641_ram_144__8_;
   wire FE_PHN3640_n3023;
   wire FE_PHN3639_n2420;
   wire FE_PHN3638_n4279;
   wire FE_PHN3637_n3133;
   wire FE_PHN3636_n847;
   wire FE_PHN3635_n2399;
   wire FE_PHN3634_n4009;
   wire FE_PHN3633_n922;
   wire FE_PHN3632_n4267;
   wire FE_PHN3631_n3055;
   wire FE_PHN3630_n4219;
   wire FE_PHN3629_n3112;
   wire FE_PHN3628_n4274;
   wire FE_PHN3627_n4245;
   wire FE_PHN3626_n1206;
   wire FE_PHN3625_n1025;
   wire FE_PHN3624_n4239;
   wire FE_PHN3623_n1018;
   wire FE_PHN3622_n2754;
   wire FE_PHN3621_n4367;
   wire FE_PHN3620_n4392;
   wire FE_PHN3619_n909;
   wire FE_PHN3618_n3073;
   wire FE_PHN3617_n2891;
   wire FE_PHN3616_n3098;
   wire FE_PHN3615_n4316;
   wire FE_PHN3614_n3003;
   wire FE_PHN3613_n2262;
   wire FE_PHN3612_n3024;
   wire FE_PHN3611_n4382;
   wire FE_PHN3610_n4334;
   wire FE_PHN3609_n3117;
   wire FE_PHN3608_n2996;
   wire FE_PHN3607_n2432;
   wire FE_PHN3606_n4116;
   wire FE_PHN3605_n2403;
   wire FE_PHN3604_n4171;
   wire FE_PHN3603_n1009;
   wire FE_PHN3602_n2727;
   wire FE_PHN3601_n3914;
   wire FE_PHN3600_n2935;
   wire FE_PHN3599_n4238;
   wire FE_PHN3598_n4299;
   wire FE_PHN3597_n4404;
   wire FE_PHN3596_n4413;
   wire FE_PHN3595_n911;
   wire FE_PHN3594_n4228;
   wire FE_PHN3593_ram_145__7_;
   wire FE_PHN3592_n3982;
   wire FE_PHN3591_n3950;
   wire FE_PHN3590_n3102;
   wire FE_PHN3589_n4188;
   wire FE_PHN3588_n3134;
   wire FE_PHN3587_n3971;
   wire FE_PHN3586_n3263;
   wire FE_PHN3585_n964;
   wire FE_PHN3584_n2994;
   wire FE_PHN3583_n3027;
   wire FE_PHN3582_n4371;
   wire FE_PHN3581_n4359;
   wire FE_PHN3580_n2951;
   wire FE_PHN3579_n901;
   wire FE_PHN3578_n3992;
   wire FE_PHN3577_n2978;
   wire FE_PHN3576_n3091;
   wire FE_PHN3575_n3044;
   wire FE_PHN3574_n4294;
   wire FE_PHN3573_n935;
   wire FE_PHN3572_n2992;
   wire FE_PHN3571_ram_133__9_;
   wire FE_PHN3570_n890;
   wire FE_PHN3569_n998;
   wire FE_PHN3568_n997;
   wire FE_PHN3567_n2431;
   wire FE_PHN3566_n927;
   wire FE_PHN3565_n3970;
   wire FE_PHN3564_n3917;
   wire FE_PHN3563_n1066;
   wire FE_PHN3562_n3095;
   wire FE_PHN3561_n3911;
   wire FE_PHN3560_n989;
   wire FE_PHN3559_n3009;
   wire FE_PHN3558_n3132;
   wire FE_PHN3557_n874;
   wire FE_PHN3556_n2987;
   wire FE_PHN3555_n849;
   wire FE_PHN3554_n2927;
   wire FE_PHN3553_n3137;
   wire FE_PHN3552_n2389;
   wire FE_PHN3551_n1870;
   wire FE_PHN3550_n4226;
   wire FE_PHN3549_n3018;
   wire FE_PHN3548_n4364;
   wire FE_PHN3547_n3140;
   wire FE_PHN3546_n984;
   wire FE_PHN3545_n1048;
   wire FE_PHN3544_n3010;
   wire FE_PHN3543_n4169;
   wire FE_PHN3542_n2932;
   wire FE_PHN3541_n4179;
   wire FE_PHN3540_n4212;
   wire FE_PHN3539_n4295;
   wire FE_PHN3538_n4211;
   wire FE_PHN3537_n4340;
   wire FE_PHN3536_n4414;
   wire FE_PHN3535_n938;
   wire FE_PHN3534_n3913;
   wire FE_PHN3533_n897;
   wire FE_PHN3532_n3052;
   wire FE_PHN3531_ram_229__12_;
   wire FE_PHN3530_n2923;
   wire FE_PHN3529_n857;
   wire FE_PHN3528_n878;
   wire FE_PHN3527_n975;
   wire FE_PHN3526_n3972;
   wire FE_PHN3525_n1056;
   wire FE_PHN3524_n3958;
   wire FE_PHN3523_n4356;
   wire FE_PHN3522_n894;
   wire FE_PHN3521_n4262;
   wire FE_PHN3520_n3002;
   wire FE_PHN3519_ram_229__3_;
   wire FE_PHN3518_n2980;
   wire FE_PHN3517_n3952;
   wire FE_PHN3516_n4034;
   wire FE_PHN3515_n3258;
   wire FE_PHN3514_n4369;
   wire FE_PHN3513_n4220;
   wire FE_PHN3512_n4292;
   wire FE_PHN3511_n982;
   wire FE_PHN3510_n4022;
   wire FE_PHN3509_n929;
   wire FE_PHN3508_n4233;
   wire FE_PHN3507_n2400;
   wire FE_PHN3506_n971;
   wire FE_PHN3505_n4412;
   wire FE_PHN3504_n914;
   wire FE_PHN3503_n4323;
   wire FE_PHN3502_ram_145__1_;
   wire FE_PHN3501_n3923;
   wire FE_PHN3500_n3948;
   wire FE_PHN3499_n4087;
   wire FE_PHN3498_n3945;
   wire FE_PHN3497_n2413;
   wire FE_PHN3496_n2703;
   wire FE_PHN3495_n4284;
   wire FE_PHN3494_n893;
   wire FE_PHN3493_n4138;
   wire FE_PHN3492_n882;
   wire FE_PHN3491_n4350;
   wire FE_PHN3490_n2964;
   wire FE_PHN3489_n3065;
   wire FE_PHN3488_ram_221__1_;
   wire FE_PHN3487_n899;
   wire FE_PHN3486_n2374;
   wire FE_PHN3485_n3089;
   wire FE_PHN3484_n2600;
   wire FE_PHN3483_n4331;
   wire FE_PHN3482_n2906;
   wire FE_PHN3481_n3078;
   wire FE_PHN3480_n4266;
   wire FE_PHN3479_n4418;
   wire FE_PHN3478_n2981;
   wire FE_PHN3477_n3910;
   wire FE_PHN3476_n1078;
   wire FE_PHN3475_n2976;
   wire FE_PHN3474_n4244;
   wire FE_PHN3473_n4419;
   wire FE_PHN3472_n3118;
   wire FE_PHN3471_n948;
   wire FE_PHN3470_n2999;
   wire FE_PHN3469_n1872;
   wire FE_PHN3468_n3123;
   wire FE_PHN3467_n4110;
   wire FE_PHN3466_n3976;
   wire FE_PHN3465_n4142;
   wire FE_PHN3464_n877;
   wire FE_PHN3463_n933;
   wire FE_PHN3462_n3930;
   wire FE_PHN3461_n3096;
   wire FE_PHN3460_n4285;
   wire FE_PHN3459_n4278;
   wire FE_PHN3458_n4327;
   wire FE_PHN3457_n4396;
   wire FE_PHN3456_n4378;
   wire FE_PHN3455_n4394;
   wire FE_PHN3454_n1017;
   wire FE_PHN3453_n3131;
   wire FE_PHN3452_n2131;
   wire FE_PHN3451_ram_17__14_;
   wire FE_PHN3450_n3944;
   wire FE_PHN3449_n3924;
   wire FE_PHN3448_n2974;
   wire FE_PHN3447_n4399;
   wire FE_PHN3446_n4023;
   wire FE_PHN3445_n2972;
   wire FE_PHN3444_n2926;
   wire FE_PHN3443_n4026;
   wire FE_PHN3442_n3979;
   wire FE_PHN3441_n861;
   wire FE_PHN3440_n994;
   wire FE_PHN3439_n946;
   wire FE_PHN3438_n3127;
   wire FE_PHN3437_n1886;
   wire FE_PHN3436_n958;
   wire FE_PHN3435_n2178;
   wire FE_PHN3434_n3103;
   wire FE_PHN3433_n3008;
   wire FE_PHN3432_n917;
   wire FE_PHN3431_n1022;
   wire FE_PHN3430_n2956;
   wire FE_PHN3429_n3936;
   wire FE_PHN3428_n4260;
   wire FE_PHN3427_n4360;
   wire FE_PHN3426_n2886;
   wire FE_PHN3425_n4375;
   wire FE_PHN3424_n2918;
   wire FE_PHN3423_n2984;
   wire FE_PHN3422_n3111;
   wire FE_PHN3421_n3093;
   wire FE_PHN3420_n1016;
   wire FE_PHN3419_n3049;
   wire FE_PHN3418_n3048;
   wire FE_PHN3417_n4363;
   wire FE_PHN3416_n3120;
   wire FE_PHN3415_n4174;
   wire FE_PHN3414_n4199;
   wire FE_PHN3413_n4146;
   wire FE_PHN3412_n4005;
   wire FE_PHN3411_n3032;
   wire FE_PHN3410_n3223;
   wire FE_PHN3409_n993;
   wire FE_PHN3408_n1093;
   wire FE_PHN3407_n3071;
   wire FE_PHN3406_n4031;
   wire FE_PHN3405_n1045;
   wire FE_PHN3404_n2904;
   wire FE_PHN3403_n3915;
   wire FE_PHN3402_n4029;
   wire FE_PHN3401_n930;
   wire FE_PHN3400_n2433;
   wire FE_PHN3399_n4206;
   wire FE_PHN3398_n3022;
   wire FE_PHN3397_n4017;
   wire FE_PHN3396_n4196;
   wire FE_PHN3395_n866;
   wire FE_PHN3394_n4417;
   wire FE_PHN3393_n1008;
   wire FE_PHN3392_n4030;
   wire FE_PHN3391_n974;
   wire FE_PHN3390_n3212;
   wire FE_PHN3389_ram_237__7_;
   wire FE_PHN3388_n3260;
   wire FE_PHN3387_n2920;
   wire FE_PHN3386_n3108;
   wire FE_PHN3385_n4421;
   wire FE_PHN3384_n4372;
   wire FE_PHN3383_n4201;
   wire FE_PHN3382_n4164;
   wire FE_PHN3381_n3038;
   wire FE_PHN3380_n4300;
   wire FE_PHN3379_n2950;
   wire FE_PHN3378_n4166;
   wire FE_PHN3377_n4408;
   wire FE_PHN3376_n848;
   wire FE_PHN3375_n1014;
   wire FE_PHN3374_ram_158__11_;
   wire FE_PHN3373_ram_153__7_;
   wire FE_PHN3372_n3116;
   wire FE_PHN3371_n2127;
   wire FE_PHN3370_n4281;
   wire FE_PHN3369_n4235;
   wire FE_PHN3368_n1090;
   wire FE_PHN3367_n2977;
   wire FE_PHN3366_n838;
   wire FE_PHN3365_n960;
   wire FE_PHN3364_n4270;
   wire FE_PHN3363_n918;
   wire FE_PHN3362_n3031;
   wire FE_PHN3361_n4028;
   wire FE_PHN3360_n4254;
   wire FE_PHN3359_n1032;
   wire FE_PHN3358_ram_145__0_;
   wire FE_PHN3357_n4251;
   wire FE_PHN3356_n3922;
   wire FE_PHN3355_n4405;
   wire FE_PHN3354_n4355;
   wire FE_PHN3353_n4214;
   wire FE_PHN3352_n3959;
   wire FE_PHN3351_n3104;
   wire FE_PHN3350_n3053;
   wire FE_PHN3349_n4307;
   wire FE_PHN3348_n2930;
   wire FE_PHN3347_ram_98__3_;
   wire FE_PHN3346_n3947;
   wire FE_PHN3345_n856;
   wire FE_PHN3344_n3138;
   wire FE_PHN3343_n2979;
   wire FE_PHN3342_n3983;
   wire FE_PHN3341_n3927;
   wire FE_PHN3340_n1005;
   wire FE_PHN3339_n3124;
   wire FE_PHN3338_n3001;
   wire FE_PHN3337_n3035;
   wire FE_PHN3336_n3115;
   wire FE_PHN3335_n869;
   wire FE_PHN3334_n3064;
   wire FE_PHN3333_n2888;
   wire FE_PHN3332_n4311;
   wire FE_PHN3331_n4398;
   wire FE_PHN3330_n1062;
   wire FE_PHN3329_n3081;
   wire FE_PHN3328_n3099;
   wire FE_PHN3327_n4001;
   wire FE_PHN3326_n4406;
   wire FE_PHN3325_n4393;
   wire FE_PHN3324_n3094;
   wire FE_PHN3323_n970;
   wire FE_PHN3322_n4342;
   wire FE_PHN3321_n4230;
   wire FE_PHN3320_n2973;
   wire FE_PHN3319_n4358;
   wire FE_PHN3318_n884;
   wire FE_PHN3317_n4194;
   wire FE_PHN3316_n4411;
   wire FE_PHN3315_n2988;
   wire FE_PHN3314_n3988;
   wire FE_PHN3313_n3937;
   wire FE_PHN3312_n3092;
   wire FE_PHN3311_n858;
   wire FE_PHN3310_n3043;
   wire FE_PHN3309_n881;
   wire FE_PHN3308_n865;
   wire FE_PHN3307_n3961;
   wire FE_PHN3306_n4286;
   wire FE_PHN3305_n879;
   wire FE_PHN3304_n4377;
   wire FE_PHN3303_n3939;
   wire FE_PHN3302_n4263;
   wire FE_PHN3301_n3014;
   wire FE_PHN3300_n3105;
   wire FE_PHN3299_n4180;
   wire FE_PHN3298_n2421;
   wire FE_PHN3297_n4402;
   wire FE_PHN3296_n4380;
   wire FE_PHN3295_n854;
   wire FE_PHN3294_n4003;
   wire FE_PHN3293_n3919;
   wire FE_PHN3292_n4386;
   wire FE_PHN3291_n3934;
   wire FE_PHN3290_n3063;
   wire FE_PHN3289_n3969;
   wire FE_PHN3288_n4167;
   wire FE_PHN3287_n4374;
   wire FE_PHN3286_ram_145__10_;
   wire FE_PHN3285_n1046;
   wire FE_PHN3284_n4014;
   wire FE_PHN3283_n2396;
   wire FE_PHN3282_n3087;
   wire FE_PHN3281_n1074;
   wire FE_PHN3280_n4379;
   wire FE_PHN3279_n864;
   wire FE_PHN3278_n3954;
   wire FE_PHN3277_n4195;
   wire FE_PHN3276_n855;
   wire FE_PHN3275_n3107;
   wire FE_PHN3274_n3998;
   wire FE_PHN3273_n3993;
   wire FE_PHN3272_n2966;
   wire FE_PHN3271_n3974;
   wire FE_PHN3270_n4123;
   wire FE_PHN3269_n1013;
   wire FE_PHN3268_n4243;
   wire FE_PHN3267_n4388;
   wire FE_PHN3266_n2158;
   wire FE_PHN3265_n2910;
   wire FE_PHN3264_n3100;
   wire FE_PHN3263_n4033;
   wire FE_PHN3262_n2141;
   wire FE_PHN3261_n4343;
   wire FE_PHN3260_n4332;
   wire FE_PHN3259_n3996;
   wire FE_PHN3258_n4391;
   wire FE_PHN3257_n2936;
   wire FE_PHN3256_n4339;
   wire FE_PHN3255_n4389;
   wire FE_PHN3254_n4384;
   wire FE_PHN3253_n2934;
   wire FE_PHN3252_n4383;
   wire FE_PHN3251_n4010;
   wire FE_PHN3250_n1064;
   wire FE_PHN3249_n4203;
   wire FE_PHN3248_n4021;
   wire FE_PHN3247_n3125;
   wire FE_PHN3246_n2391;
   wire FE_PHN3245_n3030;
   wire FE_PHN3244_n3929;
   wire FE_PHN3243_n3985;
   wire FE_PHN3242_n1026;
   wire FE_PHN3241_n4006;
   wire FE_PHN3240_n3999;
   wire FE_PHN3239_n4252;
   wire FE_PHN3238_n3987;
   wire FE_PHN3237_n4008;
   wire FE_PHN3236_n4385;
   wire FE_PHN3235_n4015;
   wire FE_PHN3234_n3931;
   wire FE_PHN3233_n4324;
   wire FE_PHN3230_n1489;
   wire FE_PHN3229_n3451;
   wire FE_PHN3228_n1773;
   wire FE_PHN3227_n649;
   wire FE_PHN3226_n2005;
   wire FE_PHN3225_n809;
   wire FE_PHN3224_n713;
   wire FE_PHN3223_n1197;
   wire FE_PHN3222_n1099;
   wire FE_PHN3221_n2104;
   wire FE_PHN3220_n1536;
   wire FE_PHN3219_n3461;
   wire FE_PHN3218_n625;
   wire FE_PHN3217_n3427;
   wire FE_PHN3216_n1425;
   wire FE_PHN3215_n1132;
   wire FE_PHN3214_n1815;
   wire FE_PHN3213_n3152;
   wire FE_PHN3212_n3520;
   wire FE_PHN3211_n1422;
   wire FE_PHN3210_n4162;
   wire FE_PHN3209_n768;
   wire FE_PHN3208_n1688;
   wire FE_PHN3207_n3284;
   wire FE_PHN3206_n3848;
   wire FE_PHN3205_n3592;
   wire FE_PHN3204_n590;
   wire FE_PHN3203_n3469;
   wire FE_PHN3202_n4541;
   wire FE_PHN3201_n1962;
   wire FE_PHN3200_n2360;
   wire FE_PHN3199_n2355;
   wire FE_PHN3198_n1324;
   wire FE_PHN3197_n3688;
   wire FE_PHN3196_n1401;
   wire FE_PHN3195_n706;
   wire FE_PHN3194_n1328;
   wire FE_PHN3193_n2012;
   wire FE_PHN3192_n3846;
   wire FE_PHN3191_n1511;
   wire FE_PHN3190_n1978;
   wire FE_PHN3189_n749;
   wire FE_PHN3188_n1780;
   wire FE_PHN3187_n1993;
   wire FE_PHN3186_n3481;
   wire FE_PHN3185_n1799;
   wire FE_PHN3184_n1601;
   wire FE_PHN3183_n3541;
   wire FE_PHN3182_n1382;
   wire FE_PHN3181_n2870;
   wire FE_PHN3180_n592;
   wire FE_PHN3179_n717;
   wire FE_PHN3178_n1825;
   wire FE_PHN3177_n4353;
   wire FE_PHN3176_n832;
   wire FE_PHN3175_n2505;
   wire FE_PHN3174_n3843;
   wire FE_PHN3173_n3519;
   wire FE_PHN3172_n3388;
   wire FE_PHN3171_n3769;
   wire FE_PHN3170_n1279;
   wire FE_PHN3169_n3483;
   wire FE_PHN3168_n3471;
   wire FE_PHN3167_n3280;
   wire FE_PHN3166_n2511;
   wire FE_PHN3165_n2196;
   wire FE_PHN3164_n594;
   wire FE_PHN3163_n2549;
   wire FE_PHN3162_n4540;
   wire FE_PHN3161_n2227;
   wire FE_PHN3160_n1277;
   wire FE_PHN3159_n1449;
   wire FE_PHN3158_n801;
   wire FE_PHN3157_n4096;
   wire FE_PHN3156_n1405;
   wire FE_PHN3155_n3891;
   wire FE_PHN3154_n1772;
   wire FE_PHN3153_n1699;
   wire FE_PHN3152_n812;
   wire FE_PHN3151_n1236;
   wire FE_PHN3150_n651;
   wire FE_PHN3149_n770;
   wire FE_PHN3148_n1254;
   wire FE_PHN3147_n2949;
   wire FE_PHN3146_n3640;
   wire FE_PHN3145_n1118;
   wire FE_PHN3144_n1676;
   wire FE_PHN3143_n1937;
   wire FE_PHN3142_n1901;
   wire FE_PHN3141_n1804;
   wire FE_PHN3140_n1529;
   wire FE_PHN3139_n3243;
   wire FE_PHN3138_n1269;
   wire FE_PHN3137_n758;
   wire FE_PHN3136_n2358;
   wire FE_PHN3135_n688;
   wire FE_PHN3134_n3797;
   wire FE_PHN3133_n715;
   wire FE_PHN3132_n1354;
   wire FE_PHN3131_n2446;
   wire FE_PHN3130_n2223;
   wire FE_PHN3129_n1203;
   wire FE_PHN3128_n2700;
   wire FE_PHN3127_n1043;
   wire FE_PHN3126_n1737;
   wire FE_PHN3125_n1593;
   wire FE_PHN3124_n4557;
   wire FE_PHN3123_n3777;
   wire FE_PHN3122_n3220;
   wire FE_PHN3121_n4173;
   wire FE_PHN3120_n2613;
   wire FE_PHN3119_n3784;
   wire FE_PHN3118_n2868;
   wire FE_PHN3117_n1714;
   wire FE_PHN3116_n3143;
   wire FE_PHN3115_n3697;
   wire FE_PHN3114_n781;
   wire FE_PHN3113_n1452;
   wire FE_PHN3112_n2773;
   wire FE_PHN3111_n1212;
   wire FE_PHN3110_n2788;
   wire FE_PHN3109_n1355;
   wire FE_PHN3108_n3535;
   wire FE_PHN3107_n3191;
   wire FE_PHN3106_n1358;
   wire FE_PHN3105_n1741;
   wire FE_PHN3104_n2802;
   wire FE_PHN3103_n1829;
   wire FE_PHN3102_n2052;
   wire FE_PHN3101_n2692;
   wire FE_PHN3100_n2112;
   wire FE_PHN3099_n2636;
   wire FE_PHN3098_n1104;
   wire FE_PHN3097_n1850;
   wire FE_PHN3096_n1470;
   wire FE_PHN3095_n3467;
   wire FE_PHN3094_n3453;
   wire FE_PHN3093_n1150;
   wire FE_PHN3092_n3854;
   wire FE_PHN3091_n2499;
   wire FE_PHN3090_n3328;
   wire FE_PHN3089_n3332;
   wire FE_PHN3088_n907;
   wire FE_PHN3087_n1935;
   wire FE_PHN3086_n4043;
   wire FE_PHN3085_n1731;
   wire FE_PHN3084_n641;
   wire FE_PHN3083_n1166;
   wire FE_PHN3082_n3459;
   wire FE_PHN3081_n2815;
   wire FE_PHN3080_n1163;
   wire FE_PHN3079_n4143;
   wire FE_PHN3078_n1426;
   wire FE_PHN3077_n1652;
   wire FE_PHN3076_n1461;
   wire FE_PHN3075_n1681;
   wire FE_PHN3074_ram_143__10_;
   wire FE_PHN3073_ram_52__15_;
   wire FE_PHN3072_n3319;
   wire FE_PHN3071_n2041;
   wire FE_PHN3070_n1229;
   wire FE_PHN3069_n2214;
   wire FE_PHN3068_n4642;
   wire FE_PHN3067_n1484;
   wire FE_PHN3066_n811;
   wire FE_PHN3065_n1101;
   wire FE_PHN3064_n1161;
   wire FE_PHN3063_n1349;
   wire FE_PHN3062_n2304;
   wire FE_PHN3061_n620;
   wire FE_PHN3060_n1134;
   wire FE_PHN3059_n1615;
   wire FE_PHN3058_n1413;
   wire FE_PHN3057_n3908;
   wire FE_PHN3056_n3487;
   wire FE_PHN3055_n1784;
   wire FE_PHN3054_n1491;
   wire FE_PHN3053_n2464;
   wire FE_PHN3052_n596;
   wire FE_PHN3051_n3634;
   wire FE_PHN3050_n1111;
   wire FE_PHN3049_n1376;
   wire FE_PHN3048_n1543;
   wire FE_PHN3047_n1600;
   wire FE_PHN3046_n2053;
   wire FE_PHN3045_n1574;
   wire FE_PHN3044_n4662;
   wire FE_PHN3043_n631;
   wire FE_PHN3042_n1618;
   wire FE_PHN3041_n1419;
   wire FE_PHN3040_n3778;
   wire FE_PHN3039_n1787;
   wire FE_PHN3038_n1726;
   wire FE_PHN3037_n585;
   wire FE_PHN3036_n721;
   wire FE_PHN3035_n2746;
   wire FE_PHN3034_n828;
   wire FE_PHN3033_n1757;
   wire FE_PHN3032_n1259;
   wire FE_PHN3031_n4510;
   wire FE_PHN3030_n3462;
   wire FE_PHN3029_n1613;
   wire FE_PHN3028_n1301;
   wire FE_PHN3027_n729;
   wire FE_PHN3026_n2055;
   wire FE_PHN3025_n3261;
   wire FE_PHN3024_n2885;
   wire FE_PHN3023_n1859;
   wire FE_PHN3022_n1941;
   wire FE_PHN3021_n4670;
   wire FE_PHN3020_n2098;
   wire FE_PHN3019_n1856;
   wire FE_PHN3018_n2665;
   wire FE_PHN3017_n1579;
   wire FE_PHN3016_n2240;
   wire FE_PHN3015_n2845;
   wire FE_PHN3014_n1417;
   wire FE_PHN3013_ram_244__10_;
   wire FE_PHN3012_n2031;
   wire FE_PHN3011_n616;
   wire FE_PHN3010_n1361;
   wire FE_PHN3009_n1540;
   wire FE_PHN3008_n3443;
   wire FE_PHN3007_n1289;
   wire FE_PHN3006_n2051;
   wire FE_PHN3005_n1451;
   wire FE_PHN3004_n4542;
   wire FE_PHN3003_n3466;
   wire FE_PHN3002_n1969;
   wire FE_PHN3001_n3639;
   wire FE_PHN3000_n4304;
   wire FE_PHN2999_n2804;
   wire FE_PHN2998_n785;
   wire FE_PHN2997_n1448;
   wire FE_PHN2996_n3816;
   wire FE_PHN2995_ram_250__1_;
   wire FE_PHN2994_n1984;
   wire FE_PHN2993_n1553;
   wire FE_PHN2992_n4208;
   wire FE_PHN2991_n1705;
   wire FE_PHN2990_n4109;
   wire FE_PHN2989_n2083;
   wire FE_PHN2988_n2217;
   wire FE_PHN2987_n1350;
   wire FE_PHN2986_n1468;
   wire FE_PHN2985_n2036;
   wire FE_PHN2984_n583;
   wire FE_PHN2983_n588;
   wire FE_PHN2982_n1609;
   wire FE_PHN2981_n1642;
   wire FE_PHN2980_n2111;
   wire FE_PHN2979_ram_46__2_;
   wire FE_PHN2978_n4104;
   wire FE_PHN2977_n3440;
   wire FE_PHN2976_n2471;
   wire FE_PHN2975_n699;
   wire FE_PHN2974_n2506;
   wire FE_PHN2973_n2030;
   wire FE_PHN2972_n1897;
   wire FE_PHN2971_n1103;
   wire FE_PHN2970_n3714;
   wire FE_PHN2969_n2105;
   wire FE_PHN2968_n2445;
   wire FE_PHN2967_n3503;
   wire FE_PHN2966_n1164;
   wire FE_PHN2965_n1336;
   wire FE_PHN2964_n1914;
   wire FE_PHN2963_n1963;
   wire FE_PHN2962_n746;
   wire FE_PHN2961_n3321;
   wire FE_PHN2960_n2869;
   wire FE_PHN2959_n3387;
   wire FE_PHN2958_n1381;
   wire FE_PHN2957_n1727;
   wire FE_PHN2956_n1147;
   wire FE_PHN2955_n2674;
   wire FE_PHN2954_n2793;
   wire FE_PHN2953_n1454;
   wire FE_PHN2952_n2630;
   wire FE_PHN2951_n655;
   wire FE_PHN2950_n1325;
   wire FE_PHN2949_n1750;
   wire FE_PHN2948_n1725;
   wire FE_PHN2947_n3392;
   wire FE_PHN2946_n4497;
   wire FE_PHN2945_n1271;
   wire FE_PHN2944_n2060;
   wire FE_PHN2943_ram_254__9_;
   wire FE_PHN2942_n4667;
   wire FE_PHN2941_n4141;
   wire FE_PHN2940_n3635;
   wire FE_PHN2939_n3540;
   wire FE_PHN2938_n1281;
   wire FE_PHN2937_n3447;
   wire FE_PHN2936_n4093;
   wire FE_PHN2935_n1213;
   wire FE_PHN2934_n4538;
   wire FE_PHN2933_n3786;
   wire FE_PHN2932_n803;
   wire FE_PHN2931_n613;
   wire FE_PHN2930_n2306;
   wire FE_PHN2929_n2546;
   wire FE_PHN2928_n1455;
   wire FE_PHN2927_n3826;
   wire FE_PHN2926_n761;
   wire FE_PHN2925_n1487;
   wire FE_PHN2924_n1407;
   wire FE_PHN2923_n2480;
   wire FE_PHN2922_n2086;
   wire FE_PHN2921_n3275;
   wire FE_PHN2920_n2103;
   wire FE_PHN2919_n3641;
   wire FE_PHN2918_n1807;
   wire FE_PHN2917_n3616;
   wire FE_PHN2916_n3674;
   wire FE_PHN2915_n3372;
   wire FE_PHN2914_n691;
   wire FE_PHN2913_n3370;
   wire FE_PHN2912_n3598;
   wire FE_PHN2911_n1752;
   wire FE_PHN2910_n1779;
   wire FE_PHN2909_n2048;
   wire FE_PHN2908_n1977;
   wire FE_PHN2907_n2320;
   wire FE_PHN2906_n1917;
   wire FE_PHN2905_n1266;
   wire FE_PHN2904_n4462;
   wire FE_PHN2903_n1533;
   wire FE_PHN2902_n1225;
   wire FE_PHN2901_n4606;
   wire FE_PHN2900_n1205;
   wire FE_PHN2899_n1488;
   wire FE_PHN2898_n1748;
   wire FE_PHN2897_n2247;
   wire FE_PHN2896_n2565;
   wire FE_PHN2895_n837;
   wire FE_PHN2894_n3343;
   wire FE_PHN2893_n2065;
   wire FE_PHN2892_n1430;
   wire FE_PHN2891_n702;
   wire FE_PHN2890_n1806;
   wire FE_PHN2889_n1133;
   wire FE_PHN2888_n1309;
   wire FE_PHN2887_n1545;
   wire FE_PHN2886_n2001;
   wire FE_PHN2885_n657;
   wire FE_PHN2884_n4575;
   wire FE_PHN2883_n2310;
   wire FE_PHN2882_n1395;
   wire FE_PHN2881_n1472;
   wire FE_PHN2880_n643;
   wire FE_PHN2879_n1107;
   wire FE_PHN2878_n650;
   wire FE_PHN2877_n2561;
   wire FE_PHN2876_n2043;
   wire FE_PHN2875_n2317;
   wire FE_PHN2874_n2522;
   wire FE_PHN2873_n4341;
   wire FE_PHN2872_n1420;
   wire FE_PHN2871_n633;
   wire FE_PHN2870_n2370;
   wire FE_PHN2869_n3426;
   wire FE_PHN2868_n2078;
   wire FE_PHN2867_n4216;
   wire FE_PHN2866_n3626;
   wire FE_PHN2865_n2093;
   wire FE_PHN2864_n1280;
   wire FE_PHN2863_n1117;
   wire FE_PHN2862_n4460;
   wire FE_PHN2861_n1083;
   wire FE_PHN2860_n684;
   wire FE_PHN2859_n1222;
   wire FE_PHN2858_n1228;
   wire FE_PHN2857_n2453;
   wire FE_PHN2856_n3433;
   wire FE_PHN2855_n3458;
   wire FE_PHN2854_n1602;
   wire FE_PHN2853_n3179;
   wire FE_PHN2852_n1596;
   wire FE_PHN2851_ram_78__8_;
   wire FE_PHN2850_n2575;
   wire FE_PHN2849_ram_104__13_;
   wire FE_PHN2848_n658;
   wire FE_PHN2847_n1848;
   wire FE_PHN2846_n795;
   wire FE_PHN2845_n754;
   wire FE_PHN2844_n2756;
   wire FE_PHN2843_n1457;
   wire FE_PHN2842_n4098;
   wire FE_PHN2841_n2215;
   wire FE_PHN2840_n3830;
   wire FE_PHN2839_n4430;
   wire FE_PHN2838_n1759;
   wire FE_PHN2837_n653;
   wire FE_PHN2836_n645;
   wire FE_PHN2835_n773;
   wire FE_PHN2834_n3631;
   wire FE_PHN2833_n1531;
   wire FE_PHN2832_n3142;
   wire FE_PHN2831_n2517;
   wire FE_PHN2830_n1363;
   wire FE_PHN2829_n623;
   wire FE_PHN2828_ram_120__14_;
   wire FE_PHN2827_n3475;
   wire FE_PHN2826_n2675;
   wire FE_PHN2825_n1290;
   wire FE_PHN2824_n652;
   wire FE_PHN2823_n2817;
   wire FE_PHN2822_n3285;
   wire FE_PHN2821_n719;
   wire FE_PHN2820_n4464;
   wire FE_PHN2819_n3518;
   wire FE_PHN2818_n3669;
   wire FE_PHN2817_n2766;
   wire FE_PHN2816_n3896;
   wire FE_PHN2815_n755;
   wire FE_PHN2814_n1162;
   wire FE_PHN2813_n1687;
   wire FE_PHN2812_n1747;
   wire FE_PHN2811_n629;
   wire FE_PHN2810_n3320;
   wire FE_PHN2809_n3455;
   wire FE_PHN2808_n1476;
   wire FE_PHN2807_n2116;
   wire FE_PHN2806_n1961;
   wire FE_PHN2805_n2109;
   wire FE_PHN2804_n1293;
   wire FE_PHN2803_n711;
   wire FE_PHN2802_ram_45__11_;
   wire FE_PHN2801_n2016;
   wire FE_PHN2800_n4176;
   wire FE_PHN2799_n1823;
   wire FE_PHN2798_n2209;
   wire FE_PHN2797_n710;
   wire FE_PHN2796_n1569;
   wire FE_PHN2795_n3860;
   wire FE_PHN2794_n2050;
   wire FE_PHN2793_n4305;
   wire FE_PHN2792_n4547;
   wire FE_PHN2791_n2479;
   wire FE_PHN2790_n2210;
   wire FE_PHN2789_n2769;
   wire FE_PHN2788_n830;
   wire FE_PHN2787_n3250;
   wire FE_PHN2786_n1264;
   wire FE_PHN2785_n1399;
   wire FE_PHN2784_n1344;
   wire FE_PHN2783_n3331;
   wire FE_PHN2782_n1866;
   wire FE_PHN2781_n1296;
   wire FE_PHN2780_n1341;
   wire FE_PHN2779_n4634;
   wire FE_PHN2778_n3448;
   wire FE_PHN2777_n2235;
   wire FE_PHN2776_n1492;
   wire FE_PHN2775_n3377;
   wire FE_PHN2774_n2282;
   wire FE_PHN2773_n1447;
   wire FE_PHN2772_n3624;
   wire FE_PHN2771_n1365;
   wire FE_PHN2770_n3205;
   wire FE_PHN2769_n4631;
   wire FE_PHN2768_n1481;
   wire FE_PHN2767_n1337;
   wire FE_PHN2766_n2362;
   wire FE_PHN2765_n1268;
   wire FE_PHN2764_n2438;
   wire FE_PHN2763_n1331;
   wire FE_PHN2762_n3272;
   wire FE_PHN2761_n3478;
   wire FE_PHN2760_n2003;
   wire FE_PHN2759_n3445;
   wire FE_PHN2758_n2102;
   wire FE_PHN2757_n1463;
   wire FE_PHN2756_n1501;
   wire FE_PHN2755_n1719;
   wire FE_PHN2754_n2004;
   wire FE_PHN2753_n2542;
   wire FE_PHN2752_n1580;
   wire FE_PHN2751_n2659;
   wire FE_PHN2750_n819;
   wire FE_PHN2749_n3668;
   wire FE_PHN2748_n2723;
   wire FE_PHN2747_n3665;
   wire FE_PHN2746_n1940;
   wire FE_PHN2745_n2037;
   wire FE_PHN2744_n778;
   wire FE_PHN2743_n2470;
   wire FE_PHN2742_n3430;
   wire FE_PHN2741_n2875;
   wire FE_PHN2740_n2256;
   wire FE_PHN2739_n1342;
   wire FE_PHN2738_n2545;
   wire FE_PHN2737_n2113;
   wire FE_PHN2736_n2500;
   wire FE_PHN2735_n1532;
   wire FE_PHN2734_n3409;
   wire FE_PHN2733_n1578;
   wire FE_PHN2732_n1109;
   wire FE_PHN2731_n2002;
   wire FE_PHN2730_n814;
   wire FE_PHN2729_n1127;
   wire FE_PHN2728_n4330;
   wire FE_PHN2727_n2326;
   wire FE_PHN2726_n2066;
   wire FE_PHN2725_n1789;
   wire FE_PHN2724_n681;
   wire FE_PHN2723_n2079;
   wire FE_PHN2722_n799;
   wire FE_PHN2721_n2757;
   wire FE_PHN2720_n664;
   wire FE_PHN2719_n937;
   wire FE_PHN2718_n1200;
   wire FE_PHN2717_n1097;
   wire FE_PHN2716_n2368;
   wire FE_PHN2715_n2351;
   wire FE_PHN2714_n2367;
   wire FE_PHN2713_n3738;
   wire FE_PHN2712_n1739;
   wire FE_PHN2711_n1467;
   wire FE_PHN2710_n4480;
   wire FE_PHN2709_n593;
   wire FE_PHN2708_n2068;
   wire FE_PHN2707_n1931;
   wire FE_PHN2706_n2760;
   wire FE_PHN2705_n1215;
   wire FE_PHN2704_n2359;
   wire FE_PHN2703_n3175;
   wire FE_PHN2702_n2581;
   wire FE_PHN2701_n2758;
   wire FE_PHN2700_n3363;
   wire FE_PHN2699_n2023;
   wire FE_PHN2698_n1912;
   wire FE_PHN2697_n2872;
   wire FE_PHN2696_n2261;
   wire FE_PHN2695_n4428;
   wire FE_PHN2694_n2101;
   wire FE_PHN2693_n1576;
   wire FE_PHN2692_n2790;
   wire FE_PHN2691_n1518;
   wire FE_PHN2690_n2798;
   wire FE_PHN2689_n2462;
   wire FE_PHN2688_n1546;
   wire FE_PHN2687_n3429;
   wire FE_PHN2686_n2059;
   wire FE_PHN2685_n1584;
   wire FE_PHN2684_n1404;
   wire FE_PHN2683_n2447;
   wire FE_PHN2682_n1959;
   wire FE_PHN2681_n1359;
   wire FE_PHN2680_n3893;
   wire FE_PHN2679_n584;
   wire FE_PHN2678_n2248;
   wire FE_PHN2677_n1774;
   wire FE_PHN2676_n2038;
   wire FE_PHN2675_n2759;
   wire FE_PHN2674_n4047;
   wire FE_PHN2673_n1868;
   wire FE_PHN2672_n831;
   wire FE_PHN2671_n1274;
   wire FE_PHN2670_n2478;
   wire FE_PHN2669_n1155;
   wire FE_PHN2668_n2069;
   wire FE_PHN2667_n1791;
   wire FE_PHN2666_n1519;
   wire FE_PHN2665_n2054;
   wire FE_PHN2664_n1927;
   wire FE_PHN2663_n3892;
   wire FE_PHN2662_n3765;
   wire FE_PHN2661_n1398;
   wire FE_PHN2660_n2039;
   wire FE_PHN2659_n2366;
   wire FE_PHN2658_ram_33__9_;
   wire FE_PHN2657_n3525;
   wire FE_PHN2656_n2670;
   wire FE_PHN2655_n2309;
   wire FE_PHN2654_n731;
   wire FE_PHN2653_n1924;
   wire FE_PHN2652_n2241;
   wire FE_PHN2651_n3394;
   wire FE_PHN2650_n2242;
   wire FE_PHN2649_n1555;
   wire FE_PHN2648_n1672;
   wire FE_PHN2647_n2629;
   wire FE_PHN2646_n3792;
   wire FE_PHN2645_n1148;
   wire FE_PHN2644_n2560;
   wire FE_PHN2643_n1744;
   wire FE_PHN2642_n3376;
   wire FE_PHN2641_n2642;
   wire FE_PHN2640_n1278;
   wire FE_PHN2639_n634;
   wire FE_PHN2638_n4605;
   wire FE_PHN2637_n1456;
   wire FE_PHN2636_n1483;
   wire FE_PHN2635_n1786;
   wire FE_PHN2634_n916;
   wire FE_PHN2633_n756;
   wire FE_PHN2632_n2501;
   wire FE_PHN2631_n3617;
   wire FE_PHN2630_n3657;
   wire FE_PHN2629_n2057;
   wire FE_PHN2628_n1216;
   wire FE_PHN2627_n3401;
   wire FE_PHN2626_n1619;
   wire FE_PHN2625_n2871;
   wire FE_PHN2624_n1428;
   wire FE_PHN2623_n4423;
   wire FE_PHN2622_n4090;
   wire FE_PHN2621_n2716;
   wire FE_PHN2620_n1374;
   wire FE_PHN2619_n2035;
   wire FE_PHN2618_n2220;
   wire FE_PHN2617_n1654;
   wire FE_PHN2616_n3782;
   wire FE_PHN2615_n742;
   wire FE_PHN2614_n4205;
   wire FE_PHN2613_n1875;
   wire FE_PHN2612_n2281;
   wire FE_PHN2611_n1436;
   wire FE_PHN2610_n1263;
   wire FE_PHN2609_n1767;
   wire FE_PHN2608_n1421;
   wire FE_PHN2607_n2115;
   wire FE_PHN2606_n2708;
   wire FE_PHN2605_n2008;
   wire FE_PHN2604_n1153;
   wire FE_PHN2603_n2882;
   wire FE_PHN2602_n3567;
   wire FE_PHN2601_n3856;
   wire FE_PHN2600_n1938;
   wire FE_PHN2599_n2117;
   wire FE_PHN2598_ram_45__0_;
   wire FE_PHN2597_ram_93__3_;
   wire FE_PHN2596_n622;
   wire FE_PHN2595_n1808;
   wire FE_PHN2594_n1458;
   wire FE_PHN2593_n1991;
   wire FE_PHN2592_n766;
   wire FE_PHN2591_n1950;
   wire FE_PHN2590_n2224;
   wire FE_PHN2589_n1135;
   wire FE_PHN2588_n598;
   wire FE_PHN2587_n3338;
   wire FE_PHN2586_n1460;
   wire FE_PHN2585_n3252;
   wire FE_PHN2584_n3182;
   wire FE_PHN2583_n1964;
   wire FE_PHN2582_n3692;
   wire FE_PHN2581_n3454;
   wire FE_PHN2580_n3622;
   wire FE_PHN2579_n3647;
   wire FE_PHN2578_n2067;
   wire FE_PHN2577_n1996;
   wire FE_PHN2576_n3878;
   wire FE_PHN2575_n2369;
   wire FE_PHN2574_n1538;
   wire FE_PHN2573_n782;
   wire FE_PHN2572_n2544;
   wire FE_PHN2571_n2535;
   wire FE_PHN2570_n4050;
   wire FE_PHN2569_n3689;
   wire FE_PHN2568_n3235;
   wire FE_PHN2567_n3302;
   wire FE_PHN2566_n1287;
   wire FE_PHN2565_n2504;
   wire FE_PHN2564_n687;
   wire FE_PHN2563_n1177;
   wire FE_PHN2562_n3157;
   wire FE_PHN2561_n3704;
   wire FE_PHN2560_n4079;
   wire FE_PHN2559_n1568;
   wire FE_PHN2558_n4560;
   wire FE_PHN2557_n1674;
   wire FE_PHN2556_n3457;
   wire FE_PHN2555_n2040;
   wire FE_PHN2554_n1551;
   wire FE_PHN2553_n1044;
   wire FE_PHN2552_n1934;
   wire FE_PHN2551_n1723;
   wire FE_PHN2550_n3422;
   wire FE_PHN2549_n1462;
   wire FE_PHN2548_n3898;
   wire FE_PHN2547_n1347;
   wire FE_PHN2546_n1465;
   wire FE_PHN2545_n4569;
   wire FE_PHN2544_n4561;
   wire FE_PHN2543_n3791;
   wire FE_PHN2542_n2669;
   wire FE_PHN2541_n3153;
   wire FE_PHN2540_n2024;
   wire FE_PHN2539_n2502;
   wire FE_PHN2538_n3185;
   wire FE_PHN2537_n3151;
   wire FE_PHN2536_n3437;
   wire FE_PHN2535_n3308;
   wire FE_PHN2534_n2314;
   wire FE_PHN2533_n2663;
   wire FE_PHN2532_n4344;
   wire FE_PHN2531_n939;
   wire FE_PHN2530_n3524;
   wire FE_PHN2529_n3795;
   wire FE_PHN2528_n1156;
   wire FE_PHN2527_n1474;
   wire FE_PHN2526_n1242;
   wire FE_PHN2525_n1343;
   wire FE_PHN2524_n2487;
   wire FE_PHN2523_n3522;
   wire FE_PHN2522_n1513;
   wire FE_PHN2521_n1438;
   wire FE_PHN2520_n3504;
   wire FE_PHN2519_n1283;
   wire FE_PHN2518_n2184;
   wire FE_PHN2517_n1389;
   wire FE_PHN2516_n1662;
   wire FE_PHN2515_n2280;
   wire FE_PHN2514_n3259;
   wire FE_PHN2513_n3654;
   wire FE_PHN2512_n3756;
   wire FE_PHN2511_n627;
   wire FE_PHN2510_n2495;
   wire FE_PHN2509_n1198;
   wire FE_PHN2508_n1383;
   wire FE_PHN2507_n1929;
   wire FE_PHN2506_n2573;
   wire FE_PHN2505_n1400;
   wire FE_PHN2504_n1403;
   wire FE_PHN2503_n3693;
   wire FE_PHN2502_n3603;
   wire FE_PHN2501_n1149;
   wire FE_PHN2500_n1958;
   wire FE_PHN2499_n1894;
   wire FE_PHN2498_n2726;
   wire FE_PHN2497_n2443;
   wire FE_PHN2496_n1070;
   wire FE_PHN2495_n2335;
   wire FE_PHN2494_ram_45__14_;
   wire FE_PHN2493_n1416;
   wire FE_PHN2492_n2448;
   wire FE_PHN2491_n1322;
   wire FE_PHN2490_n2074;
   wire FE_PHN2489_n1573;
   wire FE_PHN2488_n3638;
   wire FE_PHN2487_n3408;
   wire FE_PHN2486_n1589;
   wire FE_PHN2485_n2285;
   wire FE_PHN2484_n3844;
   wire FE_PHN2483_n3903;
   wire FE_PHN2482_n1776;
   wire FE_PHN2481_n1167;
   wire FE_PHN2480_n2534;
   wire FE_PHN2479_n3895;
   wire FE_PHN2478_n642;
   wire FE_PHN2477_n3523;
   wire FE_PHN2476_n2631;
   wire FE_PHN2475_n2483;
   wire FE_PHN2474_n2863;
   wire FE_PHN2473_n1219;
   wire FE_PHN2472_n2693;
   wire FE_PHN2471_n1992;
   wire FE_PHN2470_n1171;
   wire FE_PHN2469_n1464;
   wire FE_PHN2468_n2510;
   wire FE_PHN2467_n3722;
   wire FE_PHN2466_n3432;
   wire FE_PHN2465_n724;
   wire FE_PHN2464_n4437;
   wire FE_PHN2463_n3310;
   wire FE_PHN2462_n1983;
   wire FE_PHN2461_n1434;
   wire FE_PHN2460_n2771;
   wire FE_PHN2459_n2044;
   wire FE_PHN2458_n2706;
   wire FE_PHN2457_n3402;
   wire FE_PHN2456_n1936;
   wire FE_PHN2455_n3242;
   wire FE_PHN2454_ram_81__1_;
   wire FE_PHN2453_n692;
   wire FE_PHN2452_n4128;
   wire FE_PHN2451_n1345;
   wire FE_PHN2450_n3818;
   wire FE_PHN2449_n1469;
   wire FE_PHN2448_n2820;
   wire FE_PHN2447_n3507;
   wire FE_PHN2446_n3144;
   wire FE_PHN2445_n794;
   wire FE_PHN2444_n3500;
   wire FE_PHN2443_n3378;
   wire FE_PHN2442_n2047;
   wire FE_PHN2441_n1050;
   wire FE_PHN2440_n3149;
   wire FE_PHN2439_n2186;
   wire FE_PHN2438_n3614;
   wire FE_PHN2437_n1352;
   wire FE_PHN2436_n1614;
   wire FE_PHN2435_n4675;
   wire FE_PHN2434_n1975;
   wire FE_PHN2433_n2264;
   wire FE_PHN2432_n4615;
   wire FE_PHN2431_n1195;
   wire FE_PHN2430_n700;
   wire FE_PHN2429_n924;
   wire FE_PHN2428_n2559;
   wire FE_PHN2427_n1988;
   wire FE_PHN2426_n2063;
   wire FE_PHN2425_n2336;
   wire FE_PHN2424_n3577;
   wire FE_PHN2423_n1898;
   wire FE_PHN2422_n1994;
   wire FE_PHN2421_n3894;
   wire FE_PHN2420_n1235;
   wire FE_PHN2419_n639;
   wire FE_PHN2418_n1267;
   wire FE_PHN2417_n1486;
   wire FE_PHN2416_n1734;
   wire FE_PHN2415_n4539;
   wire FE_PHN2414_n2795;
   wire FE_PHN2413_n1883;
   wire FE_PHN2412_n2555;
   wire FE_PHN2411_n4614;
   wire FE_PHN2410_n3649;
   wire FE_PHN2409_n2022;
   wire FE_PHN2408_n2562;
   wire FE_PHN2407_n4645;
   wire FE_PHN2406_n1115;
   wire FE_PHN2405_n1284;
   wire FE_PHN2404_n3683;
   wire FE_PHN2403_n1693;
   wire FE_PHN2402_n3630;
   wire FE_PHN2401_n2543;
   wire FE_PHN2400_n738;
   wire FE_PHN2399_n1972;
   wire FE_PHN2398_n3190;
   wire FE_PHN2397_n3855;
   wire FE_PHN2396_n638;
   wire FE_PHN2395_n1778;
   wire FE_PHN2394_n2344;
   wire FE_PHN2393_n1665;
   wire FE_PHN2392_n3417;
   wire FE_PHN2391_n1157;
   wire FE_PHN2390_n3341;
   wire FE_PHN2389_n1997;
   wire FE_PHN2388_n1257;
   wire FE_PHN2387_n3656;
   wire FE_PHN2386_n595;
   wire FE_PHN2385_n834;
   wire FE_PHN2384_n1356;
   wire FE_PHN2383_n635;
   wire FE_PHN2382_n777;
   wire FE_PHN2381_n1857;
   wire FE_PHN2380_n1671;
   wire FE_PHN2379_n1437;
   wire FE_PHN2378_n1876;
   wire FE_PHN2377_n1987;
   wire FE_PHN2376_n732;
   wire FE_PHN2375_n3434;
   wire FE_PHN2374_n2829;
   wire FE_PHN2373_n2087;
   wire FE_PHN2372_n1453;
   wire FE_PHN2371_ram_241__0_;
   wire FE_PHN2370_n4077;
   wire FE_PHN2369_n1970;
   wire FE_PHN2368_n2145;
   wire FE_PHN2367_n2929;
   wire FE_PHN2366_n4309;
   wire FE_PHN2365_n4159;
   wire FE_PHN2364_ram_9__1_;
   wire FE_PHN2363_n3435;
   wire FE_PHN2362_n3723;
   wire FE_PHN2361_n1306;
   wire FE_PHN2360_n2842;
   wire FE_PHN2359_n1762;
   wire FE_PHN2358_n2883;
   wire FE_PHN2357_n1183;
   wire FE_PHN2356_n3148;
   wire FE_PHN2355_n4629;
   wire FE_PHN2354_n2029;
   wire FE_PHN2353_n789;
   wire FE_PHN2352_n3374;
   wire FE_PHN2351_n4549;
   wire FE_PHN2350_n1587;
   wire FE_PHN2349_n4596;
   wire FE_PHN2348_n1974;
   wire FE_PHN2347_n3351;
   wire FE_PHN2346_n673;
   wire FE_PHN2345_n1326;
   wire FE_PHN2344_n1366;
   wire FE_PHN2343_n3707;
   wire FE_PHN2342_n1318;
   wire FE_PHN2341_n4469;
   wire FE_PHN2340_n1530;
   wire FE_PHN2339_n2049;
   wire FE_PHN2338_n2090;
   wire FE_PHN2337_n3750;
   wire FE_PHN2336_n1256;
   wire FE_PHN2335_n1946;
   wire FE_PHN2334_n4073;
   wire FE_PHN2333_n2021;
   wire FE_PHN2332_n2569;
   wire FE_PHN2331_n4482;
   wire FE_PHN2330_n1427;
   wire FE_PHN2329_n3456;
   wire FE_PHN2328_n3849;
   wire FE_PHN2327_n1311;
   wire FE_PHN2326_ram_67__9_;
   wire FE_PHN2325_n646;
   wire FE_PHN2324_n4544;
   wire FE_PHN2323_n3298;
   wire FE_PHN2322_n3776;
   wire FE_PHN2321_n4312;
   wire FE_PHN2320_n2672;
   wire FE_PHN2319_n2550;
   wire FE_PHN2318_n3476;
   wire FE_PHN2317_n4620;
   wire FE_PHN2316_n4513;
   wire FE_PHN2315_n2541;
   wire FE_PHN2314_n1243;
   wire FE_PHN2313_n940;
   wire FE_PHN2312_n685;
   wire FE_PHN2311_n1272;
   wire FE_PHN2310_n3659;
   wire FE_PHN2309_n3858;
   wire FE_PHN2308_n4457;
   wire FE_PHN2307_n4597;
   wire FE_PHN2306_n2302;
   wire FE_PHN2305_n2234;
   wire FE_PHN2304_n955;
   wire FE_PHN2303_n4345;
   wire FE_PHN2302_n3203;
   wire FE_PHN2301_n1303;
   wire FE_PHN2300_n2662;
   wire FE_PHN2299_n4144;
   wire FE_PHN2298_n1796;
   wire FE_PHN2297_n2639;
   wire FE_PHN2296_n3506;
   wire FE_PHN2295_n1512;
   wire FE_PHN2294_n3812;
   wire FE_PHN2293_n3400;
   wire FE_PHN2292_n1591;
   wire FE_PHN2291_n1592;
   wire FE_PHN2290_n3897;
   wire FE_PHN2289_n1441;
   wire FE_PHN2288_ram_45__8_;
   wire FE_PHN2287_n2824;
   wire FE_PHN2286_ram_217__3_;
   wire FE_PHN2285_n3731;
   wire FE_PHN2284_n632;
   wire FE_PHN2283_n1520;
   wire FE_PHN2282_n1208;
   wire FE_PHN2281_n2865;
   wire FE_PHN2280_n4075;
   wire FE_PHN2279_n1294;
   wire FE_PHN2278_n739;
   wire FE_PHN2277_n1223;
   wire FE_PHN2276_n3840;
   wire FE_PHN2275_n3413;
   wire FE_PHN2274_n3701;
   wire FE_PHN2273_n2339;
   wire FE_PHN2272_n1598;
   wire FE_PHN2271_n1788;
   wire FE_PHN2270_n1684;
   wire FE_PHN2269_n2607;
   wire FE_PHN2268_n3779;
   wire FE_PHN2267_n4149;
   wire FE_PHN2266_n705;
   wire FE_PHN2265_n2100;
   wire FE_PHN2264_n1096;
   wire FE_PHN2263_n4301;
   wire FE_PHN2262_n677;
   wire FE_PHN2261_n1638;
   wire FE_PHN2260_n744;
   wire FE_PHN2259_n1482;
   wire FE_PHN2258_n1315;
   wire FE_PHN2257_n3186;
   wire FE_PHN2256_n1201;
   wire FE_PHN2255_n701;
   wire FE_PHN2254_n1224;
   wire FE_PHN2253_n589;
   wire FE_PHN2252_n2755;
   wire FE_PHN2251_n1221;
   wire FE_PHN2250_n1262;
   wire FE_PHN2249_n1517;
   wire FE_PHN2248_n3686;
   wire FE_PHN2247_n2813;
   wire FE_PHN2246_n1660;
   wire FE_PHN2245_n1926;
   wire FE_PHN2244_n1362;
   wire FE_PHN2243_n586;
   wire FE_PHN2242_n760;
   wire FE_PHN2241_n829;
   wire FE_PHN2240_n2528;
   wire FE_PHN2239_n2867;
   wire FE_PHN2238_n4536;
   wire FE_PHN2237_n1120;
   wire FE_PHN2236_n2203;
   wire FE_PHN2235_n2232;
   wire FE_PHN2234_n4100;
   wire FE_PHN2233_n3751;
   wire FE_PHN2232_n604;
   wire FE_PHN2231_n2009;
   wire FE_PHN2230_n2485;
   wire FE_PHN2229_n752;
   wire FE_PHN2228_n2091;
   wire FE_PHN2227_n3237;
   wire FE_PHN2226_n1357;
   wire FE_PHN2225_n747;
   wire FE_PHN2224_n2861;
   wire FE_PHN2223_n716;
   wire FE_PHN2222_n2061;
   wire FE_PHN2221_n3889;
   wire FE_PHN2220_n1677;
   wire FE_PHN2219_n1036;
   wire FE_PHN2218_n1968;
   wire FE_PHN2217_n2322;
   wire FE_PHN2216_n4621;
   wire FE_PHN2215_n599;
   wire FE_PHN2214_n686;
   wire FE_PHN2213_n4042;
   wire FE_PHN2212_n675;
   wire FE_PHN2211_n3405;
   wire FE_PHN2210_n1632;
   wire FE_PHN2209_n2328;
   wire FE_PHN2208_n4654;
   wire FE_PHN2207_n1314;
   wire FE_PHN2206_n3599;
   wire FE_PHN2205_n654;
   wire FE_PHN2204_n1402;
   wire FE_PHN2203_n2239;
   wire FE_PHN2202_n1915;
   wire FE_PHN2201_n1706;
   wire FE_PHN2200_n1794;
   wire FE_PHN2199_n3442;
   wire FE_PHN2198_n2627;
   wire FE_PHN2197_n1291;
   wire FE_PHN2196_n2512;
   wire FE_PHN2195_ram_199__5_;
   wire FE_PHN2194_n3597;
   wire FE_PHN2193_ram_132__8_;
   wire FE_PHN2192_n3716;
   wire FE_PHN2191_n2730;
   wire FE_PHN2190_n1397;
   wire FE_PHN2189_n2854;
   wire FE_PHN2188_n1534;
   wire FE_PHN2187_n2492;
   wire FE_PHN2186_n4314;
   wire FE_PHN2185_n1250;
   wire FE_PHN2184_n3664;
   wire FE_PHN2183_n2319;
   wire FE_PHN2182_n3727;
   wire FE_PHN2181_n1585;
   wire FE_PHN2180_n2293;
   wire FE_PHN2179_n1292;
   wire FE_PHN2178_n1033;
   wire FE_PHN2177_n1755;
   wire FE_PHN2176_n2688;
   wire FE_PHN2175_n4610;
   wire FE_PHN2174_n2551;
   wire FE_PHN2173_n2806;
   wire FE_PHN2172_n2671;
   wire FE_PHN2171_n2558;
   wire FE_PHN2170_n783;
   wire FE_PHN2169_n2694;
   wire FE_PHN2168_n2661;
   wire FE_PHN2167_n1610;
   wire FE_PHN2166_n3345;
   wire FE_PHN2165_n1193;
   wire FE_PHN2164_n1323;
   wire FE_PHN2163_n3602;
   wire FE_PHN2162_n1712;
   wire FE_PHN2161_n1514;
   wire FE_PHN2160_n2707;
   wire FE_PHN2159_n4221;
   wire FE_PHN2158_n1639;
   wire FE_PHN2157_n1199;
   wire FE_PHN2156_n1338;
   wire FE_PHN2155_n3385;
   wire FE_PHN2154_n3799;
   wire FE_PHN2153_n1304;
   wire FE_PHN2152_n4649;
   wire FE_PHN2151_n1658;
   wire FE_PHN2150_n3770;
   wire FE_PHN2149_n745;
   wire FE_PHN2148_n4321;
   wire FE_PHN2147_n3517;
   wire FE_PHN2146_n2606;
   wire FE_PHN2145_n1617;
   wire FE_PHN2144_n4671;
   wire FE_PHN2143_n1636;
   wire FE_PHN2142_n3474;
   wire FE_PHN2141_n1095;
   wire FE_PHN2140_n2814;
   wire FE_PHN2139_n1265;
   wire FE_PHN2138_n668;
   wire FE_PHN2137_n1606;
   wire FE_PHN2136_n1297;
   wire FE_PHN2135_n725;
   wire FE_PHN2134_n2475;
   wire FE_PHN2133_n3901;
   wire FE_PHN2132_n1973;
   wire FE_PHN2131_n1749;
   wire FE_PHN2130_n2513;
   wire FE_PHN2129_n3309;
   wire FE_PHN2128_n1775;
   wire FE_PHN2127_n1246;
   wire FE_PHN2126_n3872;
   wire FE_PHN2125_n4082;
   wire FE_PHN2124_n1557;
   wire FE_PHN2123_n1947;
   wire FE_PHN2122_n2013;
   wire FE_PHN2121_n1594;
   wire FE_PHN2120_n2324;
   wire FE_PHN2119_n2497;
   wire FE_PHN2118_n2291;
   wire FE_PHN2117_n637;
   wire FE_PHN2116_n1270;
   wire FE_PHN2115_n1346;
   wire FE_PHN2114_n1391;
   wire FE_PHN2113_n2216;
   wire FE_PHN2112_n628;
   wire FE_PHN2111_n2646;
   wire FE_PHN2110_n1583;
   wire FE_PHN2109_n3700;
   wire FE_PHN2108_n1151;
   wire FE_PHN2107_n2268;
   wire FE_PHN2106_n1108;
   wire FE_PHN2105_n636;
   wire FE_PHN2104_n2199;
   wire FE_PHN2103_n2096;
   wire FE_PHN2102_n1635;
   wire FE_PHN2101_n4637;
   wire FE_PHN2100_n2202;
   wire FE_PHN2099_n667;
   wire FE_PHN2098_n2509;
   wire FE_PHN2097_n1232;
   wire FE_PHN2096_n1567;
   wire FE_PHN2095_n2249;
   wire FE_PHN2094_n3357;
   wire FE_PHN2093_n4165;
   wire FE_PHN2092_n2062;
   wire FE_PHN2091_n2821;
   wire FE_PHN2090_n2734;
   wire FE_PHN2089_n3431;
   wire FE_PHN2088_n669;
   wire FE_PHN2087_n2318;
   wire FE_PHN2086_n3390;
   wire FE_PHN2085_n3655;
   wire FE_PHN2084_n1168;
   wire FE_PHN2083_n1981;
   wire FE_PHN2082_n1220;
   wire FE_PHN2081_n3594;
   wire FE_PHN2080_n1179;
   wire FE_PHN2079_n2843;
   wire FE_PHN2078_n680;
   wire FE_PHN2077_n2292;
   wire FE_PHN2076_n656;
   wire FE_PHN2075_n1169;
   wire FE_PHN2074_n1424;
   wire FE_PHN2073_n600;
   wire FE_PHN2072_n2731;
   wire FE_PHN2071_n1498;
   wire FE_PHN2070_n1210;
   wire FE_PHN2069_n1646;
   wire FE_PHN2068_n956;
   wire FE_PHN2067_n1414;
   wire FE_PHN2066_n1990;
   wire FE_PHN2065_n3410;
   wire FE_PHN2064_n1537;
   wire FE_PHN2063_n3477;
   wire FE_PHN2062_n4661;
   wire FE_PHN2061_n2056;
   wire FE_PHN2060_n1768;
   wire FE_PHN2059_n1312;
   wire FE_PHN2058_n2547;
   wire FE_PHN2057_n2287;
   wire FE_PHN2056_n3204;
   wire FE_PHN2055_n4117;
   wire FE_PHN2054_n2080;
   wire FE_PHN2053_n3729;
   wire FE_PHN2052_n2690;
   wire FE_PHN2051_n1995;
   wire FE_PHN2050_n3174;
   wire FE_PHN2049_n4585;
   wire FE_PHN2048_n621;
   wire FE_PHN2047_n3253;
   wire FE_PHN2046_n3158;
   wire FE_PHN2045_n3653;
   wire FE_PHN2044_n1659;
   wire FE_PHN2043_n2782;
   wire FE_PHN2042_n4558;
   wire FE_PHN2041_n1415;
   wire FE_PHN2040_n2033;
   wire FE_PHN2039_n2466;
   wire FE_PHN2038_n2529;
   wire FE_PHN2037_n661;
   wire FE_PHN2036_n3764;
   wire FE_PHN2035_n709;
   wire FE_PHN2034_n2237;
   wire FE_PHN2033_n3736;
   wire FE_PHN2032_n1339;
   wire FE_PHN2031_n703;
   wire FE_PHN2030_n2768;
   wire FE_PHN2029_n1209;
   wire FE_PHN2028_n759;
   wire FE_PHN2027_n2350;
   wire FE_PHN2026_n1299;
   wire FE_PHN2025_n4224;
   wire FE_PHN2024_n815;
   wire FE_PHN2023_n1736;
   wire FE_PHN2022_n3590;
   wire FE_PHN2021_n4562;
   wire FE_PHN2020_n1967;
   wire FE_PHN2019_n3269;
   wire FE_PHN2018_n4628;
   wire FE_PHN2017_n4647;
   wire FE_PHN2016_n2449;
   wire FE_PHN2015_n2884;
   wire FE_PHN2014_n2099;
   wire FE_PHN2013_n1590;
   wire FE_PHN2012_n1766;
   wire FE_PHN2011_n2110;
   wire FE_PHN2010_n597;
   wire FE_PHN2009_n1377;
   wire FE_PHN2008_n2832;
   wire FE_PHN2007_n4648;
   wire FE_PHN2006_n4640;
   wire FE_PHN2005_ram_202__13_;
   wire FE_PHN2004_n1319;
   wire FE_PHN2003_n648;
   wire FE_PHN2002_n1966;
   wire FE_PHN2001_n4346;
   wire FE_PHN2000_n1998;
   wire FE_PHN1999_n2252;
   wire FE_PHN1998_n1091;
   wire FE_PHN1997_n2556;
   wire FE_PHN1996_n762;
   wire FE_PHN1995_n2874;
   wire FE_PHN1994_n3824;
   wire FE_PHN1993_n1285;
   wire FE_PHN1992_n3775;
   wire FE_PHN1991_n3382;
   wire FE_PHN1990_n1586;
   wire FE_PHN1989_n1756;
   wire FE_PHN1988_n4298;
   wire FE_PHN1987_n1159;
   wire FE_PHN1986_n1605;
   wire FE_PHN1985_n3420;
   wire FE_PHN1984_n3671;
   wire FE_PHN1983_n1396;
   wire FE_PHN1982_n2014;
   wire FE_PHN1981_n1620;
   wire FE_PHN1980_n2076;
   wire FE_PHN1979_n1648;
   wire FE_PHN1978_n2298;
   wire FE_PHN1977_n1334;
   wire FE_PHN1976_n3715;
   wire FE_PHN1975_n822;
   wire FE_PHN1974_n2357;
   wire FE_PHN1973_n2552;
   wire FE_PHN1972_n2058;
   wire FE_PHN1971_n3416;
   wire FE_PHN1970_n3902;
   wire FE_PHN1969_n1999;
   wire FE_PHN1968_n2748;
   wire FE_PHN1967_n1527;
   wire FE_PHN1966_n1393;
   wire FE_PHN1965_n4074;
   wire FE_PHN1964_n2650;
   wire FE_PHN1963_n3790;
   wire FE_PHN1962_ram_85__10_;
   wire FE_PHN1961_n4115;
   wire FE_PHN1960_n3221;
   wire FE_PHN1959_n1136;
   wire FE_PHN1958_n4489;
   wire FE_PHN1957_n3516;
   wire FE_PHN1956_n695;
   wire FE_PHN1955_n1839;
   wire FE_PHN1954_n720;
   wire FE_PHN1953_n2286;
   wire FE_PHN1952_n714;
   wire FE_PHN1951_n2645;
   wire FE_PHN1950_n2329;
   wire FE_PHN1949_n3496;
   wire FE_PHN1948_n1141;
   wire FE_PHN1947_n2752;
   wire FE_PHN1946_n4101;
   wire FE_PHN1945_n2064;
   wire FE_PHN1944_n2372;
   wire FE_PHN1943_n1928;
   wire FE_PHN1942_n2482;
   wire FE_PHN1941_n1418;
   wire FE_PHN1940_n718;
   wire FE_PHN1939_n1979;
   wire FE_PHN1938_n2010;
   wire FE_PHN1937_n1497;
   wire FE_PHN1936_n3852;
   wire FE_PHN1935_n3884;
   wire FE_PHN1934_n722;
   wire FE_PHN1933_n4357;
   wire FE_PHN1932_n1261;
   wire FE_PHN1931_n1678;
   wire FE_PHN1930_n3719;
   wire FE_PHN1929_n4303;
   wire FE_PHN1928_n2515;
   wire FE_PHN1927_n3247;
   wire FE_PHN1926_n3637;
   wire FE_PHN1925_n1582;
   wire FE_PHN1924_n2676;
   wire FE_PHN1923_n4131;
   wire FE_PHN1922_n682;
   wire FE_PHN1921_n2106;
   wire FE_PHN1920_n1041;
   wire FE_PHN1919_n1564;
   wire FE_PHN1918_n1237;
   wire FE_PHN1917_n1954;
   wire FE_PHN1916_n4200;
   wire FE_PHN1915_n4559;
   wire FE_PHN1914_n3225;
   wire FE_PHN1913_n2316;
   wire FE_PHN1912_n3833;
   wire FE_PHN1911_n2347;
   wire FE_PHN1910_n3381;
   wire FE_PHN1909_n3290;
   wire FE_PHN1908_n2698;
   wire FE_PHN1907_n808;
   wire FE_PHN1906_n2689;
   wire FE_PHN1905_n1884;
   wire FE_PHN1904_n3181;
   wire FE_PHN1903_n1860;
   wire FE_PHN1902_n2810;
   wire FE_PHN1901_n3211;
   wire FE_PHN1900_n3177;
   wire FE_PHN1899_n923;
   wire FE_PHN1898_n2709;
   wire FE_PHN1897_n1410;
   wire FE_PHN1896_n4490;
   wire FE_PHN1895_n3502;
   wire FE_PHN1894_n1258;
   wire FE_PHN1893_n1679;
   wire FE_PHN1892_n1372;
   wire FE_PHN1891_n2830;
   wire FE_PHN1890_n3904;
   wire FE_PHN1889_n1729;
   wire FE_PHN1888_n1925;
   wire FE_PHN1887_n1986;
   wire FE_PHN1886_n2451;
   wire FE_PHN1885_n4454;
   wire FE_PHN1884_n3601;
   wire FE_PHN1883_n2450;
   wire FE_PHN1882_n1641;
   wire FE_PHN1881_n817;
   wire FE_PHN1880_n4336;
   wire FE_PHN1879_n1139;
   wire FE_PHN1878_n1388;
   wire FE_PHN1877_n3667;
   wire FE_PHN1876_n3906;
   wire FE_PHN1875_n2301;
   wire FE_PHN1874_n883;
   wire FE_PHN1873_n4351;
   wire FE_PHN1872_n787;
   wire FE_PHN1871_n3193;
   wire FE_PHN1870_n4650;
   wire FE_PHN1869_n4526;
   wire FE_PHN1868_n1539;
   wire FE_PHN1867_n1933;
   wire FE_PHN1866_n3559;
   wire FE_PHN1865_n4551;
   wire FE_PHN1864_n1234;
   wire FE_PHN1863_n2225;
   wire FE_PHN1862_n2290;
   wire FE_PHN1861_n2045;
   wire FE_PHN1860_n2371;
   wire FE_PHN1859_n2263;
   wire FE_PHN1858_n3605;
   wire FE_PHN1857_n3661;
   wire FE_PHN1856_n792;
   wire FE_PHN1855_n2772;
   wire FE_PHN1854_n2295;
   wire FE_PHN1853_n1516;
   wire FE_PHN1852_n4189;
   wire FE_PHN1851_n3369;
   wire FE_PHN1850_n1333;
   wire FE_PHN1849_n3240;
   wire FE_PHN1848_n1852;
   wire FE_PHN1847_n4674;
   wire FE_PHN1846_n2353;
   wire FE_PHN1845_n3407;
   wire FE_PHN1844_n3850;
   wire FE_PHN1843_n3642;
   wire FE_PHN1842_n2878;
   wire FE_PHN1841_n2114;
   wire FE_PHN1840_n4619;
   wire FE_PHN1839_n1649;
   wire FE_PHN1838_n3184;
   wire FE_PHN1837_n630;
   wire FE_PHN1836_n1535;
   wire FE_PHN1835_n1664;
   wire FE_PHN1834_n1011;
   wire FE_PHN1833_n2847;
   wire FE_PHN1832_n3460;
   wire FE_PHN1831_n3436;
   wire FE_PHN1830_n3444;
   wire FE_PHN1829_n1412;
   wire FE_PHN1828_n3869;
   wire FE_PHN1827_n2729;
   wire FE_PHN1826_n1473;
   wire FE_PHN1825_n3278;
   wire FE_PHN1824_n824;
   wire FE_PHN1823_n3585;
   wire FE_PHN1822_n1738;
   wire FE_PHN1821_n2742;
   wire FE_PHN1820_n1495;
   wire FE_PHN1819_n1810;
   wire FE_PHN1818_n3527;
   wire FE_PHN1817_n2182;
   wire FE_PHN1816_n2913;
   wire FE_PHN1815_n1122;
   wire FE_PHN1814_n2373;
   wire FE_PHN1813_n3787;
   wire FE_PHN1812_n1039;
   wire FE_PHN1811_n3178;
   wire FE_PHN1810_n2827;
   wire FE_PHN1809_n4491;
   wire FE_PHN1808_n2108;
   wire FE_PHN1807_n2469;
   wire FE_PHN1806_n3160;
   wire FE_PHN1805_n4520;
   wire FE_PHN1804_n690;
   wire FE_PHN1803_n726;
   wire FE_PHN1802_n3293;
   wire FE_PHN1801_n807;
   wire FE_PHN1800_n3900;
   wire FE_PHN1799_n1275;
   wire FE_PHN1798_n3593;
   wire FE_PHN1797_n1560;
   wire FE_PHN1796_n1836;
   wire FE_PHN1795_n2668;
   wire FE_PHN1794_n1173;
   wire FE_PHN1793_n2595;
   wire FE_PHN1792_n1321;
   wire FE_PHN1791_n772;
   wire FE_PHN1790_n3662;
   wire FE_PHN1789_n1305;
   wire FE_PHN1788_n1960;
   wire FE_PHN1787_n3412;
   wire FE_PHN1786_n704;
   wire FE_PHN1785_n3428;
   wire FE_PHN1784_n2028;
   wire FE_PHN1783_n4237;
   wire FE_PHN1782_n3612;
   wire FE_PHN1781_ram_63__5_;
   wire FE_PHN1780_n1842;
   wire FE_PHN1779_n4045;
   wire FE_PHN1778_ram_61__13_;
   wire FE_PHN1777_n3270;
   wire FE_PHN1776_n2686;
   wire FE_PHN1775_n1793;
   wire FE_PHN1774_n3146;
   wire FE_PHN1773_n3718;
   wire FE_PHN1772_n670;
   wire FE_PHN1771_n3452;
   wire FE_PHN1770_n4059;
   wire FE_PHN1769_n4152;
   wire FE_PHN1768_n3359;
   wire FE_PHN1767_n4122;
   wire FE_PHN1766_n4145;
   wire FE_PHN1765_n3446;
   wire FE_PHN1764_n3586;
   wire FE_PHN1763_n1477;
   wire FE_PHN1762_n4192;
   wire FE_PHN1761_n4564;
   wire FE_PHN1760_n4184;
   wire FE_PHN1759_n608;
   wire FE_PHN1758_n1724;
   wire FE_PHN1757_n4442;
   wire FE_PHN1756_n4608;
   wire FE_PHN1755_n2279;
   wire FE_PHN1754_n2879;
   wire FE_PHN1753_n1174;
   wire FE_PHN1752_n2764;
   wire FE_PHN1751_n3847;
   wire FE_PHN1750_n3695;
   wire FE_PHN1749_n4052;
   wire FE_PHN1748_n4467;
   wire FE_PHN1747_n1282;
   wire FE_PHN1746_n4484;
   wire FE_PHN1745_n2034;
   wire FE_PHN1744_n591;
   wire FE_PHN1743_n1368;
   wire FE_PHN1742_n3206;
   wire FE_PHN1741_n3256;
   wire FE_PHN1740_n1971;
   wire FE_PHN1739_n2000;
   wire FE_PHN1738_n3281;
   wire FE_PHN1737_n674;
   wire FE_PHN1736_n1549;
   wire FE_PHN1735_n4584;
   wire FE_PHN1734_n3666;
   wire FE_PHN1733_n2255;
   wire FE_PHN1732_n1244;
   wire FE_PHN1731_n2737;
   wire FE_PHN1730_n3627;
   wire FE_PHN1729_n2026;
   wire FE_PHN1728_n3439;
   wire FE_PHN1727_n644;
   wire FE_PHN1726_n1226;
   wire FE_PHN1725_n1295;
   wire FE_PHN1724_n1459;
   wire FE_PHN1723_n2097;
   wire FE_PHN1722_n3450;
   wire FE_PHN1721_n4476;
   wire FE_PHN1720_ram_117__6_;
   wire FE_PHN1719_n4041;
   wire FE_PHN1718_n4530;
   wire FE_PHN1717_n2596;
   wire FE_PHN1716_n2855;
   wire FE_PHN1715_n2015;
   wire FE_PHN1714_n836;
   wire FE_PHN1713_n1390;
   wire FE_PHN1712_n4586;
   wire FE_PHN1711_n2828;
   wire FE_PHN1710_n4591;
   wire FE_PHN1709_n757;
   wire FE_PHN1708_n3316;
   wire FE_PHN1707_n4223;
   wire FE_PHN1706_n3361;
   wire FE_PHN1705_n4529;
   wire FE_PHN1704_n3249;
   wire FE_PHN1703_n2452;
   wire FE_PHN1702_n3232;
   wire FE_PHN1701_n2496;
   wire FE_PHN1700_n3216;
   wire FE_PHN1699_n3495;
   wire FE_PHN1698_n1869;
   wire FE_PHN1697_n4463;
   wire FE_PHN1696_n676;
   wire FE_PHN1695_n3180;
   wire FE_PHN1694_n4563;
   wire FE_PHN1693_n693;
   wire FE_PHN1692_n3709;
   wire FE_PHN1691_n1252;
   wire FE_PHN1690_n3711;
   wire FE_PHN1689_n4468;
   wire FE_PHN1688_n1942;
   wire FE_PHN1687_n2088;
   wire FE_PHN1686_n2345;
   wire FE_PHN1685_n4677;
   wire FE_PHN1684_n696;
   wire FE_PHN1683_n1181;
   wire FE_PHN1682_n1276;
   wire FE_PHN1681_n821;
   wire FE_PHN1680_n1909;
   wire FE_PHN1679_n4234;
   wire FE_PHN1678_n2305;
   wire FE_PHN1677_n4069;
   wire FE_PHN1676_n2834;
   wire FE_PHN1675_n1599;
   wire FE_PHN1674_n1944;
   wire FE_PHN1673_n665;
   wire FE_PHN1672_n3620;
   wire FE_PHN1671_n1853;
   wire FE_PHN1670_n3371;
   wire FE_PHN1669_n764;
   wire FE_PHN1668_n1717;
   wire FE_PHN1667_n3199;
   wire FE_PHN1666_n1939;
   wire FE_PHN1665_n3613;
   wire FE_PHN1664_n1826;
   wire FE_PHN1663_n2191;
   wire FE_PHN1662_n2664;
   wire FE_PHN1661_n1746;
   wire FE_PHN1660_n3785;
   wire FE_PHN1659_n2095;
   wire FE_PHN1658_n771;
   wire FE_PHN1657_n3287;
   wire FE_PHN1656_n1989;
   wire FE_PHN1655_n2640;
   wire FE_PHN1654_n3419;
   wire FE_PHN1653_n1499;
   wire FE_PHN1652_n3825;
   wire FE_PHN1651_n4039;
   wire FE_PHN1650_n1129;
   wire FE_PHN1649_n1098;
   wire FE_PHN1648_n1317;
   wire FE_PHN1647_n1504;
   wire FE_PHN1646_n2666;
   wire FE_PHN1645_n1682;
   wire FE_PHN1644_n1253;
   wire FE_PHN1643_n2311;
   wire FE_PHN1642_n2327;
   wire FE_PHN1641_n2635;
   wire FE_PHN1640_n2660;
   wire FE_PHN1639_n678;
   wire FE_PHN1638_n708;
   wire FE_PHN1637_n1521;
   wire FE_PHN1636_n1631;
   wire FE_PHN1635_n3600;
   wire FE_PHN1634_n4487;
   wire FE_PHN1633_n2548;
   wire FE_PHN1632_n2007;
   wire FE_PHN1631_n2246;
   wire FE_PHN1630_n3187;
   wire FE_PHN1629_n3660;
   wire FE_PHN1628_n3793;
   wire FE_PHN1627_n4492;
   wire FE_PHN1626_n4601;
   wire FE_PHN1625_n1227;
   wire FE_PHN1624_n2323;
   wire FE_PHN1623_n2364;
   wire FE_PHN1622_n3335;
   wire FE_PHN1621_n707;
   wire FE_PHN1620_n1230;
   wire FE_PHN1619_n1544;
   wire FE_PHN1618_n1552;
   wire FE_PHN1617_n1300;
   wire FE_PHN1616_n2303;
   wire FE_PHN1615_n1888;
   wire FE_PHN1614_n2020;
   wire FE_PHN1613_n2860;
   wire FE_PHN1612_n2346;
   wire FE_PHN1611_n671;
   wire FE_PHN1610_n2275;
   wire FE_PHN1609_n1932;
   wire FE_PHN1608_n1238;
   wire FE_PHN1607_n1288;
   wire FE_PHN1606_n1743;
   wire FE_PHN1605_n4140;
   wire FE_PHN1604_n3494;
   wire FE_PHN1603_n3229;
   wire FE_PHN1602_n2525;
   wire FE_PHN1601_n1131;
   wire FE_PHN1600_n2313;
   wire FE_PHN1599_n4472;
   wire FE_PHN1598_n748;
   wire FE_PHN1597_n1505;
   wire FE_PHN1596_n2244;
   wire FE_PHN1595_n3690;
   wire FE_PHN1594_n3294;
   wire FE_PHN1593_n1251;
   wire FE_PHN1592_n3251;
   wire FE_PHN1591_n2864;
   wire FE_PHN1590_n4660;
   wire FE_PHN1589_n767;
   wire FE_PHN1588_n1172;
   wire FE_PHN1587_n786;
   wire FE_PHN1586_n1951;
   wire FE_PHN1585_n2608;
   wire FE_PHN1584_n4653;
   wire FE_PHN1583_n3379;
   wire FE_PHN1582_n3712;
   wire FE_PHN1581_n1655;
   wire FE_PHN1580_n1721;
   wire FE_PHN1579_n1189;
   wire FE_PHN1578_n1204;
   wire FE_PHN1577_n3188;
   wire FE_PHN1576_n582;
   wire FE_PHN1575_n3208;
   wire FE_PHN1574_n1637;
   wire FE_PHN1573_n776;
   wire FE_PHN1572_n835;
   wire FE_PHN1571_n1485;
   wire FE_PHN1570_n3514;
   wire FE_PHN1569_n4592;
   wire FE_PHN1568_n647;
   wire FE_PHN1567_n1822;
   wire FE_PHN1566_n1689;
   wire FE_PHN1565_n3317;
   wire FE_PHN1564_n2233;
   wire FE_PHN1563_n2468;
   wire FE_PHN1562_n3836;
   wire FE_PHN1561_n2725;
   wire FE_PHN1560_n4630;
   wire FE_PHN1559_n2762;
   wire FE_PHN1558_n1114;
   wire FE_PHN1557_n3424;
   wire FE_PHN1556_n1490;
   wire FE_PHN1555_n3314;
   wire FE_PHN1554_n4594;
   wire FE_PHN1553_n1803;
   wire FE_PHN1552_n2025;
   wire FE_PHN1551_n4126;
   wire FE_PHN1550_n698;
   wire FE_PHN1549_n3569;
   wire FE_PHN1548_n3183;
   wire FE_PHN1547_n1548;
   wire FE_PHN1546_n611;
   wire FE_PHN1545_n825;
   wire FE_PHN1544_n2568;
   wire FE_PHN1543_n3330;
   wire FE_PHN1542_n2092;
   wire FE_PHN1541_n3789;
   wire FE_PHN1540_n1478;
   wire FE_PHN1539_n2289;
   wire FE_PHN1538_n1709;
   wire FE_PHN1537_n3305;
   wire FE_PHN1536_n3173;
   wire FE_PHN1535_n2187;
   wire FE_PHN1534_n3539;
   wire FE_PHN1533_n1783;
   wire FE_PHN1532_n2593;
   wire FE_PHN1531_n3652;
   wire FE_PHN1530_n660;
   wire FE_PHN1529_n1307;
   wire FE_PHN1528_n1353;
   wire FE_PHN1527_n1542;
   wire FE_PHN1526_n2881;
   wire FE_PHN1525_n3596;
   wire FE_PHN1524_n1471;
   wire FE_PHN1523_n2539;
   wire FE_PHN1522_n3753;
   wire FE_PHN1521_n1835;
   wire FE_PHN1520_n1623;
   wire FE_PHN1519_n2780;
   wire FE_PHN1518_n3773;
   wire FE_PHN1517_n3867;
   wire FE_PHN1516_n4160;
   wire FE_PHN1515_n3425;
   wire FE_PHN1514_n3696;
   wire FE_PHN1513_n3276;
   wire FE_PHN1512_n1182;
   wire FE_PHN1511_n1556;
   wire FE_PHN1510_n4485;
   wire FE_PHN1509_n4060;
   wire FE_PHN1508_n1895;
   wire FE_PHN1507_n2321;
   wire FE_PHN1506_n816;
   wire FE_PHN1505_n1092;
   wire FE_PHN1504_n3482;
   wire FE_PHN1503_n4154;
   wire FE_PHN1502_n2840;
   wire FE_PHN1501_n1273;
   wire FE_PHN1500_n2006;
   wire FE_PHN1499_n2498;
   wire FE_PHN1498_n626;
   wire FE_PHN1497_n3282;
   wire FE_PHN1496_n1207;
   wire FE_PHN1495_n1335;
   wire FE_PHN1494_n2617;
   wire FE_PHN1493_n587;
   wire FE_PHN1492_n2877;
   wire FE_PHN1491_n3876;
   wire FE_PHN1490_n2198;
   wire FE_PHN1489_n2011;
   wire FE_PHN1488_n3399;
   wire FE_PHN1487_n3672;
   wire FE_PHN1486_n4481;
   wire FE_PHN1485_n1965;
   wire FE_PHN1484_n1830;
   wire FE_PHN1483_n3732;
   wire FE_PHN1482_n780;
   wire FE_PHN1481_n1797;
   wire FE_PHN1480_n1812;
   wire FE_PHN1479_n2656;
   wire FE_PHN1478_n3658;
   wire FE_PHN1477_n1844;
   wire FE_PHN1476_n3933;
   wire FE_PHN1475_n3336;
   wire FE_PHN1474_n4447;
   wire FE_PHN1473_n1308;
   wire FE_PHN1472_n4335;
   wire FE_PHN1471_n2774;
   wire FE_PHN1470_ram_122__2_;
   wire FE_PHN1469_n1071;
   wire FE_PHN1468_n2634;
   wire FE_PHN1467_n1819;
   wire FE_PHN1466_n3268;
   wire FE_PHN1465_n3578;
   wire FE_PHN1464_n3684;
   wire FE_PHN1463_n1625;
   wire FE_PHN1462_n2563;
   wire FE_PHN1461_n1332;
   wire FE_PHN1460_n4543;
   wire FE_PHN1459_n1854;
   wire FE_PHN1458_n3163;
   wire FE_PHN1457_n2315;
   wire FE_PHN1456_n4500;
   wire FE_PHN1455_n614;
   wire FE_PHN1454_n788;
   wire FE_PHN1453_n2490;
   wire FE_PHN1452_n2494;
   wire FE_PHN1451_n2486;
   wire FE_PHN1450_n3347;
   wire FE_PHN1449_n3334;
   wire FE_PHN1448_n2218;
   wire FE_PHN1447_n2705;
   wire FE_PHN1446_n3147;
   wire FE_PHN1445_n3755;
   wire FE_PHN1444_n1125;
   wire FE_PHN1443_n3774;
   wire FE_PHN1442_n1955;
   wire FE_PHN1441_n3393;
   wire FE_PHN1440_n4347;
   wire FE_PHN1439_n2800;
   wire FE_PHN1438_n3582;
   wire FE_PHN1437_n3383;
   wire FE_PHN1436_n3515;
   wire FE_PHN1435_n3823;
   wire FE_PHN1434_n4488;
   wire FE_PHN1433_n1423;
   wire FE_PHN1432_n712;
   wire FE_PHN1431_n1985;
   wire FE_PHN1430_n2557;
   wire FE_PHN1429_n2767;
   wire FE_PHN1428_n3713;
   wire FE_PHN1427_n3705;
   wire FE_PHN1426_n2272;
   wire FE_PHN1425_n4452;
   wire FE_PHN1424_n1138;
   wire FE_PHN1423_n3218;
   wire FE_PHN1422_n1633;
   wire FE_PHN1421_n3414;
   wire FE_PHN1420_n995;
   wire FE_PHN1419_n3886;
   wire FE_PHN1418_n1067;
   wire FE_PHN1417_n826;
   wire FE_PHN1416_n1837;
   wire FE_PHN1415_n3801;
   wire FE_PHN1414_n730;
   wire FE_PHN1413_n3741;
   wire FE_PHN1412_n2822;
   wire FE_PHN1411_n3198;
   wire FE_PHN1410_n4444;
   wire FE_PHN1409_n1541;
   wire FE_PHN1408_n1575;
   wire FE_PHN1407_n1892;
   wire FE_PHN1406_n3415;
   wire FE_PHN1405_n4657;
   wire FE_PHN1404_n2784;
   wire FE_PHN1403_n3529;
   wire FE_PHN1402_n2844;
   wire FE_PHN1401_n1327;
   wire FE_PHN1400_n790;
   wire FE_PHN1399_n774;
   wire FE_PHN1398_n624;
   wire FE_PHN1397_n2530;
   wire FE_PHN1396_n1566;
   wire FE_PHN1395_n4453;
   wire FE_PHN1394_n1211;
   wire FE_PHN1393_n2584;
   wire FE_PHN1392_n3644;
   wire FE_PHN1391_n1180;
   wire FE_PHN1390_n4306;
   wire FE_PHN1389_n4458;
   wire FE_PHN1388_n1763;
   wire FE_PHN1387_n1833;
   wire FE_PHN1386_n3397;
   wire FE_PHN1385_n765;
   wire FE_PHN1384_n3571;
   wire FE_PHN1383_n4089;
   wire FE_PHN1382_n4652;
   wire FE_PHN1381_n3266;
   wire FE_PHN1380_n3395;
   wire FE_PHN1379_n1733;
   wire FE_PHN1378_n1900;
   wire FE_PHN1377_n2537;
   wire FE_PHN1376_n4431;
   wire FE_PHN1375_n4433;
   wire FE_PHN1374_n1185;
   wire FE_PHN1373_n1858;
   wire FE_PHN1372_n2812;
   wire FE_PHN1371_n3703;
   wire FE_PHN1370_n3890;
   wire FE_PHN1369_n2230;
   wire FE_PHN1368_n4108;
   wire FE_PHN1367_n3342;
   wire FE_PHN1366_n3809;
   wire FE_PHN1365_n1202;
   wire FE_PHN1364_n1871;
   wire FE_PHN1363_n3492;
   wire FE_PHN1362_n3391;
   wire FE_PHN1361_n2503;
   wire FE_PHN1360_n2194;
   wire FE_PHN1359_n3196;
   wire FE_PHN1358_n3780;
   wire FE_PHN1357_n1515;
   wire FE_PHN1356_n3691;
   wire FE_PHN1355_n2082;
   wire FE_PHN1354_n3322;
   wire FE_PHN1353_n4432;
   wire FE_PHN1352_n1510;
   wire FE_PHN1351_n1805;
   wire FE_PHN1350_n4051;
   wire FE_PHN1349_n1847;
   wire FE_PHN1348_n2538;
   wire FE_PHN1347_n1907;
   wire FE_PHN1346_n3607;
   wire FE_PHN1345_n3837;
   wire FE_PHN1344_n2643;
   wire FE_PHN1343_n1378;
   wire FE_PHN1342_n3283;
   wire FE_PHN1341_n3834;
   wire FE_PHN1340_n2680;
   wire FE_PHN1339_n2514;
   wire FE_PHN1338_n1466;
   wire FE_PHN1337_n3949;
   wire FE_PHN1336_n4078;
   wire FE_PHN1335_n2819;
   wire FE_PHN1334_n4552;
   wire FE_PHN1333_n3811;
   wire FE_PHN1332_n1073;
   wire FE_PHN1331_n3318;
   wire FE_PHN1330_n1411;
   wire FE_PHN1329_n697;
   wire FE_PHN1328_n1982;
   wire FE_PHN1327_n1364;
   wire FE_PHN1326_n2046;
   wire FE_PHN1325_n2520;
   wire FE_PHN1324_n2940;
   wire FE_PHN1323_n4626;
   wire FE_PHN1322_ram_129__7_;
   wire FE_PHN1321_ram_65__8_;
   wire FE_PHN1320_n3650;
   wire FE_PHN1319_n3303;
   wire FE_PHN1318_ram_81__13_;
   wire FE_PHN1317_n679;
   wire FE_PHN1316_n605;
   wire FE_PHN1315_n3698;
   wire FE_PHN1314_n3488;
   wire FE_PHN1313_n1769;
   wire FE_PHN1312_n2363;
   wire FE_PHN1311_n1217;
   wire FE_PHN1310_n1214;
   wire FE_PHN1309_n3333;
   wire FE_PHN1308_n1075;
   wire FE_PHN1307_n1248;
   wire FE_PHN1306_n3464;
   wire FE_PHN1305_n798;
   wire FE_PHN1304_n1643;
   wire FE_PHN1303_n4455;
   wire FE_PHN1302_n4535;
   wire FE_PHN1301_n2267;
   wire FE_PHN1300_n3145;
   wire FE_PHN1299_n2853;
   wire FE_PHN1298_n3480;
   wire FE_PHN1297_n3717;
   wire FE_PHN1296_n1218;
   wire FE_PHN1295_n2081;
   wire FE_PHN1294_n3788;
   wire FE_PHN1293_n4612;
   wire FE_PHN1292_n3815;
   wire FE_PHN1291_n1409;
   wire FE_PHN1290_n2250;
   wire FE_PHN1289_n3880;
   wire FE_PHN1288_n659;
   wire FE_PHN1287_n1123;
   wire FE_PHN1286_n1846;
   wire FE_PHN1285_n3725;
   wire FE_PHN1284_n3162;
   wire FE_PHN1283_n1930;
   wire FE_PHN1282_n2160;
   wire FE_PHN1281_n4627;
   wire FE_PHN1280_n4157;
   wire FE_PHN1279_n3154;
   wire FE_PHN1278_n4556;
   wire FE_PHN1277_n1240;
   wire FE_PHN1276_n4531;
   wire FE_PHN1275_n1607;
   wire FE_PHN1274_n827;
   wire FE_PHN1273_n1233;
   wire FE_PHN1272_n1241;
   wire FE_PHN1271_n1340;
   wire FE_PHN1270_n1394;
   wire FE_PHN1269_n1550;
   wire FE_PHN1268_n4348;
   wire FE_PHN1267_n4656;
   wire FE_PHN1266_n2658;
   wire FE_PHN1265_n2837;
   wire FE_PHN1264_n810;
   wire FE_PHN1263_n2684;
   wire FE_PHN1262_n2296;
   wire FE_PHN1261_n3368;
   wire FE_PHN1260_n3521;
   wire FE_PHN1259_n3215;
   wire FE_PHN1258_n4127;
   wire FE_PHN1257_n1668;
   wire FE_PHN1256_n4483;
   wire FE_PHN1255_n3315;
   wire FE_PHN1254_n1140;
   wire FE_PHN1253_n2342;
   wire FE_PHN1252_n2792;
   wire FE_PHN1251_n1651;
   wire FE_PHN1250_n4354;
   wire FE_PHN1249_n1728;
   wire FE_PHN1248_n4534;
   wire FE_PHN1247_n4264;
   wire FE_PHN1246_n4611;
   wire FE_PHN1245_n2823;
   wire FE_PHN1244_n2591;
   wire FE_PHN1243_n2283;
   wire FE_PHN1242_n1758;
   wire FE_PHN1241_n4061;
   wire FE_PHN1240_n1666;
   wire FE_PHN1239_n2228;
   wire FE_PHN1238_n2620;
   wire FE_PHN1237_n3806;
   wire FE_PHN1236_n1379;
   wire FE_PHN1235_n1903;
   wire FE_PHN1234_n2641;
   wire FE_PHN1233_n2931;
   wire FE_PHN1232_n2657;
   wire FE_PHN1231_n3227;
   wire FE_PHN1230_n805;
   wire FE_PHN1229_n2745;
   wire FE_PHN1228_n3189;
   wire FE_PHN1227_n2687;
   wire FE_PHN1226_n1867;
   wire FE_PHN1225_n2491;
   wire FE_PHN1224_n2763;
   wire FE_PHN1223_n683;
   wire FE_PHN1222_n1849;
   wire FE_PHN1221_n1348;
   wire FE_PHN1220_n2699;
   wire FE_PHN1219_n2838;
   wire FE_PHN1218_n4505;
   wire FE_PHN1217_n3581;
   wire FE_PHN1216_n3615;
   wire FE_PHN1215_n3831;
   wire FE_PHN1214_n4177;
   wire FE_PHN1213_n2457;
   wire FE_PHN1212_n4546;
   wire FE_PHN1211_n3406;
   wire FE_PHN1210_n3291;
   wire FE_PHN1209_n4550;
   wire FE_PHN1208_n2794;
   wire FE_PHN1207_n1192;
   wire FE_PHN1206_n2300;
   wire FE_PHN1205_n1670;
   wire FE_PHN1204_n3200;
   wire FE_PHN1203_n3845;
   wire FE_PHN1202_n1881;
   wire FE_PHN1201_n3841;
   wire FE_PHN1200_n1685;
   wire FE_PHN1199_n3583;
   wire FE_PHN1198_n3161;
   wire FE_PHN1197_n2644;
   wire FE_PHN1196_n1385;
   wire FE_PHN1195_n3264;
   wire FE_PHN1194_n1953;
   wire FE_PHN1193_n2862;
   wire FE_PHN1192_n2579;
   wire FE_PHN1191_n1862;
   wire FE_PHN1190_n2679;
   wire FE_PHN1189_n2831;
   wire FE_PHN1188_n2677;
   wire FE_PHN1187_n3398;
   wire FE_PHN1186_n1231;
   wire FE_PHN1185_n1371;
   wire FE_PHN1184_n4617;
   wire FE_PHN1183_n963;
   wire FE_PHN1182_n2777;
   wire FE_PHN1181_n2018;
   wire FE_PHN1180_n2724;
   wire FE_PHN1179_n3851;
   wire FE_PHN1178_n2190;
   wire FE_PHN1177_n3636;
   wire FE_PHN1176_n3299;
   wire FE_PHN1175_n3873;
   wire FE_PHN1174_n3859;
   wire FE_PHN1173_n2308;
   wire FE_PHN1172_n2524;
   wire FE_PHN1171_n3197;
   wire FE_PHN1170_n1603;
   wire FE_PHN1169_n2567;
   wire FE_PHN1168_n1698;
   wire FE_PHN1167_n3728;
   wire FE_PHN1166_n3899;
   wire FE_PHN1165_n833;
   wire FE_PHN1164_n3566;
   wire FE_PHN1163_n3752;
   wire FE_PHN1162_n1840;
   wire FE_PHN1161_n2825;
   wire FE_PHN1160_n3821;
   wire FE_PHN1159_n3340;
   wire FE_PHN1158_n2833;
   wire FE_PHN1157_n3813;
   wire FE_PHN1156_n4470;
   wire FE_PHN1155_n3304;
   wire FE_PHN1154_n3325;
   wire FE_PHN1153_n3411;
   wire FE_PHN1152_n2685;
   wire FE_PHN1151_n3802;
   wire FE_PHN1150_n1732;
   wire FE_PHN1149_n2231;
   wire FE_PHN1148_n1196;
   wire FE_PHN1147_n3808;
   wire FE_PHN1146_n1370;
   wire FE_PHN1145_n3766;
   wire FE_PHN1144_n1084;
   wire FE_PHN1143_n3820;
   wire FE_PHN1142_n1588;
   wire FE_PHN1141_n4607;
   wire FE_PHN1140_n2325;
   wire FE_PHN1139_n2816;
   wire FE_PHN1138_n2472;
   wire FE_PHN1137_n1581;
   wire FE_PHN1136_n3214;
   wire FE_PHN1135_n2791;
   wire FE_PHN1134_n4673;
   wire FE_PHN1133_n4511;
   wire FE_PHN1132_n3346;
   wire FE_PHN1131_n3835;
   wire FE_PHN1130_n2738;
   wire FE_PHN1129_n3687;
   wire FE_PHN1128_n2442;
   wire FE_PHN1127_n2072;
   wire FE_PHN1126_n1877;
   wire FE_PHN1125_n1563;
   wire FE_PHN1124_n1661;
   wire FE_PHN1123_n2681;
   wire FE_PHN1122_n4133;
   wire FE_PHN1121_n3874;
   wire FE_PHN1120_n1673;
   wire FE_PHN1119_n3057;
   wire FE_PHN1118_n3192;
   wire FE_PHN1117_n1387;
   wire FE_PHN1116_n1503;
   wire FE_PHN1115_n1621;
   wire FE_PHN1114_n1558;
   wire FE_PHN1113_n672;
   wire FE_PHN1112_n1976;
   wire FE_PHN1111_n2704;
   wire FE_PHN1110_n3595;
   wire FE_PHN1109_n1949;
   wire FE_PHN1108_n3228;
   wire FE_PHN1107_n1554;
   wire FE_PHN1106_n1910;
   wire FE_PHN1105_n2188;
   wire FE_PHN1104_n2858;
   wire FE_PHN1103_n4250;
   wire FE_PHN1102_n3045;
   wire FE_PHN1101_n1386;
   wire FE_PHN1100_n2807;
   wire FE_PHN1099_n4124;
   wire FE_PHN1098_n3279;
   wire FE_PHN1097_n1245;
   wire FE_PHN1096_n3623;
   wire FE_PHN1095_n2713;
   wire FE_PHN1094_n3373;
   wire FE_PHN1093_n3588;
   wire FE_PHN1092_n2070;
   wire FE_PHN1091_n2193;
   wire FE_PHN1090_n2481;
   wire FE_PHN1089_n3348;
   wire FE_PHN1088_n4445;
   wire FE_PHN1087_n4593;
   wire FE_PHN1086_n2195;
   wire FE_PHN1085_n3039;
   wire FE_PHN1084_n1130;
   wire FE_PHN1083_n1444;
   wire FE_PHN1082_n908;
   wire FE_PHN1081_n1500;
   wire FE_PHN1080_n2785;
   wire FE_PHN1079_n1113;
   wire FE_PHN1078_n3758;
   wire FE_PHN1077_n4666;
   wire FE_PHN1076_n2226;
   wire FE_PHN1075_n2924;
   wire FE_PHN1074_n1360;
   wire FE_PHN1073_n1923;
   wire FE_PHN1072_n2682;
   wire FE_PHN1071_n1260;
   wire FE_PHN1070_n1522;
   wire FE_PHN1069_n1742;
   wire FE_PHN1068_n2189;
   wire FE_PHN1067_n3604;
   wire FE_PHN1066_n607;
   wire FE_PHN1065_n4537;
   wire FE_PHN1064_n784;
   wire FE_PHN1063_n1102;
   wire FE_PHN1062_n3721;
   wire FE_PHN1061_n4588;
   wire FE_PHN1060_n4598;
   wire FE_PHN1059_n689;
   wire FE_PHN1058_ram_201__5_;
   wire FE_PHN1057_n4427;
   wire FE_PHN1056_n4322;
   wire FE_PHN1055_n2917;
   wire FE_PHN1054_n1785;
   wire FE_PHN1053_n2027;
   wire FE_PHN1052_n4197;
   wire FE_PHN1051_n618;
   wire FE_PHN1050_n3814;
   wire FE_PHN1049_n4048;
   wire FE_PHN1048_n3706;
   wire FE_PHN1047_n3155;
   wire FE_PHN1046_n663;
   wire FE_PHN1045_n615;
   wire FE_PHN1044_n4040;
   wire FE_PHN1043_n926;
   wire FE_PHN1042_n1855;
   wire FE_PHN1041_n2493;
   wire FE_PHN1040_n3339;
   wire FE_PHN1039_n2474;
   wire FE_PHN1038_n3403;
   wire FE_PHN1037_n3396;
   wire FE_PHN1036_n4499;
   wire FE_PHN1035_n1824;
   wire FE_PHN1034_n2649;
   wire FE_PHN1033_n3449;
   wire FE_PHN1032_n4088;
   wire FE_PHN1031_n4086;
   wire FE_PHN1030_n4478;
   wire FE_PHN1029_n4429;
   wire FE_PHN1028_n2416;
   wire FE_PHN1027_n2526;
   wire FE_PHN1026_n823;
   wire FE_PHN1025_n1843;
   wire FE_PHN1024_n2075;
   wire FE_PHN1023_n2213;
   wire FE_PHN1022_n2387;
   wire FE_PHN1021_n4067;
   wire FE_PHN1020_n4112;
   wire FE_PHN1019_n1384;
   wire FE_PHN1018_n1628;
   wire FE_PHN1017_n3681;
   wire FE_PHN1016_n1718;
   wire FE_PHN1015_n2851;
   wire FE_PHN1014_n2477;
   wire FE_PHN1013_n3740;
   wire FE_PHN1012_n4672;
   wire FE_PHN1011_n1507;
   wire FE_PHN1010_n1943;
   wire FE_PHN1009_n4071;
   wire FE_PHN1008_n617;
   wire FE_PHN1007_n1432;
   wire FE_PHN1006_n2192;
   wire FE_PHN1005_n1442;
   wire FE_PHN1004_n3273;
   wire FE_PHN1003_n2019;
   wire FE_PHN1002_n3326;
   wire FE_PHN1001_n1893;
   wire FE_PHN1000_n3646;
   wire FE_PHN999_n4616;
   wire FE_PHN998_n1809;
   wire FE_PHN997_n2846;
   wire FE_PHN996_n4486;
   wire FE_PHN995_n1832;
   wire FE_PHN994_n3384;
   wire FE_PHN993_n3794;
   wire FE_PHN992_n1669;
   wire FE_PHN991_n4646;
   wire FE_PHN990_n1528;
   wire FE_PHN989_n3553;
   wire FE_PHN988_n3865;
   wire FE_PHN987_n3726;
   wire FE_PHN986_n2332;
   wire FE_PHN985_n1124;
   wire FE_PHN984_n1506;
   wire FE_PHN983_n1980;
   wire FE_PHN982_n694;
   wire FE_PHN981_n1408;
   wire FE_PHN980_n2042;
   wire FE_PHN979_n2836;
   wire FE_PHN978_n1351;
   wire FE_PHN977_n4053;
   wire FE_PHN976_n4063;
   wire FE_PHN975_n2856;
   wire FE_PHN974_n2866;
   wire FE_PHN973_n4664;
   wire FE_PHN972_n2440;
   wire FE_PHN971_n2775;
   wire FE_PHN970_n2243;
   wire FE_PHN969_n662;
   wire FE_PHN968_n1645;
   wire FE_PHN967_n1329;
   wire FE_PHN966_n1081;
   wire FE_PHN965_n3883;
   wire FE_PHN964_n2736;
   wire FE_PHN963_n3589;
   wire FE_PHN962_n2077;
   wire FE_PHN961_n4450;
   wire FE_PHN960_n3505;
   wire FE_PHN959_n1126;
   wire FE_PHN958_n4676;
   wire FE_PHN957_n3441;
   wire FE_PHN956_n1450;
   wire FE_PHN955_n3839;
   wire FE_PHN954_n4272;
   wire FE_PHN953_n4524;
   wire FE_PHN952_n3822;
   wire FE_PHN951_n1565;
   wire FE_PHN950_n1851;
   wire FE_PHN949_n2533;
   wire FE_PHN948_n3195;
   wire FE_PHN947_n4624;
   wire FE_PHN946_n2454;
   wire FE_PHN945_n3254;
   wire FE_PHN944_n3289;
   wire FE_PHN943_n4641;
   wire FE_PHN942_n3311;
   wire FE_PHN941_n779;
   wire FE_PHN940_n2848;
   wire FE_PHN939_n3202;
   wire FE_PHN938_n1446;
   wire FE_PHN937_n1152;
   wire FE_PHN936_n3648;
   wire FE_PHN935_n2128;
   wire FE_PHN934_n813;
   wire FE_PHN933_n942;
   wire FE_PHN932_n1165;
   wire FE_PHN931_n1439;
   wire FE_PHN930_n2518;
   wire FE_PHN929_n1627;
   wire FE_PHN928_n2094;
   wire FE_PHN927_n1380;
   wire FE_PHN926_n1845;
   wire FE_PHN925_n3159;
   wire FE_PHN924_n4156;
   wire FE_PHN923_n1523;
   wire FE_PHN922_n606;
   wire FE_PHN921_n4528;
   wire FE_PHN920_n2638;
   wire FE_PHN919_n3530;
   wire FE_PHN918_n1433;
   wire FE_PHN917_n3576;
   wire FE_PHN916_n1890;
   wire FE_PHN915_n1745;
   wire FE_PHN914_n1570;
   wire FE_PHN913_n3767;
   wire FE_PHN912_n3628;
   wire FE_PHN911_n1667;
   wire FE_PHN910_n2334;
   wire FE_PHN909_n3737;
   wire FE_PHN908_n1184;
   wire FE_PHN907_n1675;
   wire FE_PHN906_n3804;
   wire FE_PHN905_n1841;
   wire FE_PHN904_n3685;
   wire FE_PHN903_n3829;
   wire FE_PHN902_n4595;
   wire FE_PHN901_n2808;
   wire FE_PHN900_n4625;
   wire FE_PHN899_n1100;
   wire FE_PHN898_n3907;
   wire FE_PHN897_n2312;
   wire FE_PHN896_n2197;
   wire FE_PHN895_n1715;
   wire FE_PHN894_n3360;
   wire FE_PHN893_n800;
   wire FE_PHN892_n2849;
   wire FE_PHN891_n3761;
   wire FE_PHN890_n4422;
   wire FE_PHN889_n4498;
   wire FE_PHN888_n932;
   wire FE_PHN887_n2221;
   wire FE_PHN886_n2439;
   wire FE_PHN885_n1811;
   wire FE_PHN884_n4516;
   wire FE_PHN883_n2352;
   wire FE_PHN882_n3248;
   wire FE_PHN881_n2484;
   wire FE_PHN880_n2751;
   wire FE_PHN879_n3832;
   wire FE_PHN878_n4572;
   wire FE_PHN877_n818;
   wire FE_PHN876_n612;
   wire FE_PHN875_n1188;
   wire FE_PHN874_n775;
   wire FE_PHN873_n1801;
   wire FE_PHN872_n2809;
   wire FE_PHN871_ram_249__12_;
   wire FE_PHN870_n1128;
   wire FE_PHN869_n3745;
   wire FE_PHN868_n4253;
   wire FE_PHN867_n2776;
   wire FE_PHN866_n3828;
   wire FE_PHN865_n1777;
   wire FE_PHN864_n3404;
   wire FE_PHN863_n4136;
   wire FE_PHN862_n3879;
   wire FE_PHN861_n4545;
   wire FE_PHN860_n3486;
   wire FE_PHN859_n3176;
   wire FE_PHN858_n4293;
   wire FE_PHN857_n1191;
   wire FE_PHN856_n2253;
   wire FE_PHN855_n4337;
   wire FE_PHN854_n741;
   wire FE_PHN853_n3720;
   wire FE_PHN852_n3760;
   wire FE_PHN851_n3307;
   wire FE_PHN850_n4085;
   wire FE_PHN849_n4523;
   wire FE_PHN848_n723;
   wire FE_PHN847_n4058;
   wire FE_PHN846_n4198;
   wire FE_PHN845_n1800;
   wire FE_PHN844_n3288;
   wire FE_PHN843_n4099;
   wire FE_PHN842_n3296;
   wire FE_PHN841_n3551;
   wire FE_PHN840_n2899;
   wire FE_PHN839_n875;
   wire FE_PHN838_n3675;
   wire FE_PHN837_n1089;
   wire FE_PHN836_n3271;
   wire FE_PHN835_n1170;
   wire FE_PHN834_n1827;
   wire FE_PHN833_n2939;
   wire FE_PHN832_n1004;
   wire FE_PHN831_n1479;
   wire FE_PHN830_n2129;
   wire FE_PHN829_n3201;
   wire FE_PHN828_n3222;
   wire FE_PHN827_n3643;
   wire FE_PHN826_n2418;
   wire FE_PHN825_n3418;
   wire FE_PHN824_n3925;
   wire FE_PHN823_n1526;
   wire FE_PHN822_n1187;
   wire FE_PHN821_n3528;
   wire FE_PHN820_n2307;
   wire FE_PHN819_n4473;
   wire FE_PHN818_n2835;
   wire FE_PHN817_n1502;
   wire FE_PHN816_n859;
   wire FE_PHN815_n3423;
   wire FE_PHN814_n3485;
   wire FE_PHN813_n2717;
   wire FE_PHN812_n2797;
   wire FE_PHN811_n3724;
   wire FE_PHN810_n3871;
   wire FE_PHN809_n1440;
   wire FE_PHN808_n1524;
   wire FE_PHN807_n1882;
   wire FE_PHN806_n2947;
   wire FE_PHN805_n3168;
   wire FE_PHN804_n751;
   wire FE_PHN803_n1255;
   wire FE_PHN802_n1650;
   wire FE_PHN801_n4651;
   wire FE_PHN800_n1561;
   wire FE_PHN799_n1683;
   wire FE_PHN798_n2488;
   wire FE_PHN797_n1612;
   wire FE_PHN796_n2107;
   wire FE_PHN795_n2781;
   wire FE_PHN794_n4521;
   wire FE_PHN793_n2404;
   wire FE_PHN792_n1751;
   wire FE_PHN791_n2799;
   wire FE_PHN790_n3244;
   wire FE_PHN789_n4424;
   wire FE_PHN788_n2678;
   wire FE_PHN787_n1629;
   wire FE_PHN786_n2150;
   wire FE_PHN785_n3306;
   wire FE_PHN784_n4555;
   wire FE_PHN783_n4638;
   wire FE_PHN782_n3421;
   wire FE_PHN781_n4663;
   wire FE_PHN780_n2260;
   wire FE_PHN779_n3710;
   wire FE_PHN778_n3796;
   wire FE_PHN777_n4066;
   wire FE_PHN776_n2459;
   wire FE_PHN775_n619;
   wire FE_PHN774_n1597;
   wire FE_PHN773_n3238;
   wire FE_PHN772_n3708;
   wire FE_PHN771_n4554;
   wire FE_PHN770_n3366;
   wire FE_PHN769_n3699;
   wire FE_PHN768_n2597;
   wire FE_PHN767_n3587;
   wire FE_PHN766_n4425;
   wire FE_PHN765_n4072;
   wire FE_PHN764_n860;
   wire FE_PHN763_n3324;
   wire FE_PHN762_n3465;
   wire FE_PHN761_n4287;
   wire FE_PHN760_n1720;
   wire FE_PHN759_n3479;
   wire FE_PHN758_n4083;
   wire FE_PHN757_n603;
   wire FE_PHN756_n2436;
   wire FE_PHN755_n3349;
   wire FE_PHN754_n3645;
   wire FE_PHN753_n640;
   wire FE_PHN752_n1057;
   wire FE_PHN751_n1475;
   wire FE_PHN750_n1105;
   wire FE_PHN749_n1145;
   wire FE_PHN748_n1657;
   wire FE_PHN747_n2783;
   wire FE_PHN746_n2143;
   wire FE_PHN745_n750;
   wire FE_PHN744_n1680;
   wire FE_PHN743_n2222;
   wire FE_PHN742_n4113;
   wire FE_PHN741_n3885;
   wire FE_PHN740_n4302;
   wire FE_PHN739_n1885;
   wire FE_PHN738_n3277;
   wire FE_PHN737_n3853;
   wire FE_PHN736_n2085;
   wire FE_PHN735_n2219;
   wire FE_PHN734_n1604;
   wire FE_PHN733_n2084;
   wire FE_PHN732_n3194;
   wire FE_PHN731_n2441;
   wire FE_PHN730_n3356;
   wire FE_PHN729_n728;
   wire FE_PHN728_n1716;
   wire FE_PHN727_n2211;
   wire FE_PHN726_n3171;
   wire FE_PHN725_n4349;
   wire FE_PHN724_n4518;
   wire FE_PHN723_n3573;
   wire FE_PHN722_n4659;
   wire FE_PHN721_n4501;
   wire FE_PHN720_n4519;
   wire FE_PHN719_n1703;
   wire FE_PHN718_n733;
   wire FE_PHN717_n1052;
   wire FE_PHN716_n1608;
   wire FE_PHN715_n2173;
   wire FE_PHN714_n4091;
   wire FE_PHN713_n1144;
   wire FE_PHN712_n1298;
   wire FE_PHN711_n3511;
   wire FE_PHN710_n1820;
   wire FE_PHN709_n3733;
   wire FE_PHN708_n3941;
   wire FE_PHN707_n3651;
   wire FE_PHN706_n3061;
   wire FE_PHN705_n3267;
   wire FE_PHN704_n3575;
   wire FE_PHN703_n2739;
   wire FE_PHN702_n2271;
   wire FE_PHN701_n3875;
   wire FE_PHN700_n4495;
   wire FE_PHN699_n3759;
   wire FE_PHN698_n2911;
   wire FE_PHN697_n2905;
   wire FE_PHN696_n820;
   wire FE_PHN695_n4056;
   wire FE_PHN694_n4668;
   wire FE_PHN693_n1480;
   wire FE_PHN692_n3498;
   wire FE_PHN691_n1831;
   wire FE_PHN690_n2269;
   wire FE_PHN689_n2276;
   wire FE_PHN688_n2811;
   wire FE_PHN687_n1887;
   wire FE_PHN686_n1889;
   wire FE_PHN685_n4436;
   wire FE_PHN684_n4532;
   wire FE_PHN683_n1647;
   wire FE_PHN682_n4643;
   wire FE_PHN681_n1771;
   wire FE_PHN680_n4669;
   wire FE_PHN679_n4434;
   wire FE_PHN678_n1175;
   wire FE_PHN677_n1496;
   wire FE_PHN676_n2673;
   wire FE_PHN675_n3113;
   wire FE_PHN674_n1494;
   wire FE_PHN673_n2914;
   wire FE_PHN672_n2527;
   wire FE_PHN671_n2507;
   wire FE_PHN670_n4459;
   wire FE_PHN669_n4665;
   wire FE_PHN668_n1247;
   wire FE_PHN667_n1367;
   wire FE_PHN666_n3702;
   wire FE_PHN665_n4576;
   wire FE_PHN664_n2139;
   wire FE_PHN663_ram_109__5_;
   wire FE_PHN662_n4517;
   wire FE_PHN661_n2270;
   wire FE_PHN660_n1445;
   wire FE_PHN659_n1740;
   wire FE_PHN658_n3882;
   wire FE_PHN657_n3297;
   wire FE_PHN656_n2519;
   wire FE_PHN655_n4639;
   wire FE_PHN654_n1249;
   wire FE_PHN653_n1640;
   wire FE_PHN652_n1697;
   wire FE_PHN651_n2655;
   wire FE_PHN650_n2463;
   wire FE_PHN649_n3059;
   wire FE_PHN648_n1035;
   wire FE_PHN647_n1828;
   wire FE_PHN646_n2532;
   wire FE_PHN645_n3312;
   wire FE_PHN644_n3313;
   wire FE_PHN643_n3501;
   wire FE_PHN642_n2852;
   wire FE_PHN641_n1559;
   wire FE_PHN640_n3245;
   wire FE_PHN639_n4443;
   wire FE_PHN638_n3591;
   wire FE_PHN637_n1176;
   wire FE_PHN636_n3513;
   wire FE_PHN635_n1116;
   wire FE_PHN634_n2710;
   wire FE_PHN633_n4618;
   wire FE_PHN632_n666;
   wire FE_PHN631_n1493;
   wire FE_PHN630_n1798;
   wire FE_PHN629_n2444;
   wire FE_PHN628_n2508;
   wire FE_PHN627_n2895;
   wire FE_PHN626_n4590;
   wire FE_PHN625_n4599;
   wire FE_PHN624_n4280;
   wire FE_PHN623_n806;
   wire FE_PHN622_n2238;
   wire FE_PHN621_n3973;
   wire FE_PHN620_n2288;
   wire FE_PHN619_n2632;
   wire FE_PHN618_n4095;
   wire FE_PHN617_n1861;
   wire FE_PHN616_n4161;
   wire FE_PHN615_n3344;
   wire FE_PHN614_n1160;
   wire FE_PHN613_n2850;
   wire FE_PHN612_n2586;
   wire FE_PHN611_n1547;
   wire FE_PHN610_n3909;
   wire FE_PHN609_n4451;
   wire FE_PHN608_n2089;
   wire FE_PHN607_n3680;
   wire FE_PHN606_n1760;
   wire FE_PHN605_n1722;
   wire FE_PHN604_n4080;
   wire FE_PHN603_n1431;
   wire FE_PHN602_n1821;
   wire FE_PHN601_n602;
   wire FE_PHN600_n2265;
   wire FE_PHN599_n2585;
   wire FE_PHN598_n4466;
   wire FE_PHN597_n3468;
   wire FE_PHN596_n3663;
   wire FE_PHN595_n3438;
   wire FE_PHN594_n1834;
   wire FE_PHN593_n2284;
   wire FE_PHN592_n2553;
   wire FE_PHN591_n1702;
   wire FE_PHN590_n2229;
   wire FE_PHN589_n2721;
   wire FE_PHN588_n2859;
   wire FE_PHN587_n4623;
   wire FE_PHN586_n3509;
   wire FE_PHN585_n931;
   wire FE_PHN584_n3386;
   wire FE_PHN583_n3887;
   wire FE_PHN582_n1878;
   wire FE_PHN581_n2826;
   wire FE_PHN580_n1186;
   wire FE_PHN579_n3510;
   wire FE_PHN578_n3781;
   wire FE_PHN577_n3800;
   wire FE_PHN576_n4296;
   wire FE_PHN575_n2683;
   wire FE_PHN574_n740;
   wire FE_PHN573_n3246;
   wire FE_PHN572_n1085;
   wire FE_PHN571_n3560;
   wire FE_PHN570_n3868;
   wire FE_PHN569_n3537;
   wire FE_PHN568_n4440;
   wire FE_PHN567_n4604;
   wire FE_PHN566_n1616;
   wire FE_PHN565_n2583;
   wire FE_PHN564_n753;
   wire FE_PHN563_n2691;
   wire FE_PHN562_n3470;
   wire FE_PHN561_n3472;
   wire FE_PHN560_n3694;
   wire FE_PHN559_n1656;
   wire FE_PHN558_n3209;
   wire FE_PHN557_n4130;
   wire FE_PHN556_n2667;
   wire FE_PHN555_n4448;
   wire FE_PHN554_n2786;
   wire FE_PHN553_n3358;
   wire FE_PHN552_n802;
   wire FE_PHN551_n734;
   wire FE_PHN550_n3819;
   wire FE_PHN549_n4461;
   wire FE_PHN548_n3746;
   wire FE_PHN547_n3763;
   wire FE_PHN546_n793;
   wire FE_PHN545_n1790;
   wire FE_PHN544_n2183;
   wire FE_PHN543_n1690;
   wire FE_PHN542_n4553;
   wire FE_PHN541_n4044;
   wire FE_PHN540_n2942;
   wire FE_PHN539_n3881;
   wire FE_PHN538_n1735;
   wire FE_PHN537_n4622;
   wire FE_PHN536_n1611;
   wire FE_PHN535_n2839;
   wire FE_PHN534_n4118;
   wire FE_PHN533_n2744;
   wire FE_PHN532_n3329;
   wire FE_PHN531_n2354;
   wire FE_PHN530_n3742;
   wire FE_PHN529_n1957;
   wire FE_PHN528_n610;
   wire FE_PHN527_n1577;
   wire FE_PHN526_n2185;
   wire FE_PHN525_n2017;
   wire FE_PHN524_n2937;
   wire FE_PHN523_n1076;
   wire FE_PHN522_n2633;
   wire FE_PHN521_n3169;
   wire FE_PHN520_n3463;
   wire FE_PHN519_n1562;
   wire FE_PHN518_n4070;
   wire FE_PHN517_n3364;
   wire FE_PHN516_ram_29__14_;
   wire FE_PHN515_n3497;
   wire FE_PHN514_n3295;
   wire FE_PHN513_n4603;
   wire FE_PHN512_n736;
   wire FE_PHN511_n3838;
   wire FE_PHN510_n1443;
   wire FE_PHN509_n1055;
   wire FE_PHN508_n3323;
   wire FE_PHN507_n4441;
   wire FE_PHN506_n1700;
   wire FE_PHN505_n1816;
   wire FE_PHN504_n3337;
   wire FE_PHN503_n3676;
   wire FE_PHN502_n3327;
   wire FE_PHN501_n2456;
   wire FE_PHN500_n4275;
   wire FE_PHN499_n4609;
   wire FE_PHN498_n2948;
   wire FE_PHN497_n2915;
   wire FE_PHN496_n2718;
   wire FE_PHN495_n743;
   wire FE_PHN494_n4435;
   wire FE_PHN493_n4319;
   wire FE_PHN492_n4352;
   wire FE_PHN491_n1948;
   wire FE_PHN490_n2654;
   wire FE_PHN489_n3534;
   wire FE_PHN488_n3512;
   wire FE_PHN487_n3555;
   wire FE_PHN486_n3473;
   wire FE_PHN485_n4644;
   wire FE_PHN484_n3570;
   wire FE_PHN483_n3274;
   wire FE_PHN482_n3389;
   wire FE_PHN481_n4567;
   wire FE_PHN480_n1765;
   wire FE_PHN479_n2204;
   wire FE_PHN478_n4548;
   wire FE_PHN477_n2277;
   wire FE_PHN476_n2349;
   wire FE_PHN475_n2648;
   wire FE_PHN474_n4574;
   wire FE_PHN473_n2789;
   wire FE_PHN472_n3928;
   wire FE_PHN471_n4297;
   wire FE_PHN470_n1686;
   wire FE_PHN469_n4125;
   wire FE_PHN468_n1764;
   wire FE_PHN467_n2818;
   wire FE_PHN466_n3862;
   wire FE_PHN465_n769;
   wire FE_PHN464_n2254;
   wire FE_PHN463_n2765;
   wire FE_PHN462_n2348;
   wire FE_PHN461_n3842;
   wire FE_PHN460_n3912;
   wire FE_PHN459_n3375;
   wire FE_PHN458_n3877;
   wire FE_PHN457_n1137;
   wire FE_PHN456_n4129;
   wire FE_PHN455_n4493;
   wire FE_PHN454_n4282;
   wire FE_PHN453_n4632;
   wire FE_PHN452_n4589;
   wire FE_PHN451_n3798;
   wire FE_PHN450_n3362;
   wire FE_PHN449_n1059;
   wire FE_PHN448_n4565;
   wire FE_PHN447_n2714;
   wire FE_PHN446_n3579;
   wire FE_PHN445_n3810;
   wire FE_PHN444_n4602;
   wire FE_PHN443_n2711;
   wire FE_PHN442_n2205;
   wire FE_PHN441_n4527;
   wire FE_PHN440_n4503;
   wire FE_PHN439_n4106;
   wire FE_PHN438_n3633;
   wire FE_PHN437_n4508;
   wire FE_PHN436_n1406;
   wire FE_PHN435_n2071;
   wire FE_PHN434_n4471;
   wire FE_PHN433_n3888;
   wire FE_PHN432_n4512;
   wire FE_PHN431_n4054;
   wire FE_PHN430_n2236;
   wire FE_PHN429_n1644;
   wire FE_PHN428_n2365;
   wire FE_PHN427_n2531;
   wire FE_PHN426_n2637;
   wire FE_PHN425_n2274;
   wire FE_PHN424_n867;
   wire FE_PHN423_n990;
   wire FE_PHN422_n1710;
   wire FE_PHN421_n2356;
   wire FE_PHN420_n737;
   wire FE_PHN419_n3757;
   wire FE_PHN418_n2465;
   wire FE_PHN417_n1802;
   wire FE_PHN416_n862;
   wire FE_PHN415_n2299;
   wire FE_PHN414_n3156;
   wire FE_PHN413_n3625;
   wire FE_PHN412_n4566;
   wire FE_PHN411_n4635;
   wire FE_PHN410_n2032;
   wire FE_PHN409_n2361;
   wire FE_PHN408_n2435;
   wire FE_PHN407_n3670;
   wire FE_PHN406_n796;
   wire FE_PHN405_n3679;
   wire FE_PHN404_n1525;
   wire FE_PHN403_n3526;
   wire FE_PHN402_n1694;
   wire FE_PHN401_n804;
   wire FE_PHN400_n2245;
   wire FE_PHN399_n609;
   wire FE_PHN398_n2720;
   wire FE_PHN397_n1392;
   wire FE_PHN396_n1956;
   wire FE_PHN395_n2521;
   wire FE_PHN394_n4571;
   wire FE_PHN393_n1813;
   wire FE_PHN392_n2770;
   wire FE_PHN391_n2146;
   wire FE_PHN390_n3166;
   wire FE_PHN389_n1730;
   wire FE_PHN388_n1770;
   wire FE_PHN387_n4525;
   wire FE_PHN386_n4475;
   wire FE_PHN385_n2715;
   wire FE_PHN384_n2841;
   wire FE_PHN383_n3677;
   wire FE_PHN382_n3762;
   wire FE_PHN381_n3749;
   wire FE_PHN380_n1707;
   wire FE_PHN379_n3367;
   wire FE_PHN378_n1708;
   wire FE_PHN377_n1194;
   wire FE_PHN376_n601;
   wire FE_PHN375_n2337;
   wire FE_PHN374_n4246;
   wire FE_PHN373_n2779;
   wire FE_PHN372_n797;
   wire FE_PHN371_n4494;
   wire FE_PHN370_n3629;
   wire FE_PHN369_n4579;
   wire FE_PHN368_n4580;
   wire FE_PHN367_n4449;
   wire FE_PHN366_n4193;
   wire FE_PHN365_n987;
   wire FE_PHN364_n3236;
   wire FE_PHN363_n1509;
   wire FE_PHN362_n1711;
   wire FE_PHN361_n1065;
   wire FE_PHN360_n1330;
   wire FE_PHN359_n3531;
   wire FE_PHN358_n4326;
   wire FE_PHN357_n2473;
   wire FE_PHN356_n1653;
   wire FE_PHN355_n3354;
   wire FE_PHN354_n4581;
   wire FE_PHN353_n3608;
   wire FE_PHN352_n1063;
   wire FE_PHN351_n2647;
   wire FE_PHN350_n3805;
   wire FE_PHN349_n2294;
   wire FE_PHN348_n4474;
   wire FE_PHN347_n1792;
   wire FE_PHN346_n2801;
   wire FE_PHN345_n4257;
   wire FE_PHN344_n2787;
   wire FE_PHN343_n3165;
   wire FE_PHN342_n3233;
   wire FE_PHN341_n3743;
   wire FE_PHN340_n4038;
   wire FE_PHN339_n4613;
   wire FE_PHN338_n3783;
   wire FE_PHN337_n4318;
   wire FE_PHN336_n915;
   wire FE_PHN335_n1622;
   wire FE_PHN334_n2343;
   wire FE_PHN333_n3490;
   wire FE_PHN332_n3967;
   wire FE_PHN331_n3574;
   wire FE_PHN330_n2728;
   wire FE_PHN329_n3355;
   wire FE_PHN328_n3678;
   wire FE_PHN327_n3857;
   wire FE_PHN326_n4325;
   wire FE_PHN325_n3484;
   wire FE_PHN324_n3748;
   wire FE_PHN323_n3489;
   wire FE_PHN322_n1624;
   wire FE_PHN321_n2392;
   wire FE_PHN320_n4256;
   wire FE_PHN319_n3532;
   wire FE_PHN318_n1945;
   wire FE_PHN317_n4310;
   wire FE_PHN316_n1782;
   wire FE_PHN315_n3768;
   wire FE_PHN314_n3861;
   wire FE_PHN313_n4479;
   wire FE_PHN312_n4502;
   wire FE_PHN311_n1010;
   wire FE_PHN310_n2901;
   wire FE_PHN309_n4328;
   wire FE_PHN308_n2140;
   wire FE_PHN307_n2157;
   wire FE_PHN306_n2341;
   wire FE_PHN305_n3536;
   wire FE_PHN304_n3562;
   wire FE_PHN303_n2778;
   wire FE_PHN302_n4065;
   wire FE_PHN301_n3730;
   wire FE_PHN300_n4515;
   wire FE_PHN299_n2134;
   wire FE_PHN298_n1817;
   wire FE_PHN297_n2540;
   wire FE_PHN296_n3508;
   wire FE_PHN295_n4120;
   wire FE_PHN294_n1047;
   wire FE_PHN293_n2523;
   wire FE_PHN292_n2489;
   wire FE_PHN291_n4465;
   wire FE_PHN290_n1369;
   wire FE_PHN289_n3935;
   wire FE_PHN288_n4186;
   wire FE_PHN287_n4658;
   wire FE_PHN286_n3957;
   wire FE_PHN285_n2200;
   wire FE_PHN284_n2601;
   wire FE_PHN283_n4633;
   wire FE_PHN282_n3557;
   wire FE_PHN281_n4568;
   wire FE_PHN280_n3380;
   wire FE_PHN279_n2162;
   wire FE_PHN278_n3097;
   wire FE_PHN277_n1626;
   wire FE_PHN276_n3544;
   wire FE_PHN275_n1753;
   wire FE_PHN274_n2796;
   wire FE_PHN273_n4081;
   wire FE_PHN272_n4533;
   wire FE_PHN271_n2278;
   wire FE_PHN270_n2467;
   wire FE_PHN269_n2340;
   wire FE_PHN268_n1061;
   wire FE_PHN267_n1373;
   wire FE_PHN266_n3611;
   wire FE_PHN265_n3772;
   wire FE_PHN264_n2409;
   wire FE_PHN263_n4477;
   wire FE_PHN262_n3350;
   wire FE_PHN261_n2201;
   wire FE_PHN260_n2761;
   wire FE_PHN259_n1508;
   wire FE_PHN258_n1814;
   wire FE_PHN257_n3817;
   wire FE_PHN256_n1146;
   wire FE_PHN255_n1781;
   wire FE_PHN254_n3231;
   wire FE_PHN253_n3986;
   wire FE_PHN252_n2455;
   wire FE_PHN251_n1691;
   wire FE_PHN250_n4024;
   wire FE_PHN249_n2461;
   wire FE_PHN248_n3747;
   wire FE_PHN247_n2652;
   wire FE_PHN246_n3172;
   wire FE_PHN245_n763;
   wire FE_PHN244_n2588;
   wire FE_PHN243_n1795;
   wire FE_PHN242_n2174;
   wire FE_PHN241_n2741;
   wire FE_PHN240_n4247;
   wire FE_PHN239_n4105;
   wire FE_PHN238_n3572;
   wire FE_PHN237_n4317;
   wire FE_PHN236_n3863;
   wire FE_PHN235_n1761;
   wire FE_PHN234_n4191;
   wire FE_PHN233_n4092;
   wire FE_PHN232_n791;
   wire FE_PHN231_n3991;
   wire FE_PHN230_n3543;
   wire FE_PHN229_n2333;
   wire FE_PHN228_n3632;
   wire FE_PHN227_n4600;
   wire FE_PHN226_n1239;
   wire FE_PHN225_n2212;
   wire FE_PHN224_n3735;
   wire FE_PHN223_n4020;
   wire FE_PHN222_n2803;
   wire FE_PHN221_n2651;
   wire FE_PHN220_n4636;
   wire FE_PHN219_n2805;
   wire FE_PHN218_n3610;
   wire FE_PHN217_n3239;
   wire FE_PHN216_n2266;
   wire FE_PHN215_n3997;
   wire FE_PHN214_n3565;
   wire FE_PHN213_n3170;
   wire FE_PHN212_n4426;
   wire FE_PHN211_n1121;
   wire FE_PHN210_n4132;
   wire FE_PHN209_n3938;
   wire FE_PHN208_n3744;
   wire FE_PHN207_n3673;
   wire FE_PHN206_n1818;
   wire FE_PHN205_n3352;
   wire FE_PHN204_n1754;
   wire FE_PHN203_n1701;
   wire FE_PHN202_n2338;
   wire FE_PHN201_n3990;
   wire FE_PHN200_n4288;
   wire FE_PHN199_n3101;
   wire FE_PHN198_n2208;
   wire FE_PHN197_n4315;
   wire FE_PHN196_n3905;
   wire FE_PHN195_n4587;
   wire FE_PHN194_n2476;
   wire FE_PHN193_n3493;
   wire FE_PHN192_n735;
   wire FE_PHN191_n3682;
   wire FE_PHN190_n4182;
   wire FE_PHN189_n2712;
   wire FE_PHN188_n3213;
   wire FE_PHN187_n4084;
   wire FE_PHN186_n4320;
   wire FE_PHN185_n4376;
   wire FE_PHN184_n1696;
   wire FE_PHN183_n3491;
   wire FE_PHN182_n1053;
   wire FE_PHN181_n3292;
   wire FE_PHN180_n4456;
   wire FE_PHN179_n3754;
   wire FE_PHN178_n3353;
   wire FE_PHN177_n3300;
   wire FE_PHN176_n1112;
   wire FE_PHN175_n3167;
   wire FE_PHN174_n3734;
   wire FE_PHN173_n4004;
   wire FE_PHN172_n4570;
   wire FE_PHN171_n4190;
   wire FE_PHN170_n3561;
   wire FE_PHN169_n4582;
   wire FE_PHN168_n1435;
   wire FE_PHN167_n3580;
   wire FE_PHN166_n4514;
   wire FE_PHN165_ram_241__1_;
   wire FE_PHN164_n3164;
   wire FE_PHN163_n2458;
   wire FE_PHN162_n3234;
   wire FE_PHN161_n3548;
   wire FE_PHN160_n3618;
   wire FE_PHN159_n3224;
   wire FE_PHN158_n3563;
   wire FE_PHN157_n3286;
   wire FE_PHN156_n3499;
   wire FE_PHN155_n4055;
   wire FE_PHN154_n3365;
   wire FE_PHN153_n3550;
   wire FE_PHN152_n1049;
   wire FE_PHN151_n1572;
   wire FE_PHN150_n3564;
   wire FE_PHN149_n3621;
   wire FE_PHN148_n4522;
   wire FE_PHN147_n3556;
   wire FE_PHN146_n3609;
   wire FE_PHN145_n2330;
   wire FE_PHN144_n1634;
   wire FE_PHN143_n1704;
   wire FE_PHN142_n3864;
   wire FE_PHN141_n2206;
   wire FE_PHN140_n4313;
   wire FE_PHN139_n4506;
   wire FE_PHN138_n1713;
   wire FE_PHN137_n2142;
   wire FE_PHN136_n4573;
   wire FE_PHN135_n4064;
   wire FE_PHN134_n3606;
   wire FE_PHN133_n2136;
   wire FE_PHN132_n3106;
   wire FE_PHN131_n3870;
   wire FE_PHN130_n4068;
   wire FE_PHN129_n2147;
   wire FE_PHN128_n1695;
   wire FE_PHN127_n4507;
   wire FE_PHN126_n3866;
   wire FE_PHN125_n3546;
   wire FE_PHN124_n2273;
   wire FE_PHN123_n1058;
   wire FE_PHN122_n3226;
   wire FE_PHN121_n3995;
   wire FE_PHN120_n4509;
   wire FE_PHN119_n3538;
   wire FE_PHN118_n4446;
   wire FE_PHN117_n3301;
   wire FE_PHN116_n2207;
   wire FE_PHN115_n3739;
   wire FE_PHN114_n3807;
   wire FE_PHN113_n3533;
   wire FE_PHN112_n4577;
   wire FE_PHN111_n3584;
   wire FE_PHN110_n4504;
   wire FE_PHN109_n3549;
   wire FE_PHN108_n3568;
   wire FE_PHN107_n1692;
   wire FE_PHN106_n3619;
   wire FE_PHN105_n3552;
   wire FE_PHN104_n3545;
   wire FE_PHN103_n3558;
   wire FE_PHN102_n3554;
   wire FE_PHN101_n3547;
   wire FE_PHN100_n3542;
   wire FE_OFN94_mem_write;
   wire FE_OFN93_mem_write;
   wire FE_OFN92_mem_write;
   wire FE_OFN91_n23;
   wire FE_OFN90_n23;
   wire FE_OFN89_n23;
   wire FE_OFN88_n22;
   wire FE_OFN87_n22;
   wire FE_OFN86_n22;
   wire FE_OFN85_n21;
   wire FE_OFN84_n21;
   wire FE_OFN83_n21;
   wire FE_OFN82_n20;
   wire FE_OFN81_n20;
   wire FE_OFN80_n20;
   wire FE_OFN79_n20;
   wire FE_OFN78_n19;
   wire FE_OFN77_n19;
   wire FE_OFN76_n19;
   wire FE_OFN75_n18;
   wire FE_OFN74_n18;
   wire FE_OFN73_n18;
   wire FE_OFN72_n17;
   wire FE_OFN71_n17;
   wire FE_OFN70_n17;
   wire FE_OFN69_n16;
   wire FE_OFN68_n16;
   wire FE_OFN67_n16;
   wire FE_OFN66_n16;
   wire FE_OFN65_n15;
   wire FE_OFN64_n15;
   wire FE_OFN63_n15;
   wire FE_OFN62_n14;
   wire FE_OFN61_n14;
   wire FE_OFN60_n14;
   wire FE_OFN59_n14;
   wire FE_OFN58_n13;
   wire FE_OFN57_n13;
   wire FE_OFN56_n13;
   wire FE_OFN55_n12;
   wire FE_OFN54_n12;
   wire FE_OFN53_n12;
   wire FE_OFN52_n11;
   wire FE_OFN51_n11;
   wire FE_OFN50_n11;
   wire FE_OFN49_n10;
   wire FE_OFN48_n10;
   wire FE_OFN47_n10;
   wire FE_OFN46_n9;
   wire FE_OFN45_n9;
   wire FE_OFN44_n9;
   wire FE_OFN43_n6;
   wire FE_OFN42_n6;
   wire FE_OFN41_n6;
   wire FE_OFN40_n6459;
   wire FE_OFN39_n6459;
   wire FE_OFN38_n6459;
   wire FE_OFN37_n6459;
   wire FE_OFN36_n6459;
   wire FE_OFN35_n6459;
   wire FE_OFN34_n6459;
   wire FE_OFN33_n6459;
   wire FE_OFN32_n6459;
   wire FE_OFN31_n6459;
   wire FE_OFN30_n6459;
   wire FE_OFN29_n6459;
   wire FE_OFN28_n6459;
   wire FE_OFN27_n6459;
   wire FE_OFN26_n6459;
   wire FE_OFN25_n6459;
   wire FE_OFN24_n6136;
   wire FE_OFN23_n6136;
   wire FE_OFN22_n6136;
   wire FE_OFN21_n7440;
   wire FE_OFN20_n7440;
   wire FE_OFN19_n7440;
   wire FE_OFN18_n7440;
   wire FE_OFN17_n7440;
   wire FE_OFN16_n7440;
   wire FE_OFN15_n7440;
   wire FE_OFN14_n7440;
   wire FE_OFN13_n7440;
   wire FE_OFN12_n7440;
   wire FE_OFN11_n7440;
   wire FE_OFN10_n7440;
   wire FE_OFN9_n7440;
   wire FE_OFN8_n7440;
   wire FE_OFN7_n7440;
   wire FE_OFN6_n7440;
   wire FE_OFN5_n7440;
   wire FE_OFN4_n7442;
   wire FE_OFN3_n7442;
   wire FE_OFN2_n7442;
   wire FE_OFN1_n7442;
   wire FE_OFN0_n7442;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire \ram[255][15] ;
   wire \ram[255][14] ;
   wire \ram[255][13] ;
   wire \ram[255][12] ;
   wire \ram[255][11] ;
   wire \ram[255][10] ;
   wire \ram[255][9] ;
   wire \ram[255][8] ;
   wire \ram[255][7] ;
   wire \ram[255][6] ;
   wire \ram[255][5] ;
   wire \ram[255][4] ;
   wire \ram[255][3] ;
   wire \ram[255][2] ;
   wire \ram[255][1] ;
   wire \ram[255][0] ;
   wire \ram[254][15] ;
   wire \ram[254][14] ;
   wire \ram[254][13] ;
   wire \ram[254][12] ;
   wire \ram[254][11] ;
   wire \ram[254][10] ;
   wire \ram[254][9] ;
   wire \ram[254][8] ;
   wire \ram[254][7] ;
   wire \ram[254][6] ;
   wire \ram[254][5] ;
   wire \ram[254][4] ;
   wire \ram[254][3] ;
   wire \ram[254][2] ;
   wire \ram[254][1] ;
   wire \ram[254][0] ;
   wire \ram[253][15] ;
   wire \ram[253][14] ;
   wire \ram[253][13] ;
   wire \ram[253][12] ;
   wire \ram[253][11] ;
   wire \ram[253][10] ;
   wire \ram[253][9] ;
   wire \ram[253][8] ;
   wire \ram[253][7] ;
   wire \ram[253][6] ;
   wire \ram[253][5] ;
   wire \ram[253][4] ;
   wire \ram[253][3] ;
   wire \ram[253][2] ;
   wire \ram[253][1] ;
   wire \ram[253][0] ;
   wire \ram[252][15] ;
   wire \ram[252][14] ;
   wire \ram[252][13] ;
   wire \ram[252][12] ;
   wire \ram[252][11] ;
   wire \ram[252][10] ;
   wire \ram[252][9] ;
   wire \ram[252][8] ;
   wire \ram[252][7] ;
   wire \ram[252][6] ;
   wire \ram[252][5] ;
   wire \ram[252][4] ;
   wire \ram[252][3] ;
   wire \ram[252][2] ;
   wire \ram[252][1] ;
   wire \ram[252][0] ;
   wire \ram[251][15] ;
   wire \ram[251][14] ;
   wire \ram[251][13] ;
   wire \ram[251][12] ;
   wire \ram[251][11] ;
   wire \ram[251][10] ;
   wire \ram[251][9] ;
   wire \ram[251][8] ;
   wire \ram[251][7] ;
   wire \ram[251][6] ;
   wire \ram[251][5] ;
   wire \ram[251][4] ;
   wire \ram[251][3] ;
   wire \ram[251][2] ;
   wire \ram[251][1] ;
   wire \ram[251][0] ;
   wire \ram[250][15] ;
   wire \ram[250][14] ;
   wire \ram[250][13] ;
   wire \ram[250][12] ;
   wire \ram[250][11] ;
   wire \ram[250][10] ;
   wire \ram[250][9] ;
   wire \ram[250][8] ;
   wire \ram[250][7] ;
   wire \ram[250][6] ;
   wire \ram[250][5] ;
   wire \ram[250][4] ;
   wire \ram[250][3] ;
   wire \ram[250][2] ;
   wire \ram[250][1] ;
   wire \ram[250][0] ;
   wire \ram[249][15] ;
   wire \ram[249][14] ;
   wire \ram[249][13] ;
   wire \ram[249][12] ;
   wire \ram[249][11] ;
   wire \ram[249][10] ;
   wire \ram[249][9] ;
   wire \ram[249][8] ;
   wire \ram[249][7] ;
   wire \ram[249][6] ;
   wire \ram[249][5] ;
   wire \ram[249][4] ;
   wire \ram[249][3] ;
   wire \ram[249][2] ;
   wire \ram[249][1] ;
   wire \ram[249][0] ;
   wire \ram[248][15] ;
   wire \ram[248][14] ;
   wire \ram[248][13] ;
   wire \ram[248][12] ;
   wire \ram[248][11] ;
   wire \ram[248][10] ;
   wire \ram[248][9] ;
   wire \ram[248][8] ;
   wire \ram[248][7] ;
   wire \ram[248][6] ;
   wire \ram[248][5] ;
   wire \ram[248][4] ;
   wire \ram[248][3] ;
   wire \ram[248][2] ;
   wire \ram[248][1] ;
   wire \ram[248][0] ;
   wire \ram[247][15] ;
   wire \ram[247][14] ;
   wire \ram[247][13] ;
   wire \ram[247][12] ;
   wire \ram[247][11] ;
   wire \ram[247][10] ;
   wire \ram[247][9] ;
   wire \ram[247][8] ;
   wire \ram[247][7] ;
   wire \ram[247][6] ;
   wire \ram[247][5] ;
   wire \ram[247][4] ;
   wire \ram[247][3] ;
   wire \ram[247][2] ;
   wire \ram[247][1] ;
   wire \ram[247][0] ;
   wire \ram[246][15] ;
   wire \ram[246][14] ;
   wire \ram[246][13] ;
   wire \ram[246][12] ;
   wire \ram[246][11] ;
   wire \ram[246][10] ;
   wire \ram[246][9] ;
   wire \ram[246][8] ;
   wire \ram[246][7] ;
   wire \ram[246][6] ;
   wire \ram[246][5] ;
   wire \ram[246][4] ;
   wire \ram[246][3] ;
   wire \ram[246][2] ;
   wire \ram[246][1] ;
   wire \ram[246][0] ;
   wire \ram[245][15] ;
   wire \ram[245][14] ;
   wire \ram[245][13] ;
   wire \ram[245][12] ;
   wire \ram[245][11] ;
   wire \ram[245][10] ;
   wire \ram[245][9] ;
   wire \ram[245][8] ;
   wire \ram[245][7] ;
   wire \ram[245][6] ;
   wire \ram[245][5] ;
   wire \ram[245][4] ;
   wire \ram[245][3] ;
   wire \ram[245][2] ;
   wire \ram[245][1] ;
   wire \ram[245][0] ;
   wire \ram[244][15] ;
   wire \ram[244][14] ;
   wire \ram[244][13] ;
   wire \ram[244][12] ;
   wire \ram[244][11] ;
   wire \ram[244][10] ;
   wire \ram[244][9] ;
   wire \ram[244][8] ;
   wire \ram[244][7] ;
   wire \ram[244][6] ;
   wire \ram[244][5] ;
   wire \ram[244][4] ;
   wire \ram[244][3] ;
   wire \ram[244][2] ;
   wire \ram[244][1] ;
   wire \ram[244][0] ;
   wire \ram[243][15] ;
   wire \ram[243][14] ;
   wire \ram[243][13] ;
   wire \ram[243][12] ;
   wire \ram[243][11] ;
   wire \ram[243][10] ;
   wire \ram[243][9] ;
   wire \ram[243][8] ;
   wire \ram[243][7] ;
   wire \ram[243][6] ;
   wire \ram[243][5] ;
   wire \ram[243][4] ;
   wire \ram[243][3] ;
   wire \ram[243][2] ;
   wire \ram[243][1] ;
   wire \ram[243][0] ;
   wire \ram[242][15] ;
   wire \ram[242][14] ;
   wire \ram[242][13] ;
   wire \ram[242][12] ;
   wire \ram[242][11] ;
   wire \ram[242][10] ;
   wire \ram[242][9] ;
   wire \ram[242][8] ;
   wire \ram[242][7] ;
   wire \ram[242][6] ;
   wire \ram[242][5] ;
   wire \ram[242][4] ;
   wire \ram[242][3] ;
   wire \ram[242][2] ;
   wire \ram[242][1] ;
   wire \ram[242][0] ;
   wire \ram[241][15] ;
   wire \ram[241][14] ;
   wire \ram[241][13] ;
   wire \ram[241][12] ;
   wire \ram[241][11] ;
   wire \ram[241][10] ;
   wire \ram[241][9] ;
   wire \ram[241][8] ;
   wire \ram[241][7] ;
   wire \ram[241][6] ;
   wire \ram[241][5] ;
   wire \ram[241][4] ;
   wire \ram[241][3] ;
   wire \ram[241][2] ;
   wire \ram[241][1] ;
   wire \ram[241][0] ;
   wire \ram[240][15] ;
   wire \ram[240][14] ;
   wire \ram[240][13] ;
   wire \ram[240][12] ;
   wire \ram[240][11] ;
   wire \ram[240][10] ;
   wire \ram[240][9] ;
   wire \ram[240][8] ;
   wire \ram[240][7] ;
   wire \ram[240][6] ;
   wire \ram[240][5] ;
   wire \ram[240][4] ;
   wire \ram[240][3] ;
   wire \ram[240][2] ;
   wire \ram[240][1] ;
   wire \ram[240][0] ;
   wire \ram[239][15] ;
   wire \ram[239][14] ;
   wire \ram[239][13] ;
   wire \ram[239][12] ;
   wire \ram[239][11] ;
   wire \ram[239][10] ;
   wire \ram[239][9] ;
   wire \ram[239][8] ;
   wire \ram[239][7] ;
   wire \ram[239][6] ;
   wire \ram[239][5] ;
   wire \ram[239][4] ;
   wire \ram[239][3] ;
   wire \ram[239][2] ;
   wire \ram[239][1] ;
   wire \ram[239][0] ;
   wire \ram[238][15] ;
   wire \ram[238][14] ;
   wire \ram[238][13] ;
   wire \ram[238][12] ;
   wire \ram[238][11] ;
   wire \ram[238][10] ;
   wire \ram[238][9] ;
   wire \ram[238][8] ;
   wire \ram[238][7] ;
   wire \ram[238][6] ;
   wire \ram[238][5] ;
   wire \ram[238][4] ;
   wire \ram[238][3] ;
   wire \ram[238][2] ;
   wire \ram[238][1] ;
   wire \ram[238][0] ;
   wire \ram[237][15] ;
   wire \ram[237][14] ;
   wire \ram[237][13] ;
   wire \ram[237][12] ;
   wire \ram[237][11] ;
   wire \ram[237][10] ;
   wire \ram[237][9] ;
   wire \ram[237][8] ;
   wire \ram[237][7] ;
   wire \ram[237][6] ;
   wire \ram[237][5] ;
   wire \ram[237][4] ;
   wire \ram[237][3] ;
   wire \ram[237][2] ;
   wire \ram[237][1] ;
   wire \ram[237][0] ;
   wire \ram[236][15] ;
   wire \ram[236][14] ;
   wire \ram[236][13] ;
   wire \ram[236][12] ;
   wire \ram[236][11] ;
   wire \ram[236][10] ;
   wire \ram[236][9] ;
   wire \ram[236][8] ;
   wire \ram[236][7] ;
   wire \ram[236][6] ;
   wire \ram[236][5] ;
   wire \ram[236][4] ;
   wire \ram[236][3] ;
   wire \ram[236][2] ;
   wire \ram[236][1] ;
   wire \ram[236][0] ;
   wire \ram[235][15] ;
   wire \ram[235][14] ;
   wire \ram[235][13] ;
   wire \ram[235][12] ;
   wire \ram[235][11] ;
   wire \ram[235][10] ;
   wire \ram[235][9] ;
   wire \ram[235][8] ;
   wire \ram[235][7] ;
   wire \ram[235][6] ;
   wire \ram[235][5] ;
   wire \ram[235][4] ;
   wire \ram[235][3] ;
   wire \ram[235][2] ;
   wire \ram[235][1] ;
   wire \ram[235][0] ;
   wire \ram[234][15] ;
   wire \ram[234][14] ;
   wire \ram[234][13] ;
   wire \ram[234][12] ;
   wire \ram[234][11] ;
   wire \ram[234][10] ;
   wire \ram[234][9] ;
   wire \ram[234][8] ;
   wire \ram[234][7] ;
   wire \ram[234][6] ;
   wire \ram[234][5] ;
   wire \ram[234][4] ;
   wire \ram[234][3] ;
   wire \ram[234][2] ;
   wire \ram[234][1] ;
   wire \ram[234][0] ;
   wire \ram[233][15] ;
   wire \ram[233][14] ;
   wire \ram[233][13] ;
   wire \ram[233][12] ;
   wire \ram[233][11] ;
   wire \ram[233][10] ;
   wire \ram[233][9] ;
   wire \ram[233][8] ;
   wire \ram[233][7] ;
   wire \ram[233][6] ;
   wire \ram[233][5] ;
   wire \ram[233][4] ;
   wire \ram[233][3] ;
   wire \ram[233][2] ;
   wire \ram[233][1] ;
   wire \ram[233][0] ;
   wire \ram[232][15] ;
   wire \ram[232][14] ;
   wire \ram[232][13] ;
   wire \ram[232][12] ;
   wire \ram[232][11] ;
   wire \ram[232][10] ;
   wire \ram[232][9] ;
   wire \ram[232][8] ;
   wire \ram[232][7] ;
   wire \ram[232][6] ;
   wire \ram[232][5] ;
   wire \ram[232][4] ;
   wire \ram[232][3] ;
   wire \ram[232][2] ;
   wire \ram[232][1] ;
   wire \ram[232][0] ;
   wire \ram[231][15] ;
   wire \ram[231][14] ;
   wire \ram[231][13] ;
   wire \ram[231][12] ;
   wire \ram[231][11] ;
   wire \ram[231][10] ;
   wire \ram[231][9] ;
   wire \ram[231][8] ;
   wire \ram[231][7] ;
   wire \ram[231][6] ;
   wire \ram[231][5] ;
   wire \ram[231][4] ;
   wire \ram[231][3] ;
   wire \ram[231][2] ;
   wire \ram[231][1] ;
   wire \ram[231][0] ;
   wire \ram[230][15] ;
   wire \ram[230][14] ;
   wire \ram[230][13] ;
   wire \ram[230][12] ;
   wire \ram[230][11] ;
   wire \ram[230][10] ;
   wire \ram[230][9] ;
   wire \ram[230][8] ;
   wire \ram[230][7] ;
   wire \ram[230][6] ;
   wire \ram[230][5] ;
   wire \ram[230][4] ;
   wire \ram[230][3] ;
   wire \ram[230][2] ;
   wire \ram[230][1] ;
   wire \ram[230][0] ;
   wire \ram[229][15] ;
   wire \ram[229][14] ;
   wire \ram[229][13] ;
   wire \ram[229][12] ;
   wire \ram[229][11] ;
   wire \ram[229][10] ;
   wire \ram[229][9] ;
   wire \ram[229][8] ;
   wire \ram[229][7] ;
   wire \ram[229][6] ;
   wire \ram[229][5] ;
   wire \ram[229][4] ;
   wire \ram[229][3] ;
   wire \ram[229][2] ;
   wire \ram[229][1] ;
   wire \ram[229][0] ;
   wire \ram[228][15] ;
   wire \ram[228][14] ;
   wire \ram[228][13] ;
   wire \ram[228][12] ;
   wire \ram[228][11] ;
   wire \ram[228][10] ;
   wire \ram[228][9] ;
   wire \ram[228][8] ;
   wire \ram[228][7] ;
   wire \ram[228][6] ;
   wire \ram[228][5] ;
   wire \ram[228][4] ;
   wire \ram[228][3] ;
   wire \ram[228][2] ;
   wire \ram[228][1] ;
   wire \ram[228][0] ;
   wire \ram[227][15] ;
   wire \ram[227][14] ;
   wire \ram[227][13] ;
   wire \ram[227][12] ;
   wire \ram[227][11] ;
   wire \ram[227][10] ;
   wire \ram[227][9] ;
   wire \ram[227][8] ;
   wire \ram[227][7] ;
   wire \ram[227][6] ;
   wire \ram[227][5] ;
   wire \ram[227][4] ;
   wire \ram[227][3] ;
   wire \ram[227][2] ;
   wire \ram[227][1] ;
   wire \ram[227][0] ;
   wire \ram[226][15] ;
   wire \ram[226][14] ;
   wire \ram[226][13] ;
   wire \ram[226][12] ;
   wire \ram[226][11] ;
   wire \ram[226][10] ;
   wire \ram[226][9] ;
   wire \ram[226][8] ;
   wire \ram[226][7] ;
   wire \ram[226][6] ;
   wire \ram[226][5] ;
   wire \ram[226][4] ;
   wire \ram[226][3] ;
   wire \ram[226][2] ;
   wire \ram[226][1] ;
   wire \ram[226][0] ;
   wire \ram[225][15] ;
   wire \ram[225][14] ;
   wire \ram[225][13] ;
   wire \ram[225][12] ;
   wire \ram[225][11] ;
   wire \ram[225][10] ;
   wire \ram[225][9] ;
   wire \ram[225][8] ;
   wire \ram[225][7] ;
   wire \ram[225][6] ;
   wire \ram[225][5] ;
   wire \ram[225][4] ;
   wire \ram[225][3] ;
   wire \ram[225][2] ;
   wire \ram[225][1] ;
   wire \ram[225][0] ;
   wire \ram[224][15] ;
   wire \ram[224][14] ;
   wire \ram[224][13] ;
   wire \ram[224][12] ;
   wire \ram[224][11] ;
   wire \ram[224][10] ;
   wire \ram[224][9] ;
   wire \ram[224][8] ;
   wire \ram[224][7] ;
   wire \ram[224][6] ;
   wire \ram[224][5] ;
   wire \ram[224][4] ;
   wire \ram[224][3] ;
   wire \ram[224][2] ;
   wire \ram[224][1] ;
   wire \ram[224][0] ;
   wire \ram[223][15] ;
   wire \ram[223][14] ;
   wire \ram[223][13] ;
   wire \ram[223][12] ;
   wire \ram[223][11] ;
   wire \ram[223][10] ;
   wire \ram[223][9] ;
   wire \ram[223][8] ;
   wire \ram[223][7] ;
   wire \ram[223][6] ;
   wire \ram[223][5] ;
   wire \ram[223][4] ;
   wire \ram[223][3] ;
   wire \ram[223][2] ;
   wire \ram[223][1] ;
   wire \ram[223][0] ;
   wire \ram[222][15] ;
   wire \ram[222][14] ;
   wire \ram[222][13] ;
   wire \ram[222][12] ;
   wire \ram[222][11] ;
   wire \ram[222][10] ;
   wire \ram[222][9] ;
   wire \ram[222][8] ;
   wire \ram[222][7] ;
   wire \ram[222][6] ;
   wire \ram[222][5] ;
   wire \ram[222][4] ;
   wire \ram[222][3] ;
   wire \ram[222][2] ;
   wire \ram[222][1] ;
   wire \ram[222][0] ;
   wire \ram[221][15] ;
   wire \ram[221][14] ;
   wire \ram[221][13] ;
   wire \ram[221][12] ;
   wire \ram[221][11] ;
   wire \ram[221][10] ;
   wire \ram[221][9] ;
   wire \ram[221][8] ;
   wire \ram[221][7] ;
   wire \ram[221][6] ;
   wire \ram[221][5] ;
   wire \ram[221][4] ;
   wire \ram[221][3] ;
   wire \ram[221][2] ;
   wire \ram[221][1] ;
   wire \ram[221][0] ;
   wire \ram[220][15] ;
   wire \ram[220][14] ;
   wire \ram[220][13] ;
   wire \ram[220][12] ;
   wire \ram[220][11] ;
   wire \ram[220][10] ;
   wire \ram[220][9] ;
   wire \ram[220][8] ;
   wire \ram[220][7] ;
   wire \ram[220][6] ;
   wire \ram[220][5] ;
   wire \ram[220][4] ;
   wire \ram[220][3] ;
   wire \ram[220][2] ;
   wire \ram[220][1] ;
   wire \ram[220][0] ;
   wire \ram[219][15] ;
   wire \ram[219][14] ;
   wire \ram[219][13] ;
   wire \ram[219][12] ;
   wire \ram[219][11] ;
   wire \ram[219][10] ;
   wire \ram[219][9] ;
   wire \ram[219][8] ;
   wire \ram[219][7] ;
   wire \ram[219][6] ;
   wire \ram[219][5] ;
   wire \ram[219][4] ;
   wire \ram[219][3] ;
   wire \ram[219][2] ;
   wire \ram[219][1] ;
   wire \ram[219][0] ;
   wire \ram[218][15] ;
   wire \ram[218][14] ;
   wire \ram[218][13] ;
   wire \ram[218][12] ;
   wire \ram[218][11] ;
   wire \ram[218][10] ;
   wire \ram[218][9] ;
   wire \ram[218][8] ;
   wire \ram[218][7] ;
   wire \ram[218][6] ;
   wire \ram[218][5] ;
   wire \ram[218][4] ;
   wire \ram[218][3] ;
   wire \ram[218][2] ;
   wire \ram[218][1] ;
   wire \ram[218][0] ;
   wire \ram[217][15] ;
   wire \ram[217][14] ;
   wire \ram[217][13] ;
   wire \ram[217][12] ;
   wire \ram[217][11] ;
   wire \ram[217][10] ;
   wire \ram[217][9] ;
   wire \ram[217][8] ;
   wire \ram[217][7] ;
   wire \ram[217][6] ;
   wire \ram[217][5] ;
   wire \ram[217][4] ;
   wire \ram[217][3] ;
   wire \ram[217][2] ;
   wire \ram[217][1] ;
   wire \ram[217][0] ;
   wire \ram[216][15] ;
   wire \ram[216][14] ;
   wire \ram[216][13] ;
   wire \ram[216][12] ;
   wire \ram[216][11] ;
   wire \ram[216][10] ;
   wire \ram[216][9] ;
   wire \ram[216][8] ;
   wire \ram[216][7] ;
   wire \ram[216][6] ;
   wire \ram[216][5] ;
   wire \ram[216][4] ;
   wire \ram[216][3] ;
   wire \ram[216][2] ;
   wire \ram[216][1] ;
   wire \ram[216][0] ;
   wire \ram[215][15] ;
   wire \ram[215][14] ;
   wire \ram[215][13] ;
   wire \ram[215][12] ;
   wire \ram[215][11] ;
   wire \ram[215][10] ;
   wire \ram[215][9] ;
   wire \ram[215][8] ;
   wire \ram[215][7] ;
   wire \ram[215][6] ;
   wire \ram[215][5] ;
   wire \ram[215][4] ;
   wire \ram[215][3] ;
   wire \ram[215][2] ;
   wire \ram[215][1] ;
   wire \ram[215][0] ;
   wire \ram[214][15] ;
   wire \ram[214][14] ;
   wire \ram[214][13] ;
   wire \ram[214][12] ;
   wire \ram[214][11] ;
   wire \ram[214][10] ;
   wire \ram[214][9] ;
   wire \ram[214][8] ;
   wire \ram[214][7] ;
   wire \ram[214][6] ;
   wire \ram[214][5] ;
   wire \ram[214][4] ;
   wire \ram[214][3] ;
   wire \ram[214][2] ;
   wire \ram[214][1] ;
   wire \ram[214][0] ;
   wire \ram[213][15] ;
   wire \ram[213][14] ;
   wire \ram[213][13] ;
   wire \ram[213][12] ;
   wire \ram[213][11] ;
   wire \ram[213][10] ;
   wire \ram[213][9] ;
   wire \ram[213][8] ;
   wire \ram[213][7] ;
   wire \ram[213][6] ;
   wire \ram[213][5] ;
   wire \ram[213][4] ;
   wire \ram[213][3] ;
   wire \ram[213][2] ;
   wire \ram[213][1] ;
   wire \ram[213][0] ;
   wire \ram[212][15] ;
   wire \ram[212][14] ;
   wire \ram[212][13] ;
   wire \ram[212][12] ;
   wire \ram[212][11] ;
   wire \ram[212][10] ;
   wire \ram[212][9] ;
   wire \ram[212][8] ;
   wire \ram[212][7] ;
   wire \ram[212][6] ;
   wire \ram[212][5] ;
   wire \ram[212][4] ;
   wire \ram[212][3] ;
   wire \ram[212][2] ;
   wire \ram[212][1] ;
   wire \ram[212][0] ;
   wire \ram[211][15] ;
   wire \ram[211][14] ;
   wire \ram[211][13] ;
   wire \ram[211][12] ;
   wire \ram[211][11] ;
   wire \ram[211][10] ;
   wire \ram[211][9] ;
   wire \ram[211][8] ;
   wire \ram[211][7] ;
   wire \ram[211][6] ;
   wire \ram[211][5] ;
   wire \ram[211][4] ;
   wire \ram[211][3] ;
   wire \ram[211][2] ;
   wire \ram[211][1] ;
   wire \ram[211][0] ;
   wire \ram[210][15] ;
   wire \ram[210][14] ;
   wire \ram[210][13] ;
   wire \ram[210][12] ;
   wire \ram[210][11] ;
   wire \ram[210][10] ;
   wire \ram[210][9] ;
   wire \ram[210][8] ;
   wire \ram[210][7] ;
   wire \ram[210][6] ;
   wire \ram[210][5] ;
   wire \ram[210][4] ;
   wire \ram[210][3] ;
   wire \ram[210][2] ;
   wire \ram[210][1] ;
   wire \ram[210][0] ;
   wire \ram[209][15] ;
   wire \ram[209][14] ;
   wire \ram[209][13] ;
   wire \ram[209][12] ;
   wire \ram[209][11] ;
   wire \ram[209][10] ;
   wire \ram[209][9] ;
   wire \ram[209][8] ;
   wire \ram[209][7] ;
   wire \ram[209][6] ;
   wire \ram[209][5] ;
   wire \ram[209][4] ;
   wire \ram[209][3] ;
   wire \ram[209][2] ;
   wire \ram[209][1] ;
   wire \ram[209][0] ;
   wire \ram[208][15] ;
   wire \ram[208][14] ;
   wire \ram[208][13] ;
   wire \ram[208][12] ;
   wire \ram[208][11] ;
   wire \ram[208][10] ;
   wire \ram[208][9] ;
   wire \ram[208][8] ;
   wire \ram[208][7] ;
   wire \ram[208][6] ;
   wire \ram[208][5] ;
   wire \ram[208][4] ;
   wire \ram[208][3] ;
   wire \ram[208][2] ;
   wire \ram[208][1] ;
   wire \ram[208][0] ;
   wire \ram[207][15] ;
   wire \ram[207][14] ;
   wire \ram[207][13] ;
   wire \ram[207][12] ;
   wire \ram[207][11] ;
   wire \ram[207][10] ;
   wire \ram[207][9] ;
   wire \ram[207][8] ;
   wire \ram[207][7] ;
   wire \ram[207][6] ;
   wire \ram[207][5] ;
   wire \ram[207][4] ;
   wire \ram[207][3] ;
   wire \ram[207][2] ;
   wire \ram[207][1] ;
   wire \ram[207][0] ;
   wire \ram[206][15] ;
   wire \ram[206][14] ;
   wire \ram[206][13] ;
   wire \ram[206][12] ;
   wire \ram[206][11] ;
   wire \ram[206][10] ;
   wire \ram[206][9] ;
   wire \ram[206][8] ;
   wire \ram[206][7] ;
   wire \ram[206][6] ;
   wire \ram[206][5] ;
   wire \ram[206][4] ;
   wire \ram[206][3] ;
   wire \ram[206][2] ;
   wire \ram[206][1] ;
   wire \ram[206][0] ;
   wire \ram[205][15] ;
   wire \ram[205][14] ;
   wire \ram[205][13] ;
   wire \ram[205][12] ;
   wire \ram[205][11] ;
   wire \ram[205][10] ;
   wire \ram[205][9] ;
   wire \ram[205][8] ;
   wire \ram[205][7] ;
   wire \ram[205][6] ;
   wire \ram[205][5] ;
   wire \ram[205][4] ;
   wire \ram[205][3] ;
   wire \ram[205][2] ;
   wire \ram[205][1] ;
   wire \ram[205][0] ;
   wire \ram[204][15] ;
   wire \ram[204][14] ;
   wire \ram[204][13] ;
   wire \ram[204][12] ;
   wire \ram[204][11] ;
   wire \ram[204][10] ;
   wire \ram[204][9] ;
   wire \ram[204][8] ;
   wire \ram[204][7] ;
   wire \ram[204][6] ;
   wire \ram[204][5] ;
   wire \ram[204][4] ;
   wire \ram[204][3] ;
   wire \ram[204][2] ;
   wire \ram[204][1] ;
   wire \ram[204][0] ;
   wire \ram[203][15] ;
   wire \ram[203][14] ;
   wire \ram[203][13] ;
   wire \ram[203][12] ;
   wire \ram[203][11] ;
   wire \ram[203][10] ;
   wire \ram[203][9] ;
   wire \ram[203][8] ;
   wire \ram[203][7] ;
   wire \ram[203][6] ;
   wire \ram[203][5] ;
   wire \ram[203][4] ;
   wire \ram[203][3] ;
   wire \ram[203][2] ;
   wire \ram[203][1] ;
   wire \ram[203][0] ;
   wire \ram[202][15] ;
   wire \ram[202][14] ;
   wire \ram[202][13] ;
   wire \ram[202][12] ;
   wire \ram[202][11] ;
   wire \ram[202][10] ;
   wire \ram[202][9] ;
   wire \ram[202][8] ;
   wire \ram[202][7] ;
   wire \ram[202][6] ;
   wire \ram[202][5] ;
   wire \ram[202][4] ;
   wire \ram[202][3] ;
   wire \ram[202][2] ;
   wire \ram[202][1] ;
   wire \ram[202][0] ;
   wire \ram[201][15] ;
   wire \ram[201][14] ;
   wire \ram[201][13] ;
   wire \ram[201][12] ;
   wire \ram[201][11] ;
   wire \ram[201][10] ;
   wire \ram[201][9] ;
   wire \ram[201][8] ;
   wire \ram[201][7] ;
   wire \ram[201][6] ;
   wire \ram[201][5] ;
   wire \ram[201][4] ;
   wire \ram[201][3] ;
   wire \ram[201][2] ;
   wire \ram[201][1] ;
   wire \ram[201][0] ;
   wire \ram[200][15] ;
   wire \ram[200][14] ;
   wire \ram[200][13] ;
   wire \ram[200][12] ;
   wire \ram[200][11] ;
   wire \ram[200][10] ;
   wire \ram[200][9] ;
   wire \ram[200][8] ;
   wire \ram[200][7] ;
   wire \ram[200][6] ;
   wire \ram[200][5] ;
   wire \ram[200][4] ;
   wire \ram[200][3] ;
   wire \ram[200][2] ;
   wire \ram[200][1] ;
   wire \ram[200][0] ;
   wire \ram[199][15] ;
   wire \ram[199][14] ;
   wire \ram[199][13] ;
   wire \ram[199][12] ;
   wire \ram[199][11] ;
   wire \ram[199][10] ;
   wire \ram[199][9] ;
   wire \ram[199][8] ;
   wire \ram[199][7] ;
   wire \ram[199][6] ;
   wire \ram[199][5] ;
   wire \ram[199][4] ;
   wire \ram[199][3] ;
   wire \ram[199][2] ;
   wire \ram[199][1] ;
   wire \ram[199][0] ;
   wire \ram[198][15] ;
   wire \ram[198][14] ;
   wire \ram[198][13] ;
   wire \ram[198][12] ;
   wire \ram[198][11] ;
   wire \ram[198][10] ;
   wire \ram[198][9] ;
   wire \ram[198][8] ;
   wire \ram[198][7] ;
   wire \ram[198][6] ;
   wire \ram[198][5] ;
   wire \ram[198][4] ;
   wire \ram[198][3] ;
   wire \ram[198][2] ;
   wire \ram[198][1] ;
   wire \ram[198][0] ;
   wire \ram[197][15] ;
   wire \ram[197][14] ;
   wire \ram[197][13] ;
   wire \ram[197][12] ;
   wire \ram[197][11] ;
   wire \ram[197][10] ;
   wire \ram[197][9] ;
   wire \ram[197][8] ;
   wire \ram[197][7] ;
   wire \ram[197][6] ;
   wire \ram[197][5] ;
   wire \ram[197][4] ;
   wire \ram[197][3] ;
   wire \ram[197][2] ;
   wire \ram[197][1] ;
   wire \ram[197][0] ;
   wire \ram[196][15] ;
   wire \ram[196][14] ;
   wire \ram[196][13] ;
   wire \ram[196][12] ;
   wire \ram[196][11] ;
   wire \ram[196][10] ;
   wire \ram[196][9] ;
   wire \ram[196][8] ;
   wire \ram[196][7] ;
   wire \ram[196][6] ;
   wire \ram[196][5] ;
   wire \ram[196][4] ;
   wire \ram[196][3] ;
   wire \ram[196][2] ;
   wire \ram[196][1] ;
   wire \ram[196][0] ;
   wire \ram[195][15] ;
   wire \ram[195][14] ;
   wire \ram[195][13] ;
   wire \ram[195][12] ;
   wire \ram[195][11] ;
   wire \ram[195][10] ;
   wire \ram[195][9] ;
   wire \ram[195][8] ;
   wire \ram[195][7] ;
   wire \ram[195][6] ;
   wire \ram[195][5] ;
   wire \ram[195][4] ;
   wire \ram[195][3] ;
   wire \ram[195][2] ;
   wire \ram[195][1] ;
   wire \ram[195][0] ;
   wire \ram[194][15] ;
   wire \ram[194][14] ;
   wire \ram[194][13] ;
   wire \ram[194][12] ;
   wire \ram[194][11] ;
   wire \ram[194][10] ;
   wire \ram[194][9] ;
   wire \ram[194][8] ;
   wire \ram[194][7] ;
   wire \ram[194][6] ;
   wire \ram[194][5] ;
   wire \ram[194][4] ;
   wire \ram[194][3] ;
   wire \ram[194][2] ;
   wire \ram[194][1] ;
   wire \ram[194][0] ;
   wire \ram[193][15] ;
   wire \ram[193][14] ;
   wire \ram[193][13] ;
   wire \ram[193][12] ;
   wire \ram[193][11] ;
   wire \ram[193][10] ;
   wire \ram[193][9] ;
   wire \ram[193][8] ;
   wire \ram[193][7] ;
   wire \ram[193][6] ;
   wire \ram[193][5] ;
   wire \ram[193][4] ;
   wire \ram[193][3] ;
   wire \ram[193][2] ;
   wire \ram[193][1] ;
   wire \ram[193][0] ;
   wire \ram[192][15] ;
   wire \ram[192][14] ;
   wire \ram[192][13] ;
   wire \ram[192][12] ;
   wire \ram[192][11] ;
   wire \ram[192][10] ;
   wire \ram[192][9] ;
   wire \ram[192][8] ;
   wire \ram[192][7] ;
   wire \ram[192][6] ;
   wire \ram[192][5] ;
   wire \ram[192][4] ;
   wire \ram[192][3] ;
   wire \ram[192][2] ;
   wire \ram[192][1] ;
   wire \ram[192][0] ;
   wire \ram[191][15] ;
   wire \ram[191][14] ;
   wire \ram[191][13] ;
   wire \ram[191][12] ;
   wire \ram[191][11] ;
   wire \ram[191][10] ;
   wire \ram[191][9] ;
   wire \ram[191][8] ;
   wire \ram[191][7] ;
   wire \ram[191][6] ;
   wire \ram[191][5] ;
   wire \ram[191][4] ;
   wire \ram[191][3] ;
   wire \ram[191][2] ;
   wire \ram[191][1] ;
   wire \ram[191][0] ;
   wire \ram[190][15] ;
   wire \ram[190][14] ;
   wire \ram[190][13] ;
   wire \ram[190][12] ;
   wire \ram[190][11] ;
   wire \ram[190][10] ;
   wire \ram[190][9] ;
   wire \ram[190][8] ;
   wire \ram[190][7] ;
   wire \ram[190][6] ;
   wire \ram[190][5] ;
   wire \ram[190][4] ;
   wire \ram[190][3] ;
   wire \ram[190][2] ;
   wire \ram[190][1] ;
   wire \ram[190][0] ;
   wire \ram[189][15] ;
   wire \ram[189][14] ;
   wire \ram[189][13] ;
   wire \ram[189][12] ;
   wire \ram[189][11] ;
   wire \ram[189][10] ;
   wire \ram[189][9] ;
   wire \ram[189][8] ;
   wire \ram[189][7] ;
   wire \ram[189][6] ;
   wire \ram[189][5] ;
   wire \ram[189][4] ;
   wire \ram[189][3] ;
   wire \ram[189][2] ;
   wire \ram[189][1] ;
   wire \ram[189][0] ;
   wire \ram[188][15] ;
   wire \ram[188][14] ;
   wire \ram[188][13] ;
   wire \ram[188][12] ;
   wire \ram[188][11] ;
   wire \ram[188][10] ;
   wire \ram[188][9] ;
   wire \ram[188][8] ;
   wire \ram[188][7] ;
   wire \ram[188][6] ;
   wire \ram[188][5] ;
   wire \ram[188][4] ;
   wire \ram[188][3] ;
   wire \ram[188][2] ;
   wire \ram[188][1] ;
   wire \ram[188][0] ;
   wire \ram[187][15] ;
   wire \ram[187][14] ;
   wire \ram[187][13] ;
   wire \ram[187][12] ;
   wire \ram[187][11] ;
   wire \ram[187][10] ;
   wire \ram[187][9] ;
   wire \ram[187][8] ;
   wire \ram[187][7] ;
   wire \ram[187][6] ;
   wire \ram[187][5] ;
   wire \ram[187][4] ;
   wire \ram[187][3] ;
   wire \ram[187][2] ;
   wire \ram[187][1] ;
   wire \ram[187][0] ;
   wire \ram[186][15] ;
   wire \ram[186][14] ;
   wire \ram[186][13] ;
   wire \ram[186][12] ;
   wire \ram[186][11] ;
   wire \ram[186][10] ;
   wire \ram[186][9] ;
   wire \ram[186][8] ;
   wire \ram[186][7] ;
   wire \ram[186][6] ;
   wire \ram[186][5] ;
   wire \ram[186][4] ;
   wire \ram[186][3] ;
   wire \ram[186][2] ;
   wire \ram[186][1] ;
   wire \ram[186][0] ;
   wire \ram[185][15] ;
   wire \ram[185][14] ;
   wire \ram[185][13] ;
   wire \ram[185][12] ;
   wire \ram[185][11] ;
   wire \ram[185][10] ;
   wire \ram[185][9] ;
   wire \ram[185][8] ;
   wire \ram[185][7] ;
   wire \ram[185][6] ;
   wire \ram[185][5] ;
   wire \ram[185][4] ;
   wire \ram[185][3] ;
   wire \ram[185][2] ;
   wire \ram[185][1] ;
   wire \ram[185][0] ;
   wire \ram[184][15] ;
   wire \ram[184][14] ;
   wire \ram[184][13] ;
   wire \ram[184][12] ;
   wire \ram[184][11] ;
   wire \ram[184][10] ;
   wire \ram[184][9] ;
   wire \ram[184][8] ;
   wire \ram[184][7] ;
   wire \ram[184][6] ;
   wire \ram[184][5] ;
   wire \ram[184][4] ;
   wire \ram[184][3] ;
   wire \ram[184][2] ;
   wire \ram[184][1] ;
   wire \ram[184][0] ;
   wire \ram[183][15] ;
   wire \ram[183][14] ;
   wire \ram[183][13] ;
   wire \ram[183][12] ;
   wire \ram[183][11] ;
   wire \ram[183][10] ;
   wire \ram[183][9] ;
   wire \ram[183][8] ;
   wire \ram[183][7] ;
   wire \ram[183][6] ;
   wire \ram[183][5] ;
   wire \ram[183][4] ;
   wire \ram[183][3] ;
   wire \ram[183][2] ;
   wire \ram[183][1] ;
   wire \ram[183][0] ;
   wire \ram[182][15] ;
   wire \ram[182][14] ;
   wire \ram[182][13] ;
   wire \ram[182][12] ;
   wire \ram[182][11] ;
   wire \ram[182][10] ;
   wire \ram[182][9] ;
   wire \ram[182][8] ;
   wire \ram[182][7] ;
   wire \ram[182][6] ;
   wire \ram[182][5] ;
   wire \ram[182][4] ;
   wire \ram[182][3] ;
   wire \ram[182][2] ;
   wire \ram[182][1] ;
   wire \ram[182][0] ;
   wire \ram[181][15] ;
   wire \ram[181][14] ;
   wire \ram[181][13] ;
   wire \ram[181][12] ;
   wire \ram[181][11] ;
   wire \ram[181][10] ;
   wire \ram[181][9] ;
   wire \ram[181][8] ;
   wire \ram[181][7] ;
   wire \ram[181][6] ;
   wire \ram[181][5] ;
   wire \ram[181][4] ;
   wire \ram[181][3] ;
   wire \ram[181][2] ;
   wire \ram[181][1] ;
   wire \ram[181][0] ;
   wire \ram[180][15] ;
   wire \ram[180][14] ;
   wire \ram[180][13] ;
   wire \ram[180][12] ;
   wire \ram[180][11] ;
   wire \ram[180][10] ;
   wire \ram[180][9] ;
   wire \ram[180][8] ;
   wire \ram[180][7] ;
   wire \ram[180][6] ;
   wire \ram[180][5] ;
   wire \ram[180][4] ;
   wire \ram[180][3] ;
   wire \ram[180][2] ;
   wire \ram[180][1] ;
   wire \ram[180][0] ;
   wire \ram[179][15] ;
   wire \ram[179][14] ;
   wire \ram[179][13] ;
   wire \ram[179][12] ;
   wire \ram[179][11] ;
   wire \ram[179][10] ;
   wire \ram[179][9] ;
   wire \ram[179][8] ;
   wire \ram[179][7] ;
   wire \ram[179][6] ;
   wire \ram[179][5] ;
   wire \ram[179][4] ;
   wire \ram[179][3] ;
   wire \ram[179][2] ;
   wire \ram[179][1] ;
   wire \ram[179][0] ;
   wire \ram[178][15] ;
   wire \ram[178][14] ;
   wire \ram[178][13] ;
   wire \ram[178][12] ;
   wire \ram[178][11] ;
   wire \ram[178][10] ;
   wire \ram[178][9] ;
   wire \ram[178][8] ;
   wire \ram[178][7] ;
   wire \ram[178][6] ;
   wire \ram[178][5] ;
   wire \ram[178][4] ;
   wire \ram[178][3] ;
   wire \ram[178][2] ;
   wire \ram[178][1] ;
   wire \ram[178][0] ;
   wire \ram[177][15] ;
   wire \ram[177][14] ;
   wire \ram[177][13] ;
   wire \ram[177][12] ;
   wire \ram[177][11] ;
   wire \ram[177][10] ;
   wire \ram[177][9] ;
   wire \ram[177][8] ;
   wire \ram[177][7] ;
   wire \ram[177][6] ;
   wire \ram[177][5] ;
   wire \ram[177][4] ;
   wire \ram[177][3] ;
   wire \ram[177][2] ;
   wire \ram[177][1] ;
   wire \ram[177][0] ;
   wire \ram[176][15] ;
   wire \ram[176][14] ;
   wire \ram[176][13] ;
   wire \ram[176][12] ;
   wire \ram[176][11] ;
   wire \ram[176][10] ;
   wire \ram[176][9] ;
   wire \ram[176][8] ;
   wire \ram[176][7] ;
   wire \ram[176][6] ;
   wire \ram[176][5] ;
   wire \ram[176][4] ;
   wire \ram[176][3] ;
   wire \ram[176][2] ;
   wire \ram[176][1] ;
   wire \ram[176][0] ;
   wire \ram[175][15] ;
   wire \ram[175][14] ;
   wire \ram[175][13] ;
   wire \ram[175][12] ;
   wire \ram[175][11] ;
   wire \ram[175][10] ;
   wire \ram[175][9] ;
   wire \ram[175][8] ;
   wire \ram[175][7] ;
   wire \ram[175][6] ;
   wire \ram[175][5] ;
   wire \ram[175][4] ;
   wire \ram[175][3] ;
   wire \ram[175][2] ;
   wire \ram[175][1] ;
   wire \ram[175][0] ;
   wire \ram[174][15] ;
   wire \ram[174][14] ;
   wire \ram[174][13] ;
   wire \ram[174][12] ;
   wire \ram[174][11] ;
   wire \ram[174][10] ;
   wire \ram[174][9] ;
   wire \ram[174][8] ;
   wire \ram[174][7] ;
   wire \ram[174][6] ;
   wire \ram[174][5] ;
   wire \ram[174][4] ;
   wire \ram[174][3] ;
   wire \ram[174][2] ;
   wire \ram[174][1] ;
   wire \ram[174][0] ;
   wire \ram[173][15] ;
   wire \ram[173][14] ;
   wire \ram[173][13] ;
   wire \ram[173][12] ;
   wire \ram[173][11] ;
   wire \ram[173][10] ;
   wire \ram[173][9] ;
   wire \ram[173][8] ;
   wire \ram[173][7] ;
   wire \ram[173][6] ;
   wire \ram[173][5] ;
   wire \ram[173][4] ;
   wire \ram[173][3] ;
   wire \ram[173][2] ;
   wire \ram[173][1] ;
   wire \ram[173][0] ;
   wire \ram[172][15] ;
   wire \ram[172][14] ;
   wire \ram[172][13] ;
   wire \ram[172][12] ;
   wire \ram[172][11] ;
   wire \ram[172][10] ;
   wire \ram[172][9] ;
   wire \ram[172][8] ;
   wire \ram[172][7] ;
   wire \ram[172][6] ;
   wire \ram[172][5] ;
   wire \ram[172][4] ;
   wire \ram[172][3] ;
   wire \ram[172][2] ;
   wire \ram[172][1] ;
   wire \ram[172][0] ;
   wire \ram[171][15] ;
   wire \ram[171][14] ;
   wire \ram[171][13] ;
   wire \ram[171][12] ;
   wire \ram[171][11] ;
   wire \ram[171][10] ;
   wire \ram[171][9] ;
   wire \ram[171][8] ;
   wire \ram[171][7] ;
   wire \ram[171][6] ;
   wire \ram[171][5] ;
   wire \ram[171][4] ;
   wire \ram[171][3] ;
   wire \ram[171][2] ;
   wire \ram[171][1] ;
   wire \ram[171][0] ;
   wire \ram[170][15] ;
   wire \ram[170][14] ;
   wire \ram[170][13] ;
   wire \ram[170][12] ;
   wire \ram[170][11] ;
   wire \ram[170][10] ;
   wire \ram[170][9] ;
   wire \ram[170][8] ;
   wire \ram[170][7] ;
   wire \ram[170][6] ;
   wire \ram[170][5] ;
   wire \ram[170][4] ;
   wire \ram[170][3] ;
   wire \ram[170][2] ;
   wire \ram[170][1] ;
   wire \ram[170][0] ;
   wire \ram[169][15] ;
   wire \ram[169][14] ;
   wire \ram[169][13] ;
   wire \ram[169][12] ;
   wire \ram[169][11] ;
   wire \ram[169][10] ;
   wire \ram[169][9] ;
   wire \ram[169][8] ;
   wire \ram[169][7] ;
   wire \ram[169][6] ;
   wire \ram[169][5] ;
   wire \ram[169][4] ;
   wire \ram[169][3] ;
   wire \ram[169][2] ;
   wire \ram[169][1] ;
   wire \ram[169][0] ;
   wire \ram[168][15] ;
   wire \ram[168][14] ;
   wire \ram[168][13] ;
   wire \ram[168][12] ;
   wire \ram[168][11] ;
   wire \ram[168][10] ;
   wire \ram[168][9] ;
   wire \ram[168][8] ;
   wire \ram[168][7] ;
   wire \ram[168][6] ;
   wire \ram[168][5] ;
   wire \ram[168][4] ;
   wire \ram[168][3] ;
   wire \ram[168][2] ;
   wire \ram[168][1] ;
   wire \ram[168][0] ;
   wire \ram[167][15] ;
   wire \ram[167][14] ;
   wire \ram[167][13] ;
   wire \ram[167][12] ;
   wire \ram[167][11] ;
   wire \ram[167][10] ;
   wire \ram[167][9] ;
   wire \ram[167][8] ;
   wire \ram[167][7] ;
   wire \ram[167][6] ;
   wire \ram[167][5] ;
   wire \ram[167][4] ;
   wire \ram[167][3] ;
   wire \ram[167][2] ;
   wire \ram[167][1] ;
   wire \ram[167][0] ;
   wire \ram[166][15] ;
   wire \ram[166][14] ;
   wire \ram[166][13] ;
   wire \ram[166][12] ;
   wire \ram[166][11] ;
   wire \ram[166][10] ;
   wire \ram[166][9] ;
   wire \ram[166][8] ;
   wire \ram[166][7] ;
   wire \ram[166][6] ;
   wire \ram[166][5] ;
   wire \ram[166][4] ;
   wire \ram[166][3] ;
   wire \ram[166][2] ;
   wire \ram[166][1] ;
   wire \ram[166][0] ;
   wire \ram[165][15] ;
   wire \ram[165][14] ;
   wire \ram[165][13] ;
   wire \ram[165][12] ;
   wire \ram[165][11] ;
   wire \ram[165][10] ;
   wire \ram[165][9] ;
   wire \ram[165][8] ;
   wire \ram[165][7] ;
   wire \ram[165][6] ;
   wire \ram[165][5] ;
   wire \ram[165][4] ;
   wire \ram[165][3] ;
   wire \ram[165][2] ;
   wire \ram[165][1] ;
   wire \ram[165][0] ;
   wire \ram[164][15] ;
   wire \ram[164][14] ;
   wire \ram[164][13] ;
   wire \ram[164][12] ;
   wire \ram[164][11] ;
   wire \ram[164][10] ;
   wire \ram[164][9] ;
   wire \ram[164][8] ;
   wire \ram[164][7] ;
   wire \ram[164][6] ;
   wire \ram[164][5] ;
   wire \ram[164][4] ;
   wire \ram[164][3] ;
   wire \ram[164][2] ;
   wire \ram[164][1] ;
   wire \ram[164][0] ;
   wire \ram[163][15] ;
   wire \ram[163][14] ;
   wire \ram[163][13] ;
   wire \ram[163][12] ;
   wire \ram[163][11] ;
   wire \ram[163][10] ;
   wire \ram[163][9] ;
   wire \ram[163][8] ;
   wire \ram[163][7] ;
   wire \ram[163][6] ;
   wire \ram[163][5] ;
   wire \ram[163][4] ;
   wire \ram[163][3] ;
   wire \ram[163][2] ;
   wire \ram[163][1] ;
   wire \ram[163][0] ;
   wire \ram[162][15] ;
   wire \ram[162][14] ;
   wire \ram[162][13] ;
   wire \ram[162][12] ;
   wire \ram[162][11] ;
   wire \ram[162][10] ;
   wire \ram[162][9] ;
   wire \ram[162][8] ;
   wire \ram[162][7] ;
   wire \ram[162][6] ;
   wire \ram[162][5] ;
   wire \ram[162][4] ;
   wire \ram[162][3] ;
   wire \ram[162][2] ;
   wire \ram[162][1] ;
   wire \ram[162][0] ;
   wire \ram[161][15] ;
   wire \ram[161][14] ;
   wire \ram[161][13] ;
   wire \ram[161][12] ;
   wire \ram[161][11] ;
   wire \ram[161][10] ;
   wire \ram[161][9] ;
   wire \ram[161][8] ;
   wire \ram[161][7] ;
   wire \ram[161][6] ;
   wire \ram[161][5] ;
   wire \ram[161][4] ;
   wire \ram[161][3] ;
   wire \ram[161][2] ;
   wire \ram[161][1] ;
   wire \ram[161][0] ;
   wire \ram[160][15] ;
   wire \ram[160][14] ;
   wire \ram[160][13] ;
   wire \ram[160][12] ;
   wire \ram[160][11] ;
   wire \ram[160][10] ;
   wire \ram[160][9] ;
   wire \ram[160][8] ;
   wire \ram[160][7] ;
   wire \ram[160][6] ;
   wire \ram[160][5] ;
   wire \ram[160][4] ;
   wire \ram[160][3] ;
   wire \ram[160][2] ;
   wire \ram[160][1] ;
   wire \ram[160][0] ;
   wire \ram[159][15] ;
   wire \ram[159][14] ;
   wire \ram[159][13] ;
   wire \ram[159][12] ;
   wire \ram[159][11] ;
   wire \ram[159][10] ;
   wire \ram[159][9] ;
   wire \ram[159][8] ;
   wire \ram[159][7] ;
   wire \ram[159][6] ;
   wire \ram[159][5] ;
   wire \ram[159][4] ;
   wire \ram[159][3] ;
   wire \ram[159][2] ;
   wire \ram[159][1] ;
   wire \ram[159][0] ;
   wire \ram[158][15] ;
   wire \ram[158][14] ;
   wire \ram[158][13] ;
   wire \ram[158][12] ;
   wire \ram[158][11] ;
   wire \ram[158][10] ;
   wire \ram[158][9] ;
   wire \ram[158][8] ;
   wire \ram[158][7] ;
   wire \ram[158][6] ;
   wire \ram[158][5] ;
   wire \ram[158][4] ;
   wire \ram[158][3] ;
   wire \ram[158][2] ;
   wire \ram[158][1] ;
   wire \ram[158][0] ;
   wire \ram[157][15] ;
   wire \ram[157][14] ;
   wire \ram[157][13] ;
   wire \ram[157][12] ;
   wire \ram[157][11] ;
   wire \ram[157][10] ;
   wire \ram[157][9] ;
   wire \ram[157][8] ;
   wire \ram[157][7] ;
   wire \ram[157][6] ;
   wire \ram[157][5] ;
   wire \ram[157][4] ;
   wire \ram[157][3] ;
   wire \ram[157][2] ;
   wire \ram[157][1] ;
   wire \ram[157][0] ;
   wire \ram[156][15] ;
   wire \ram[156][14] ;
   wire \ram[156][13] ;
   wire \ram[156][12] ;
   wire \ram[156][11] ;
   wire \ram[156][10] ;
   wire \ram[156][9] ;
   wire \ram[156][8] ;
   wire \ram[156][7] ;
   wire \ram[156][6] ;
   wire \ram[156][5] ;
   wire \ram[156][4] ;
   wire \ram[156][3] ;
   wire \ram[156][2] ;
   wire \ram[156][1] ;
   wire \ram[156][0] ;
   wire \ram[155][15] ;
   wire \ram[155][14] ;
   wire \ram[155][13] ;
   wire \ram[155][12] ;
   wire \ram[155][11] ;
   wire \ram[155][10] ;
   wire \ram[155][9] ;
   wire \ram[155][8] ;
   wire \ram[155][7] ;
   wire \ram[155][6] ;
   wire \ram[155][5] ;
   wire \ram[155][4] ;
   wire \ram[155][3] ;
   wire \ram[155][2] ;
   wire \ram[155][1] ;
   wire \ram[155][0] ;
   wire \ram[154][15] ;
   wire \ram[154][14] ;
   wire \ram[154][13] ;
   wire \ram[154][12] ;
   wire \ram[154][11] ;
   wire \ram[154][10] ;
   wire \ram[154][9] ;
   wire \ram[154][8] ;
   wire \ram[154][7] ;
   wire \ram[154][6] ;
   wire \ram[154][5] ;
   wire \ram[154][4] ;
   wire \ram[154][3] ;
   wire \ram[154][2] ;
   wire \ram[154][1] ;
   wire \ram[154][0] ;
   wire \ram[153][15] ;
   wire \ram[153][14] ;
   wire \ram[153][13] ;
   wire \ram[153][12] ;
   wire \ram[153][11] ;
   wire \ram[153][10] ;
   wire \ram[153][9] ;
   wire \ram[153][8] ;
   wire \ram[153][7] ;
   wire \ram[153][6] ;
   wire \ram[153][5] ;
   wire \ram[153][4] ;
   wire \ram[153][3] ;
   wire \ram[153][2] ;
   wire \ram[153][1] ;
   wire \ram[153][0] ;
   wire \ram[152][15] ;
   wire \ram[152][14] ;
   wire \ram[152][13] ;
   wire \ram[152][12] ;
   wire \ram[152][11] ;
   wire \ram[152][10] ;
   wire \ram[152][9] ;
   wire \ram[152][8] ;
   wire \ram[152][7] ;
   wire \ram[152][6] ;
   wire \ram[152][5] ;
   wire \ram[152][4] ;
   wire \ram[152][3] ;
   wire \ram[152][2] ;
   wire \ram[152][1] ;
   wire \ram[152][0] ;
   wire \ram[151][15] ;
   wire \ram[151][14] ;
   wire \ram[151][13] ;
   wire \ram[151][12] ;
   wire \ram[151][11] ;
   wire \ram[151][10] ;
   wire \ram[151][9] ;
   wire \ram[151][8] ;
   wire \ram[151][7] ;
   wire \ram[151][6] ;
   wire \ram[151][5] ;
   wire \ram[151][4] ;
   wire \ram[151][3] ;
   wire \ram[151][2] ;
   wire \ram[151][1] ;
   wire \ram[151][0] ;
   wire \ram[150][15] ;
   wire \ram[150][14] ;
   wire \ram[150][13] ;
   wire \ram[150][12] ;
   wire \ram[150][11] ;
   wire \ram[150][10] ;
   wire \ram[150][9] ;
   wire \ram[150][8] ;
   wire \ram[150][7] ;
   wire \ram[150][6] ;
   wire \ram[150][5] ;
   wire \ram[150][4] ;
   wire \ram[150][3] ;
   wire \ram[150][2] ;
   wire \ram[150][1] ;
   wire \ram[150][0] ;
   wire \ram[149][15] ;
   wire \ram[149][14] ;
   wire \ram[149][13] ;
   wire \ram[149][12] ;
   wire \ram[149][11] ;
   wire \ram[149][10] ;
   wire \ram[149][9] ;
   wire \ram[149][8] ;
   wire \ram[149][7] ;
   wire \ram[149][6] ;
   wire \ram[149][5] ;
   wire \ram[149][4] ;
   wire \ram[149][3] ;
   wire \ram[149][2] ;
   wire \ram[149][1] ;
   wire \ram[149][0] ;
   wire \ram[148][15] ;
   wire \ram[148][14] ;
   wire \ram[148][13] ;
   wire \ram[148][12] ;
   wire \ram[148][11] ;
   wire \ram[148][10] ;
   wire \ram[148][9] ;
   wire \ram[148][8] ;
   wire \ram[148][7] ;
   wire \ram[148][6] ;
   wire \ram[148][5] ;
   wire \ram[148][4] ;
   wire \ram[148][3] ;
   wire \ram[148][2] ;
   wire \ram[148][1] ;
   wire \ram[148][0] ;
   wire \ram[147][15] ;
   wire \ram[147][14] ;
   wire \ram[147][13] ;
   wire \ram[147][12] ;
   wire \ram[147][11] ;
   wire \ram[147][10] ;
   wire \ram[147][9] ;
   wire \ram[147][8] ;
   wire \ram[147][7] ;
   wire \ram[147][6] ;
   wire \ram[147][5] ;
   wire \ram[147][4] ;
   wire \ram[147][3] ;
   wire \ram[147][2] ;
   wire \ram[147][1] ;
   wire \ram[147][0] ;
   wire \ram[146][15] ;
   wire \ram[146][14] ;
   wire \ram[146][13] ;
   wire \ram[146][12] ;
   wire \ram[146][11] ;
   wire \ram[146][10] ;
   wire \ram[146][9] ;
   wire \ram[146][8] ;
   wire \ram[146][7] ;
   wire \ram[146][6] ;
   wire \ram[146][5] ;
   wire \ram[146][4] ;
   wire \ram[146][3] ;
   wire \ram[146][2] ;
   wire \ram[146][1] ;
   wire \ram[146][0] ;
   wire \ram[145][15] ;
   wire \ram[145][14] ;
   wire \ram[145][13] ;
   wire \ram[145][12] ;
   wire \ram[145][11] ;
   wire \ram[145][10] ;
   wire \ram[145][9] ;
   wire \ram[145][8] ;
   wire \ram[145][7] ;
   wire \ram[145][6] ;
   wire \ram[145][5] ;
   wire \ram[145][4] ;
   wire \ram[145][3] ;
   wire \ram[145][2] ;
   wire \ram[145][1] ;
   wire \ram[145][0] ;
   wire \ram[144][15] ;
   wire \ram[144][14] ;
   wire \ram[144][13] ;
   wire \ram[144][12] ;
   wire \ram[144][11] ;
   wire \ram[144][10] ;
   wire \ram[144][9] ;
   wire \ram[144][8] ;
   wire \ram[144][7] ;
   wire \ram[144][6] ;
   wire \ram[144][5] ;
   wire \ram[144][4] ;
   wire \ram[144][3] ;
   wire \ram[144][2] ;
   wire \ram[144][1] ;
   wire \ram[144][0] ;
   wire \ram[143][15] ;
   wire \ram[143][14] ;
   wire \ram[143][13] ;
   wire \ram[143][12] ;
   wire \ram[143][11] ;
   wire \ram[143][10] ;
   wire \ram[143][9] ;
   wire \ram[143][8] ;
   wire \ram[143][7] ;
   wire \ram[143][6] ;
   wire \ram[143][5] ;
   wire \ram[143][4] ;
   wire \ram[143][3] ;
   wire \ram[143][2] ;
   wire \ram[143][1] ;
   wire \ram[143][0] ;
   wire \ram[142][15] ;
   wire \ram[142][14] ;
   wire \ram[142][13] ;
   wire \ram[142][12] ;
   wire \ram[142][11] ;
   wire \ram[142][10] ;
   wire \ram[142][9] ;
   wire \ram[142][8] ;
   wire \ram[142][7] ;
   wire \ram[142][6] ;
   wire \ram[142][5] ;
   wire \ram[142][4] ;
   wire \ram[142][3] ;
   wire \ram[142][2] ;
   wire \ram[142][1] ;
   wire \ram[142][0] ;
   wire \ram[141][15] ;
   wire \ram[141][14] ;
   wire \ram[141][13] ;
   wire \ram[141][12] ;
   wire \ram[141][11] ;
   wire \ram[141][10] ;
   wire \ram[141][9] ;
   wire \ram[141][8] ;
   wire \ram[141][7] ;
   wire \ram[141][6] ;
   wire \ram[141][5] ;
   wire \ram[141][4] ;
   wire \ram[141][3] ;
   wire \ram[141][2] ;
   wire \ram[141][1] ;
   wire \ram[141][0] ;
   wire \ram[140][15] ;
   wire \ram[140][14] ;
   wire \ram[140][13] ;
   wire \ram[140][12] ;
   wire \ram[140][11] ;
   wire \ram[140][10] ;
   wire \ram[140][9] ;
   wire \ram[140][8] ;
   wire \ram[140][7] ;
   wire \ram[140][6] ;
   wire \ram[140][5] ;
   wire \ram[140][4] ;
   wire \ram[140][3] ;
   wire \ram[140][2] ;
   wire \ram[140][1] ;
   wire \ram[140][0] ;
   wire \ram[139][15] ;
   wire \ram[139][14] ;
   wire \ram[139][13] ;
   wire \ram[139][12] ;
   wire \ram[139][11] ;
   wire \ram[139][10] ;
   wire \ram[139][9] ;
   wire \ram[139][8] ;
   wire \ram[139][7] ;
   wire \ram[139][6] ;
   wire \ram[139][5] ;
   wire \ram[139][4] ;
   wire \ram[139][3] ;
   wire \ram[139][2] ;
   wire \ram[139][1] ;
   wire \ram[139][0] ;
   wire \ram[138][15] ;
   wire \ram[138][14] ;
   wire \ram[138][13] ;
   wire \ram[138][12] ;
   wire \ram[138][11] ;
   wire \ram[138][10] ;
   wire \ram[138][9] ;
   wire \ram[138][8] ;
   wire \ram[138][7] ;
   wire \ram[138][6] ;
   wire \ram[138][5] ;
   wire \ram[138][4] ;
   wire \ram[138][3] ;
   wire \ram[138][2] ;
   wire \ram[138][1] ;
   wire \ram[138][0] ;
   wire \ram[137][15] ;
   wire \ram[137][14] ;
   wire \ram[137][13] ;
   wire \ram[137][12] ;
   wire \ram[137][11] ;
   wire \ram[137][10] ;
   wire \ram[137][9] ;
   wire \ram[137][8] ;
   wire \ram[137][7] ;
   wire \ram[137][6] ;
   wire \ram[137][5] ;
   wire \ram[137][4] ;
   wire \ram[137][3] ;
   wire \ram[137][2] ;
   wire \ram[137][1] ;
   wire \ram[137][0] ;
   wire \ram[136][15] ;
   wire \ram[136][14] ;
   wire \ram[136][13] ;
   wire \ram[136][12] ;
   wire \ram[136][11] ;
   wire \ram[136][10] ;
   wire \ram[136][9] ;
   wire \ram[136][8] ;
   wire \ram[136][7] ;
   wire \ram[136][6] ;
   wire \ram[136][5] ;
   wire \ram[136][4] ;
   wire \ram[136][3] ;
   wire \ram[136][2] ;
   wire \ram[136][1] ;
   wire \ram[136][0] ;
   wire \ram[135][15] ;
   wire \ram[135][14] ;
   wire \ram[135][13] ;
   wire \ram[135][12] ;
   wire \ram[135][11] ;
   wire \ram[135][10] ;
   wire \ram[135][9] ;
   wire \ram[135][8] ;
   wire \ram[135][7] ;
   wire \ram[135][6] ;
   wire \ram[135][5] ;
   wire \ram[135][4] ;
   wire \ram[135][3] ;
   wire \ram[135][2] ;
   wire \ram[135][1] ;
   wire \ram[135][0] ;
   wire \ram[134][15] ;
   wire \ram[134][14] ;
   wire \ram[134][13] ;
   wire \ram[134][12] ;
   wire \ram[134][11] ;
   wire \ram[134][10] ;
   wire \ram[134][9] ;
   wire \ram[134][8] ;
   wire \ram[134][7] ;
   wire \ram[134][6] ;
   wire \ram[134][5] ;
   wire \ram[134][4] ;
   wire \ram[134][3] ;
   wire \ram[134][2] ;
   wire \ram[134][1] ;
   wire \ram[134][0] ;
   wire \ram[133][15] ;
   wire \ram[133][14] ;
   wire \ram[133][13] ;
   wire \ram[133][12] ;
   wire \ram[133][11] ;
   wire \ram[133][10] ;
   wire \ram[133][9] ;
   wire \ram[133][8] ;
   wire \ram[133][7] ;
   wire \ram[133][6] ;
   wire \ram[133][5] ;
   wire \ram[133][4] ;
   wire \ram[133][3] ;
   wire \ram[133][2] ;
   wire \ram[133][1] ;
   wire \ram[133][0] ;
   wire \ram[132][15] ;
   wire \ram[132][14] ;
   wire \ram[132][13] ;
   wire \ram[132][12] ;
   wire \ram[132][11] ;
   wire \ram[132][10] ;
   wire \ram[132][9] ;
   wire \ram[132][8] ;
   wire \ram[132][7] ;
   wire \ram[132][6] ;
   wire \ram[132][5] ;
   wire \ram[132][4] ;
   wire \ram[132][3] ;
   wire \ram[132][2] ;
   wire \ram[132][1] ;
   wire \ram[132][0] ;
   wire \ram[131][15] ;
   wire \ram[131][14] ;
   wire \ram[131][13] ;
   wire \ram[131][12] ;
   wire \ram[131][11] ;
   wire \ram[131][10] ;
   wire \ram[131][9] ;
   wire \ram[131][8] ;
   wire \ram[131][7] ;
   wire \ram[131][6] ;
   wire \ram[131][5] ;
   wire \ram[131][4] ;
   wire \ram[131][3] ;
   wire \ram[131][2] ;
   wire \ram[131][1] ;
   wire \ram[131][0] ;
   wire \ram[130][15] ;
   wire \ram[130][14] ;
   wire \ram[130][13] ;
   wire \ram[130][12] ;
   wire \ram[130][11] ;
   wire \ram[130][10] ;
   wire \ram[130][9] ;
   wire \ram[130][8] ;
   wire \ram[130][7] ;
   wire \ram[130][6] ;
   wire \ram[130][5] ;
   wire \ram[130][4] ;
   wire \ram[130][3] ;
   wire \ram[130][2] ;
   wire \ram[130][1] ;
   wire \ram[130][0] ;
   wire \ram[129][15] ;
   wire \ram[129][14] ;
   wire \ram[129][13] ;
   wire \ram[129][12] ;
   wire \ram[129][11] ;
   wire \ram[129][10] ;
   wire \ram[129][9] ;
   wire \ram[129][8] ;
   wire \ram[129][7] ;
   wire \ram[129][6] ;
   wire \ram[129][5] ;
   wire \ram[129][4] ;
   wire \ram[129][3] ;
   wire \ram[129][2] ;
   wire \ram[129][1] ;
   wire \ram[129][0] ;
   wire \ram[128][15] ;
   wire \ram[128][14] ;
   wire \ram[128][13] ;
   wire \ram[128][12] ;
   wire \ram[128][11] ;
   wire \ram[128][10] ;
   wire \ram[128][9] ;
   wire \ram[128][8] ;
   wire \ram[128][7] ;
   wire \ram[128][6] ;
   wire \ram[128][5] ;
   wire \ram[128][4] ;
   wire \ram[128][3] ;
   wire \ram[128][2] ;
   wire \ram[128][1] ;
   wire \ram[128][0] ;
   wire \ram[127][15] ;
   wire \ram[127][14] ;
   wire \ram[127][13] ;
   wire \ram[127][12] ;
   wire \ram[127][11] ;
   wire \ram[127][10] ;
   wire \ram[127][9] ;
   wire \ram[127][8] ;
   wire \ram[127][7] ;
   wire \ram[127][6] ;
   wire \ram[127][5] ;
   wire \ram[127][4] ;
   wire \ram[127][3] ;
   wire \ram[127][2] ;
   wire \ram[127][1] ;
   wire \ram[127][0] ;
   wire \ram[126][15] ;
   wire \ram[126][14] ;
   wire \ram[126][13] ;
   wire \ram[126][12] ;
   wire \ram[126][11] ;
   wire \ram[126][10] ;
   wire \ram[126][9] ;
   wire \ram[126][8] ;
   wire \ram[126][7] ;
   wire \ram[126][6] ;
   wire \ram[126][5] ;
   wire \ram[126][4] ;
   wire \ram[126][3] ;
   wire \ram[126][2] ;
   wire \ram[126][1] ;
   wire \ram[126][0] ;
   wire \ram[125][15] ;
   wire \ram[125][14] ;
   wire \ram[125][13] ;
   wire \ram[125][12] ;
   wire \ram[125][11] ;
   wire \ram[125][10] ;
   wire \ram[125][9] ;
   wire \ram[125][8] ;
   wire \ram[125][7] ;
   wire \ram[125][6] ;
   wire \ram[125][5] ;
   wire \ram[125][4] ;
   wire \ram[125][3] ;
   wire \ram[125][2] ;
   wire \ram[125][1] ;
   wire \ram[125][0] ;
   wire \ram[124][15] ;
   wire \ram[124][14] ;
   wire \ram[124][13] ;
   wire \ram[124][12] ;
   wire \ram[124][11] ;
   wire \ram[124][10] ;
   wire \ram[124][9] ;
   wire \ram[124][8] ;
   wire \ram[124][7] ;
   wire \ram[124][6] ;
   wire \ram[124][5] ;
   wire \ram[124][4] ;
   wire \ram[124][3] ;
   wire \ram[124][2] ;
   wire \ram[124][1] ;
   wire \ram[124][0] ;
   wire \ram[123][15] ;
   wire \ram[123][14] ;
   wire \ram[123][13] ;
   wire \ram[123][12] ;
   wire \ram[123][11] ;
   wire \ram[123][10] ;
   wire \ram[123][9] ;
   wire \ram[123][8] ;
   wire \ram[123][7] ;
   wire \ram[123][6] ;
   wire \ram[123][5] ;
   wire \ram[123][4] ;
   wire \ram[123][3] ;
   wire \ram[123][2] ;
   wire \ram[123][1] ;
   wire \ram[123][0] ;
   wire \ram[122][15] ;
   wire \ram[122][14] ;
   wire \ram[122][13] ;
   wire \ram[122][12] ;
   wire \ram[122][11] ;
   wire \ram[122][10] ;
   wire \ram[122][9] ;
   wire \ram[122][8] ;
   wire \ram[122][7] ;
   wire \ram[122][6] ;
   wire \ram[122][5] ;
   wire \ram[122][4] ;
   wire \ram[122][3] ;
   wire \ram[122][2] ;
   wire \ram[122][1] ;
   wire \ram[122][0] ;
   wire \ram[121][15] ;
   wire \ram[121][14] ;
   wire \ram[121][13] ;
   wire \ram[121][12] ;
   wire \ram[121][11] ;
   wire \ram[121][10] ;
   wire \ram[121][9] ;
   wire \ram[121][8] ;
   wire \ram[121][7] ;
   wire \ram[121][6] ;
   wire \ram[121][5] ;
   wire \ram[121][4] ;
   wire \ram[121][3] ;
   wire \ram[121][2] ;
   wire \ram[121][1] ;
   wire \ram[121][0] ;
   wire \ram[120][15] ;
   wire \ram[120][14] ;
   wire \ram[120][13] ;
   wire \ram[120][12] ;
   wire \ram[120][11] ;
   wire \ram[120][10] ;
   wire \ram[120][9] ;
   wire \ram[120][8] ;
   wire \ram[120][7] ;
   wire \ram[120][6] ;
   wire \ram[120][5] ;
   wire \ram[120][4] ;
   wire \ram[120][3] ;
   wire \ram[120][2] ;
   wire \ram[120][1] ;
   wire \ram[120][0] ;
   wire \ram[119][15] ;
   wire \ram[119][14] ;
   wire \ram[119][13] ;
   wire \ram[119][12] ;
   wire \ram[119][11] ;
   wire \ram[119][10] ;
   wire \ram[119][9] ;
   wire \ram[119][8] ;
   wire \ram[119][7] ;
   wire \ram[119][6] ;
   wire \ram[119][5] ;
   wire \ram[119][4] ;
   wire \ram[119][3] ;
   wire \ram[119][2] ;
   wire \ram[119][1] ;
   wire \ram[119][0] ;
   wire \ram[118][15] ;
   wire \ram[118][14] ;
   wire \ram[118][13] ;
   wire \ram[118][12] ;
   wire \ram[118][11] ;
   wire \ram[118][10] ;
   wire \ram[118][9] ;
   wire \ram[118][8] ;
   wire \ram[118][7] ;
   wire \ram[118][6] ;
   wire \ram[118][5] ;
   wire \ram[118][4] ;
   wire \ram[118][3] ;
   wire \ram[118][2] ;
   wire \ram[118][1] ;
   wire \ram[118][0] ;
   wire \ram[117][15] ;
   wire \ram[117][14] ;
   wire \ram[117][13] ;
   wire \ram[117][12] ;
   wire \ram[117][11] ;
   wire \ram[117][10] ;
   wire \ram[117][9] ;
   wire \ram[117][8] ;
   wire \ram[117][7] ;
   wire \ram[117][6] ;
   wire \ram[117][5] ;
   wire \ram[117][4] ;
   wire \ram[117][3] ;
   wire \ram[117][2] ;
   wire \ram[117][1] ;
   wire \ram[117][0] ;
   wire \ram[116][15] ;
   wire \ram[116][14] ;
   wire \ram[116][13] ;
   wire \ram[116][12] ;
   wire \ram[116][11] ;
   wire \ram[116][10] ;
   wire \ram[116][9] ;
   wire \ram[116][8] ;
   wire \ram[116][7] ;
   wire \ram[116][6] ;
   wire \ram[116][5] ;
   wire \ram[116][4] ;
   wire \ram[116][3] ;
   wire \ram[116][2] ;
   wire \ram[116][1] ;
   wire \ram[116][0] ;
   wire \ram[115][15] ;
   wire \ram[115][14] ;
   wire \ram[115][13] ;
   wire \ram[115][12] ;
   wire \ram[115][11] ;
   wire \ram[115][10] ;
   wire \ram[115][9] ;
   wire \ram[115][8] ;
   wire \ram[115][7] ;
   wire \ram[115][6] ;
   wire \ram[115][5] ;
   wire \ram[115][4] ;
   wire \ram[115][3] ;
   wire \ram[115][2] ;
   wire \ram[115][1] ;
   wire \ram[115][0] ;
   wire \ram[114][15] ;
   wire \ram[114][14] ;
   wire \ram[114][13] ;
   wire \ram[114][12] ;
   wire \ram[114][11] ;
   wire \ram[114][10] ;
   wire \ram[114][9] ;
   wire \ram[114][8] ;
   wire \ram[114][7] ;
   wire \ram[114][6] ;
   wire \ram[114][5] ;
   wire \ram[114][4] ;
   wire \ram[114][3] ;
   wire \ram[114][2] ;
   wire \ram[114][1] ;
   wire \ram[114][0] ;
   wire \ram[113][15] ;
   wire \ram[113][14] ;
   wire \ram[113][13] ;
   wire \ram[113][12] ;
   wire \ram[113][11] ;
   wire \ram[113][10] ;
   wire \ram[113][9] ;
   wire \ram[113][8] ;
   wire \ram[113][7] ;
   wire \ram[113][6] ;
   wire \ram[113][5] ;
   wire \ram[113][4] ;
   wire \ram[113][3] ;
   wire \ram[113][2] ;
   wire \ram[113][1] ;
   wire \ram[113][0] ;
   wire \ram[112][15] ;
   wire \ram[112][14] ;
   wire \ram[112][13] ;
   wire \ram[112][12] ;
   wire \ram[112][11] ;
   wire \ram[112][10] ;
   wire \ram[112][9] ;
   wire \ram[112][8] ;
   wire \ram[112][7] ;
   wire \ram[112][6] ;
   wire \ram[112][5] ;
   wire \ram[112][4] ;
   wire \ram[112][3] ;
   wire \ram[112][2] ;
   wire \ram[112][1] ;
   wire \ram[112][0] ;
   wire \ram[111][15] ;
   wire \ram[111][14] ;
   wire \ram[111][13] ;
   wire \ram[111][12] ;
   wire \ram[111][11] ;
   wire \ram[111][10] ;
   wire \ram[111][9] ;
   wire \ram[111][8] ;
   wire \ram[111][7] ;
   wire \ram[111][6] ;
   wire \ram[111][5] ;
   wire \ram[111][4] ;
   wire \ram[111][3] ;
   wire \ram[111][2] ;
   wire \ram[111][1] ;
   wire \ram[111][0] ;
   wire \ram[110][15] ;
   wire \ram[110][14] ;
   wire \ram[110][13] ;
   wire \ram[110][12] ;
   wire \ram[110][11] ;
   wire \ram[110][10] ;
   wire \ram[110][9] ;
   wire \ram[110][8] ;
   wire \ram[110][7] ;
   wire \ram[110][6] ;
   wire \ram[110][5] ;
   wire \ram[110][4] ;
   wire \ram[110][3] ;
   wire \ram[110][2] ;
   wire \ram[110][1] ;
   wire \ram[110][0] ;
   wire \ram[109][15] ;
   wire \ram[109][14] ;
   wire \ram[109][13] ;
   wire \ram[109][12] ;
   wire \ram[109][11] ;
   wire \ram[109][10] ;
   wire \ram[109][9] ;
   wire \ram[109][8] ;
   wire \ram[109][7] ;
   wire \ram[109][6] ;
   wire \ram[109][5] ;
   wire \ram[109][4] ;
   wire \ram[109][3] ;
   wire \ram[109][2] ;
   wire \ram[109][1] ;
   wire \ram[109][0] ;
   wire \ram[108][15] ;
   wire \ram[108][14] ;
   wire \ram[108][13] ;
   wire \ram[108][12] ;
   wire \ram[108][11] ;
   wire \ram[108][10] ;
   wire \ram[108][9] ;
   wire \ram[108][8] ;
   wire \ram[108][7] ;
   wire \ram[108][6] ;
   wire \ram[108][5] ;
   wire \ram[108][4] ;
   wire \ram[108][3] ;
   wire \ram[108][2] ;
   wire \ram[108][1] ;
   wire \ram[108][0] ;
   wire \ram[107][15] ;
   wire \ram[107][14] ;
   wire \ram[107][13] ;
   wire \ram[107][12] ;
   wire \ram[107][11] ;
   wire \ram[107][10] ;
   wire \ram[107][9] ;
   wire \ram[107][8] ;
   wire \ram[107][7] ;
   wire \ram[107][6] ;
   wire \ram[107][5] ;
   wire \ram[107][4] ;
   wire \ram[107][3] ;
   wire \ram[107][2] ;
   wire \ram[107][1] ;
   wire \ram[107][0] ;
   wire \ram[106][15] ;
   wire \ram[106][14] ;
   wire \ram[106][13] ;
   wire \ram[106][12] ;
   wire \ram[106][11] ;
   wire \ram[106][10] ;
   wire \ram[106][9] ;
   wire \ram[106][8] ;
   wire \ram[106][7] ;
   wire \ram[106][6] ;
   wire \ram[106][5] ;
   wire \ram[106][4] ;
   wire \ram[106][3] ;
   wire \ram[106][2] ;
   wire \ram[106][1] ;
   wire \ram[106][0] ;
   wire \ram[105][15] ;
   wire \ram[105][14] ;
   wire \ram[105][13] ;
   wire \ram[105][12] ;
   wire \ram[105][11] ;
   wire \ram[105][10] ;
   wire \ram[105][9] ;
   wire \ram[105][8] ;
   wire \ram[105][7] ;
   wire \ram[105][6] ;
   wire \ram[105][5] ;
   wire \ram[105][4] ;
   wire \ram[105][3] ;
   wire \ram[105][2] ;
   wire \ram[105][1] ;
   wire \ram[105][0] ;
   wire \ram[104][15] ;
   wire \ram[104][14] ;
   wire \ram[104][13] ;
   wire \ram[104][12] ;
   wire \ram[104][11] ;
   wire \ram[104][10] ;
   wire \ram[104][9] ;
   wire \ram[104][8] ;
   wire \ram[104][7] ;
   wire \ram[104][6] ;
   wire \ram[104][5] ;
   wire \ram[104][4] ;
   wire \ram[104][3] ;
   wire \ram[104][2] ;
   wire \ram[104][1] ;
   wire \ram[104][0] ;
   wire \ram[103][15] ;
   wire \ram[103][14] ;
   wire \ram[103][13] ;
   wire \ram[103][12] ;
   wire \ram[103][11] ;
   wire \ram[103][10] ;
   wire \ram[103][9] ;
   wire \ram[103][8] ;
   wire \ram[103][7] ;
   wire \ram[103][6] ;
   wire \ram[103][5] ;
   wire \ram[103][4] ;
   wire \ram[103][3] ;
   wire \ram[103][2] ;
   wire \ram[103][1] ;
   wire \ram[103][0] ;
   wire \ram[102][15] ;
   wire \ram[102][14] ;
   wire \ram[102][13] ;
   wire \ram[102][12] ;
   wire \ram[102][11] ;
   wire \ram[102][10] ;
   wire \ram[102][9] ;
   wire \ram[102][8] ;
   wire \ram[102][7] ;
   wire \ram[102][6] ;
   wire \ram[102][5] ;
   wire \ram[102][4] ;
   wire \ram[102][3] ;
   wire \ram[102][2] ;
   wire \ram[102][1] ;
   wire \ram[102][0] ;
   wire \ram[101][15] ;
   wire \ram[101][14] ;
   wire \ram[101][13] ;
   wire \ram[101][12] ;
   wire \ram[101][11] ;
   wire \ram[101][10] ;
   wire \ram[101][9] ;
   wire \ram[101][8] ;
   wire \ram[101][7] ;
   wire \ram[101][6] ;
   wire \ram[101][5] ;
   wire \ram[101][4] ;
   wire \ram[101][3] ;
   wire \ram[101][2] ;
   wire \ram[101][1] ;
   wire \ram[101][0] ;
   wire \ram[100][15] ;
   wire \ram[100][14] ;
   wire \ram[100][13] ;
   wire \ram[100][12] ;
   wire \ram[100][11] ;
   wire \ram[100][10] ;
   wire \ram[100][9] ;
   wire \ram[100][8] ;
   wire \ram[100][7] ;
   wire \ram[100][6] ;
   wire \ram[100][5] ;
   wire \ram[100][4] ;
   wire \ram[100][3] ;
   wire \ram[100][2] ;
   wire \ram[100][1] ;
   wire \ram[100][0] ;
   wire \ram[99][15] ;
   wire \ram[99][14] ;
   wire \ram[99][13] ;
   wire \ram[99][12] ;
   wire \ram[99][11] ;
   wire \ram[99][10] ;
   wire \ram[99][9] ;
   wire \ram[99][8] ;
   wire \ram[99][7] ;
   wire \ram[99][6] ;
   wire \ram[99][5] ;
   wire \ram[99][4] ;
   wire \ram[99][3] ;
   wire \ram[99][2] ;
   wire \ram[99][1] ;
   wire \ram[99][0] ;
   wire \ram[98][15] ;
   wire \ram[98][14] ;
   wire \ram[98][13] ;
   wire \ram[98][12] ;
   wire \ram[98][11] ;
   wire \ram[98][10] ;
   wire \ram[98][9] ;
   wire \ram[98][8] ;
   wire \ram[98][7] ;
   wire \ram[98][6] ;
   wire \ram[98][5] ;
   wire \ram[98][4] ;
   wire \ram[98][3] ;
   wire \ram[98][2] ;
   wire \ram[98][1] ;
   wire \ram[98][0] ;
   wire \ram[97][15] ;
   wire \ram[97][14] ;
   wire \ram[97][13] ;
   wire \ram[97][12] ;
   wire \ram[97][11] ;
   wire \ram[97][10] ;
   wire \ram[97][9] ;
   wire \ram[97][8] ;
   wire \ram[97][7] ;
   wire \ram[97][6] ;
   wire \ram[97][5] ;
   wire \ram[97][4] ;
   wire \ram[97][3] ;
   wire \ram[97][2] ;
   wire \ram[97][1] ;
   wire \ram[97][0] ;
   wire \ram[96][15] ;
   wire \ram[96][14] ;
   wire \ram[96][13] ;
   wire \ram[96][12] ;
   wire \ram[96][11] ;
   wire \ram[96][10] ;
   wire \ram[96][9] ;
   wire \ram[96][8] ;
   wire \ram[96][7] ;
   wire \ram[96][6] ;
   wire \ram[96][5] ;
   wire \ram[96][4] ;
   wire \ram[96][3] ;
   wire \ram[96][2] ;
   wire \ram[96][1] ;
   wire \ram[96][0] ;
   wire \ram[95][15] ;
   wire \ram[95][14] ;
   wire \ram[95][13] ;
   wire \ram[95][12] ;
   wire \ram[95][11] ;
   wire \ram[95][10] ;
   wire \ram[95][9] ;
   wire \ram[95][8] ;
   wire \ram[95][7] ;
   wire \ram[95][6] ;
   wire \ram[95][5] ;
   wire \ram[95][4] ;
   wire \ram[95][3] ;
   wire \ram[95][2] ;
   wire \ram[95][1] ;
   wire \ram[95][0] ;
   wire \ram[94][15] ;
   wire \ram[94][14] ;
   wire \ram[94][13] ;
   wire \ram[94][12] ;
   wire \ram[94][11] ;
   wire \ram[94][10] ;
   wire \ram[94][9] ;
   wire \ram[94][8] ;
   wire \ram[94][7] ;
   wire \ram[94][6] ;
   wire \ram[94][5] ;
   wire \ram[94][4] ;
   wire \ram[94][3] ;
   wire \ram[94][2] ;
   wire \ram[94][1] ;
   wire \ram[94][0] ;
   wire \ram[93][15] ;
   wire \ram[93][14] ;
   wire \ram[93][13] ;
   wire \ram[93][12] ;
   wire \ram[93][11] ;
   wire \ram[93][10] ;
   wire \ram[93][9] ;
   wire \ram[93][8] ;
   wire \ram[93][7] ;
   wire \ram[93][6] ;
   wire \ram[93][5] ;
   wire \ram[93][4] ;
   wire \ram[93][3] ;
   wire \ram[93][2] ;
   wire \ram[93][1] ;
   wire \ram[93][0] ;
   wire \ram[92][15] ;
   wire \ram[92][14] ;
   wire \ram[92][13] ;
   wire \ram[92][12] ;
   wire \ram[92][11] ;
   wire \ram[92][10] ;
   wire \ram[92][9] ;
   wire \ram[92][8] ;
   wire \ram[92][7] ;
   wire \ram[92][6] ;
   wire \ram[92][5] ;
   wire \ram[92][4] ;
   wire \ram[92][3] ;
   wire \ram[92][2] ;
   wire \ram[92][1] ;
   wire \ram[92][0] ;
   wire \ram[91][15] ;
   wire \ram[91][14] ;
   wire \ram[91][13] ;
   wire \ram[91][12] ;
   wire \ram[91][11] ;
   wire \ram[91][10] ;
   wire \ram[91][9] ;
   wire \ram[91][8] ;
   wire \ram[91][7] ;
   wire \ram[91][6] ;
   wire \ram[91][5] ;
   wire \ram[91][4] ;
   wire \ram[91][3] ;
   wire \ram[91][2] ;
   wire \ram[91][1] ;
   wire \ram[91][0] ;
   wire \ram[90][15] ;
   wire \ram[90][14] ;
   wire \ram[90][13] ;
   wire \ram[90][12] ;
   wire \ram[90][11] ;
   wire \ram[90][10] ;
   wire \ram[90][9] ;
   wire \ram[90][8] ;
   wire \ram[90][7] ;
   wire \ram[90][6] ;
   wire \ram[90][5] ;
   wire \ram[90][4] ;
   wire \ram[90][3] ;
   wire \ram[90][2] ;
   wire \ram[90][1] ;
   wire \ram[90][0] ;
   wire \ram[89][15] ;
   wire \ram[89][14] ;
   wire \ram[89][13] ;
   wire \ram[89][12] ;
   wire \ram[89][11] ;
   wire \ram[89][10] ;
   wire \ram[89][9] ;
   wire \ram[89][8] ;
   wire \ram[89][7] ;
   wire \ram[89][6] ;
   wire \ram[89][5] ;
   wire \ram[89][4] ;
   wire \ram[89][3] ;
   wire \ram[89][2] ;
   wire \ram[89][1] ;
   wire \ram[89][0] ;
   wire \ram[88][15] ;
   wire \ram[88][14] ;
   wire \ram[88][13] ;
   wire \ram[88][12] ;
   wire \ram[88][11] ;
   wire \ram[88][10] ;
   wire \ram[88][9] ;
   wire \ram[88][8] ;
   wire \ram[88][7] ;
   wire \ram[88][6] ;
   wire \ram[88][5] ;
   wire \ram[88][4] ;
   wire \ram[88][3] ;
   wire \ram[88][2] ;
   wire \ram[88][1] ;
   wire \ram[88][0] ;
   wire \ram[87][15] ;
   wire \ram[87][14] ;
   wire \ram[87][13] ;
   wire \ram[87][12] ;
   wire \ram[87][11] ;
   wire \ram[87][10] ;
   wire \ram[87][9] ;
   wire \ram[87][8] ;
   wire \ram[87][7] ;
   wire \ram[87][6] ;
   wire \ram[87][5] ;
   wire \ram[87][4] ;
   wire \ram[87][3] ;
   wire \ram[87][2] ;
   wire \ram[87][1] ;
   wire \ram[87][0] ;
   wire \ram[86][15] ;
   wire \ram[86][14] ;
   wire \ram[86][13] ;
   wire \ram[86][12] ;
   wire \ram[86][11] ;
   wire \ram[86][10] ;
   wire \ram[86][9] ;
   wire \ram[86][8] ;
   wire \ram[86][7] ;
   wire \ram[86][6] ;
   wire \ram[86][5] ;
   wire \ram[86][4] ;
   wire \ram[86][3] ;
   wire \ram[86][2] ;
   wire \ram[86][1] ;
   wire \ram[86][0] ;
   wire \ram[85][15] ;
   wire \ram[85][14] ;
   wire \ram[85][13] ;
   wire \ram[85][12] ;
   wire \ram[85][11] ;
   wire \ram[85][10] ;
   wire \ram[85][9] ;
   wire \ram[85][8] ;
   wire \ram[85][7] ;
   wire \ram[85][6] ;
   wire \ram[85][5] ;
   wire \ram[85][4] ;
   wire \ram[85][3] ;
   wire \ram[85][2] ;
   wire \ram[85][1] ;
   wire \ram[85][0] ;
   wire \ram[84][15] ;
   wire \ram[84][14] ;
   wire \ram[84][13] ;
   wire \ram[84][12] ;
   wire \ram[84][11] ;
   wire \ram[84][10] ;
   wire \ram[84][9] ;
   wire \ram[84][8] ;
   wire \ram[84][7] ;
   wire \ram[84][6] ;
   wire \ram[84][5] ;
   wire \ram[84][4] ;
   wire \ram[84][3] ;
   wire \ram[84][2] ;
   wire \ram[84][1] ;
   wire \ram[84][0] ;
   wire \ram[83][15] ;
   wire \ram[83][14] ;
   wire \ram[83][13] ;
   wire \ram[83][12] ;
   wire \ram[83][11] ;
   wire \ram[83][10] ;
   wire \ram[83][9] ;
   wire \ram[83][8] ;
   wire \ram[83][7] ;
   wire \ram[83][6] ;
   wire \ram[83][5] ;
   wire \ram[83][4] ;
   wire \ram[83][3] ;
   wire \ram[83][2] ;
   wire \ram[83][1] ;
   wire \ram[83][0] ;
   wire \ram[82][15] ;
   wire \ram[82][14] ;
   wire \ram[82][13] ;
   wire \ram[82][12] ;
   wire \ram[82][11] ;
   wire \ram[82][10] ;
   wire \ram[82][9] ;
   wire \ram[82][8] ;
   wire \ram[82][7] ;
   wire \ram[82][6] ;
   wire \ram[82][5] ;
   wire \ram[82][4] ;
   wire \ram[82][3] ;
   wire \ram[82][2] ;
   wire \ram[82][1] ;
   wire \ram[82][0] ;
   wire \ram[81][15] ;
   wire \ram[81][14] ;
   wire \ram[81][13] ;
   wire \ram[81][12] ;
   wire \ram[81][11] ;
   wire \ram[81][10] ;
   wire \ram[81][9] ;
   wire \ram[81][8] ;
   wire \ram[81][7] ;
   wire \ram[81][6] ;
   wire \ram[81][5] ;
   wire \ram[81][4] ;
   wire \ram[81][3] ;
   wire \ram[81][2] ;
   wire \ram[81][1] ;
   wire \ram[81][0] ;
   wire \ram[80][15] ;
   wire \ram[80][14] ;
   wire \ram[80][13] ;
   wire \ram[80][12] ;
   wire \ram[80][11] ;
   wire \ram[80][10] ;
   wire \ram[80][9] ;
   wire \ram[80][8] ;
   wire \ram[80][7] ;
   wire \ram[80][6] ;
   wire \ram[80][5] ;
   wire \ram[80][4] ;
   wire \ram[80][3] ;
   wire \ram[80][2] ;
   wire \ram[80][1] ;
   wire \ram[80][0] ;
   wire \ram[79][15] ;
   wire \ram[79][14] ;
   wire \ram[79][13] ;
   wire \ram[79][12] ;
   wire \ram[79][11] ;
   wire \ram[79][10] ;
   wire \ram[79][9] ;
   wire \ram[79][8] ;
   wire \ram[79][7] ;
   wire \ram[79][6] ;
   wire \ram[79][5] ;
   wire \ram[79][4] ;
   wire \ram[79][3] ;
   wire \ram[79][2] ;
   wire \ram[79][1] ;
   wire \ram[79][0] ;
   wire \ram[78][15] ;
   wire \ram[78][14] ;
   wire \ram[78][13] ;
   wire \ram[78][12] ;
   wire \ram[78][11] ;
   wire \ram[78][10] ;
   wire \ram[78][9] ;
   wire \ram[78][8] ;
   wire \ram[78][7] ;
   wire \ram[78][6] ;
   wire \ram[78][5] ;
   wire \ram[78][4] ;
   wire \ram[78][3] ;
   wire \ram[78][2] ;
   wire \ram[78][1] ;
   wire \ram[78][0] ;
   wire \ram[77][15] ;
   wire \ram[77][14] ;
   wire \ram[77][13] ;
   wire \ram[77][12] ;
   wire \ram[77][11] ;
   wire \ram[77][10] ;
   wire \ram[77][9] ;
   wire \ram[77][8] ;
   wire \ram[77][7] ;
   wire \ram[77][6] ;
   wire \ram[77][5] ;
   wire \ram[77][4] ;
   wire \ram[77][3] ;
   wire \ram[77][2] ;
   wire \ram[77][1] ;
   wire \ram[77][0] ;
   wire \ram[76][15] ;
   wire \ram[76][14] ;
   wire \ram[76][13] ;
   wire \ram[76][12] ;
   wire \ram[76][11] ;
   wire \ram[76][10] ;
   wire \ram[76][9] ;
   wire \ram[76][8] ;
   wire \ram[76][7] ;
   wire \ram[76][6] ;
   wire \ram[76][5] ;
   wire \ram[76][4] ;
   wire \ram[76][3] ;
   wire \ram[76][2] ;
   wire \ram[76][1] ;
   wire \ram[76][0] ;
   wire \ram[75][15] ;
   wire \ram[75][14] ;
   wire \ram[75][13] ;
   wire \ram[75][12] ;
   wire \ram[75][11] ;
   wire \ram[75][10] ;
   wire \ram[75][9] ;
   wire \ram[75][8] ;
   wire \ram[75][7] ;
   wire \ram[75][6] ;
   wire \ram[75][5] ;
   wire \ram[75][4] ;
   wire \ram[75][3] ;
   wire \ram[75][2] ;
   wire \ram[75][1] ;
   wire \ram[75][0] ;
   wire \ram[74][15] ;
   wire \ram[74][14] ;
   wire \ram[74][13] ;
   wire \ram[74][12] ;
   wire \ram[74][11] ;
   wire \ram[74][10] ;
   wire \ram[74][9] ;
   wire \ram[74][8] ;
   wire \ram[74][7] ;
   wire \ram[74][6] ;
   wire \ram[74][5] ;
   wire \ram[74][4] ;
   wire \ram[74][3] ;
   wire \ram[74][2] ;
   wire \ram[74][1] ;
   wire \ram[74][0] ;
   wire \ram[73][15] ;
   wire \ram[73][14] ;
   wire \ram[73][13] ;
   wire \ram[73][12] ;
   wire \ram[73][11] ;
   wire \ram[73][10] ;
   wire \ram[73][9] ;
   wire \ram[73][8] ;
   wire \ram[73][7] ;
   wire \ram[73][6] ;
   wire \ram[73][5] ;
   wire \ram[73][4] ;
   wire \ram[73][3] ;
   wire \ram[73][2] ;
   wire \ram[73][1] ;
   wire \ram[73][0] ;
   wire \ram[72][15] ;
   wire \ram[72][14] ;
   wire \ram[72][13] ;
   wire \ram[72][12] ;
   wire \ram[72][11] ;
   wire \ram[72][10] ;
   wire \ram[72][9] ;
   wire \ram[72][8] ;
   wire \ram[72][7] ;
   wire \ram[72][6] ;
   wire \ram[72][5] ;
   wire \ram[72][4] ;
   wire \ram[72][3] ;
   wire \ram[72][2] ;
   wire \ram[72][1] ;
   wire \ram[72][0] ;
   wire \ram[71][15] ;
   wire \ram[71][14] ;
   wire \ram[71][13] ;
   wire \ram[71][12] ;
   wire \ram[71][11] ;
   wire \ram[71][10] ;
   wire \ram[71][9] ;
   wire \ram[71][8] ;
   wire \ram[71][7] ;
   wire \ram[71][6] ;
   wire \ram[71][5] ;
   wire \ram[71][4] ;
   wire \ram[71][3] ;
   wire \ram[71][2] ;
   wire \ram[71][1] ;
   wire \ram[71][0] ;
   wire \ram[70][15] ;
   wire \ram[70][14] ;
   wire \ram[70][13] ;
   wire \ram[70][12] ;
   wire \ram[70][11] ;
   wire \ram[70][10] ;
   wire \ram[70][9] ;
   wire \ram[70][8] ;
   wire \ram[70][7] ;
   wire \ram[70][6] ;
   wire \ram[70][5] ;
   wire \ram[70][4] ;
   wire \ram[70][3] ;
   wire \ram[70][2] ;
   wire \ram[70][1] ;
   wire \ram[70][0] ;
   wire \ram[69][15] ;
   wire \ram[69][14] ;
   wire \ram[69][13] ;
   wire \ram[69][12] ;
   wire \ram[69][11] ;
   wire \ram[69][10] ;
   wire \ram[69][9] ;
   wire \ram[69][8] ;
   wire \ram[69][7] ;
   wire \ram[69][6] ;
   wire \ram[69][5] ;
   wire \ram[69][4] ;
   wire \ram[69][3] ;
   wire \ram[69][2] ;
   wire \ram[69][1] ;
   wire \ram[69][0] ;
   wire \ram[68][15] ;
   wire \ram[68][14] ;
   wire \ram[68][13] ;
   wire \ram[68][12] ;
   wire \ram[68][11] ;
   wire \ram[68][10] ;
   wire \ram[68][9] ;
   wire \ram[68][8] ;
   wire \ram[68][7] ;
   wire \ram[68][6] ;
   wire \ram[68][5] ;
   wire \ram[68][4] ;
   wire \ram[68][3] ;
   wire \ram[68][2] ;
   wire \ram[68][1] ;
   wire \ram[68][0] ;
   wire \ram[67][15] ;
   wire \ram[67][14] ;
   wire \ram[67][13] ;
   wire \ram[67][12] ;
   wire \ram[67][11] ;
   wire \ram[67][10] ;
   wire \ram[67][9] ;
   wire \ram[67][8] ;
   wire \ram[67][7] ;
   wire \ram[67][6] ;
   wire \ram[67][5] ;
   wire \ram[67][4] ;
   wire \ram[67][3] ;
   wire \ram[67][2] ;
   wire \ram[67][1] ;
   wire \ram[67][0] ;
   wire \ram[66][15] ;
   wire \ram[66][14] ;
   wire \ram[66][13] ;
   wire \ram[66][12] ;
   wire \ram[66][11] ;
   wire \ram[66][10] ;
   wire \ram[66][9] ;
   wire \ram[66][8] ;
   wire \ram[66][7] ;
   wire \ram[66][6] ;
   wire \ram[66][5] ;
   wire \ram[66][4] ;
   wire \ram[66][3] ;
   wire \ram[66][2] ;
   wire \ram[66][1] ;
   wire \ram[66][0] ;
   wire \ram[65][15] ;
   wire \ram[65][14] ;
   wire \ram[65][13] ;
   wire \ram[65][12] ;
   wire \ram[65][11] ;
   wire \ram[65][10] ;
   wire \ram[65][9] ;
   wire \ram[65][8] ;
   wire \ram[65][7] ;
   wire \ram[65][6] ;
   wire \ram[65][5] ;
   wire \ram[65][4] ;
   wire \ram[65][3] ;
   wire \ram[65][2] ;
   wire \ram[65][1] ;
   wire \ram[65][0] ;
   wire \ram[64][15] ;
   wire \ram[64][14] ;
   wire \ram[64][13] ;
   wire \ram[64][12] ;
   wire \ram[64][11] ;
   wire \ram[64][10] ;
   wire \ram[64][9] ;
   wire \ram[64][8] ;
   wire \ram[64][7] ;
   wire \ram[64][6] ;
   wire \ram[64][5] ;
   wire \ram[64][4] ;
   wire \ram[64][3] ;
   wire \ram[64][2] ;
   wire \ram[64][1] ;
   wire \ram[64][0] ;
   wire \ram[63][15] ;
   wire \ram[63][14] ;
   wire \ram[63][13] ;
   wire \ram[63][12] ;
   wire \ram[63][11] ;
   wire \ram[63][10] ;
   wire \ram[63][9] ;
   wire \ram[63][8] ;
   wire \ram[63][7] ;
   wire \ram[63][6] ;
   wire \ram[63][5] ;
   wire \ram[63][4] ;
   wire \ram[63][3] ;
   wire \ram[63][2] ;
   wire \ram[63][1] ;
   wire \ram[63][0] ;
   wire \ram[62][15] ;
   wire \ram[62][14] ;
   wire \ram[62][13] ;
   wire \ram[62][12] ;
   wire \ram[62][11] ;
   wire \ram[62][10] ;
   wire \ram[62][9] ;
   wire \ram[62][8] ;
   wire \ram[62][7] ;
   wire \ram[62][6] ;
   wire \ram[62][5] ;
   wire \ram[62][4] ;
   wire \ram[62][3] ;
   wire \ram[62][2] ;
   wire \ram[62][1] ;
   wire \ram[62][0] ;
   wire \ram[61][15] ;
   wire \ram[61][14] ;
   wire \ram[61][13] ;
   wire \ram[61][12] ;
   wire \ram[61][11] ;
   wire \ram[61][10] ;
   wire \ram[61][9] ;
   wire \ram[61][8] ;
   wire \ram[61][7] ;
   wire \ram[61][6] ;
   wire \ram[61][5] ;
   wire \ram[61][4] ;
   wire \ram[61][3] ;
   wire \ram[61][2] ;
   wire \ram[61][1] ;
   wire \ram[61][0] ;
   wire \ram[60][15] ;
   wire \ram[60][14] ;
   wire \ram[60][13] ;
   wire \ram[60][12] ;
   wire \ram[60][11] ;
   wire \ram[60][10] ;
   wire \ram[60][9] ;
   wire \ram[60][8] ;
   wire \ram[60][7] ;
   wire \ram[60][6] ;
   wire \ram[60][5] ;
   wire \ram[60][4] ;
   wire \ram[60][3] ;
   wire \ram[60][2] ;
   wire \ram[60][1] ;
   wire \ram[60][0] ;
   wire \ram[59][15] ;
   wire \ram[59][14] ;
   wire \ram[59][13] ;
   wire \ram[59][12] ;
   wire \ram[59][11] ;
   wire \ram[59][10] ;
   wire \ram[59][9] ;
   wire \ram[59][8] ;
   wire \ram[59][7] ;
   wire \ram[59][6] ;
   wire \ram[59][5] ;
   wire \ram[59][4] ;
   wire \ram[59][3] ;
   wire \ram[59][2] ;
   wire \ram[59][1] ;
   wire \ram[59][0] ;
   wire \ram[58][15] ;
   wire \ram[58][14] ;
   wire \ram[58][13] ;
   wire \ram[58][12] ;
   wire \ram[58][11] ;
   wire \ram[58][10] ;
   wire \ram[58][9] ;
   wire \ram[58][8] ;
   wire \ram[58][7] ;
   wire \ram[58][6] ;
   wire \ram[58][5] ;
   wire \ram[58][4] ;
   wire \ram[58][3] ;
   wire \ram[58][2] ;
   wire \ram[58][1] ;
   wire \ram[58][0] ;
   wire \ram[57][15] ;
   wire \ram[57][14] ;
   wire \ram[57][13] ;
   wire \ram[57][12] ;
   wire \ram[57][11] ;
   wire \ram[57][10] ;
   wire \ram[57][9] ;
   wire \ram[57][8] ;
   wire \ram[57][7] ;
   wire \ram[57][6] ;
   wire \ram[57][5] ;
   wire \ram[57][4] ;
   wire \ram[57][3] ;
   wire \ram[57][2] ;
   wire \ram[57][1] ;
   wire \ram[57][0] ;
   wire \ram[56][15] ;
   wire \ram[56][14] ;
   wire \ram[56][13] ;
   wire \ram[56][12] ;
   wire \ram[56][11] ;
   wire \ram[56][10] ;
   wire \ram[56][9] ;
   wire \ram[56][8] ;
   wire \ram[56][7] ;
   wire \ram[56][6] ;
   wire \ram[56][5] ;
   wire \ram[56][4] ;
   wire \ram[56][3] ;
   wire \ram[56][2] ;
   wire \ram[56][1] ;
   wire \ram[56][0] ;
   wire \ram[55][15] ;
   wire \ram[55][14] ;
   wire \ram[55][13] ;
   wire \ram[55][12] ;
   wire \ram[55][11] ;
   wire \ram[55][10] ;
   wire \ram[55][9] ;
   wire \ram[55][8] ;
   wire \ram[55][7] ;
   wire \ram[55][6] ;
   wire \ram[55][5] ;
   wire \ram[55][4] ;
   wire \ram[55][3] ;
   wire \ram[55][2] ;
   wire \ram[55][1] ;
   wire \ram[55][0] ;
   wire \ram[54][15] ;
   wire \ram[54][14] ;
   wire \ram[54][13] ;
   wire \ram[54][12] ;
   wire \ram[54][11] ;
   wire \ram[54][10] ;
   wire \ram[54][9] ;
   wire \ram[54][8] ;
   wire \ram[54][7] ;
   wire \ram[54][6] ;
   wire \ram[54][5] ;
   wire \ram[54][4] ;
   wire \ram[54][3] ;
   wire \ram[54][2] ;
   wire \ram[54][1] ;
   wire \ram[54][0] ;
   wire \ram[53][15] ;
   wire \ram[53][14] ;
   wire \ram[53][13] ;
   wire \ram[53][12] ;
   wire \ram[53][11] ;
   wire \ram[53][10] ;
   wire \ram[53][9] ;
   wire \ram[53][8] ;
   wire \ram[53][7] ;
   wire \ram[53][6] ;
   wire \ram[53][5] ;
   wire \ram[53][4] ;
   wire \ram[53][3] ;
   wire \ram[53][2] ;
   wire \ram[53][1] ;
   wire \ram[53][0] ;
   wire \ram[52][15] ;
   wire \ram[52][14] ;
   wire \ram[52][13] ;
   wire \ram[52][12] ;
   wire \ram[52][11] ;
   wire \ram[52][10] ;
   wire \ram[52][9] ;
   wire \ram[52][8] ;
   wire \ram[52][7] ;
   wire \ram[52][6] ;
   wire \ram[52][5] ;
   wire \ram[52][4] ;
   wire \ram[52][3] ;
   wire \ram[52][2] ;
   wire \ram[52][1] ;
   wire \ram[52][0] ;
   wire \ram[51][15] ;
   wire \ram[51][14] ;
   wire \ram[51][13] ;
   wire \ram[51][12] ;
   wire \ram[51][11] ;
   wire \ram[51][10] ;
   wire \ram[51][9] ;
   wire \ram[51][8] ;
   wire \ram[51][7] ;
   wire \ram[51][6] ;
   wire \ram[51][5] ;
   wire \ram[51][4] ;
   wire \ram[51][3] ;
   wire \ram[51][2] ;
   wire \ram[51][1] ;
   wire \ram[51][0] ;
   wire \ram[50][15] ;
   wire \ram[50][14] ;
   wire \ram[50][13] ;
   wire \ram[50][12] ;
   wire \ram[50][11] ;
   wire \ram[50][10] ;
   wire \ram[50][9] ;
   wire \ram[50][8] ;
   wire \ram[50][7] ;
   wire \ram[50][6] ;
   wire \ram[50][5] ;
   wire \ram[50][4] ;
   wire \ram[50][3] ;
   wire \ram[50][2] ;
   wire \ram[50][1] ;
   wire \ram[50][0] ;
   wire \ram[49][15] ;
   wire \ram[49][14] ;
   wire \ram[49][13] ;
   wire \ram[49][12] ;
   wire \ram[49][11] ;
   wire \ram[49][10] ;
   wire \ram[49][9] ;
   wire \ram[49][8] ;
   wire \ram[49][7] ;
   wire \ram[49][6] ;
   wire \ram[49][5] ;
   wire \ram[49][4] ;
   wire \ram[49][3] ;
   wire \ram[49][2] ;
   wire \ram[49][1] ;
   wire \ram[49][0] ;
   wire \ram[48][15] ;
   wire \ram[48][14] ;
   wire \ram[48][13] ;
   wire \ram[48][12] ;
   wire \ram[48][11] ;
   wire \ram[48][10] ;
   wire \ram[48][9] ;
   wire \ram[48][8] ;
   wire \ram[48][7] ;
   wire \ram[48][6] ;
   wire \ram[48][5] ;
   wire \ram[48][4] ;
   wire \ram[48][3] ;
   wire \ram[48][2] ;
   wire \ram[48][1] ;
   wire \ram[48][0] ;
   wire \ram[47][15] ;
   wire \ram[47][14] ;
   wire \ram[47][13] ;
   wire \ram[47][12] ;
   wire \ram[47][11] ;
   wire \ram[47][10] ;
   wire \ram[47][9] ;
   wire \ram[47][8] ;
   wire \ram[47][7] ;
   wire \ram[47][6] ;
   wire \ram[47][5] ;
   wire \ram[47][4] ;
   wire \ram[47][3] ;
   wire \ram[47][2] ;
   wire \ram[47][1] ;
   wire \ram[47][0] ;
   wire \ram[46][15] ;
   wire \ram[46][14] ;
   wire \ram[46][13] ;
   wire \ram[46][12] ;
   wire \ram[46][11] ;
   wire \ram[46][10] ;
   wire \ram[46][9] ;
   wire \ram[46][8] ;
   wire \ram[46][7] ;
   wire \ram[46][6] ;
   wire \ram[46][5] ;
   wire \ram[46][4] ;
   wire \ram[46][3] ;
   wire \ram[46][2] ;
   wire \ram[46][1] ;
   wire \ram[46][0] ;
   wire \ram[45][15] ;
   wire \ram[45][14] ;
   wire \ram[45][13] ;
   wire \ram[45][12] ;
   wire \ram[45][11] ;
   wire \ram[45][10] ;
   wire \ram[45][9] ;
   wire \ram[45][8] ;
   wire \ram[45][7] ;
   wire \ram[45][6] ;
   wire \ram[45][5] ;
   wire \ram[45][4] ;
   wire \ram[45][3] ;
   wire \ram[45][2] ;
   wire \ram[45][1] ;
   wire \ram[45][0] ;
   wire \ram[44][15] ;
   wire \ram[44][14] ;
   wire \ram[44][13] ;
   wire \ram[44][12] ;
   wire \ram[44][11] ;
   wire \ram[44][10] ;
   wire \ram[44][9] ;
   wire \ram[44][8] ;
   wire \ram[44][7] ;
   wire \ram[44][6] ;
   wire \ram[44][5] ;
   wire \ram[44][4] ;
   wire \ram[44][3] ;
   wire \ram[44][2] ;
   wire \ram[44][1] ;
   wire \ram[44][0] ;
   wire \ram[43][15] ;
   wire \ram[43][14] ;
   wire \ram[43][13] ;
   wire \ram[43][12] ;
   wire \ram[43][11] ;
   wire \ram[43][10] ;
   wire \ram[43][9] ;
   wire \ram[43][8] ;
   wire \ram[43][7] ;
   wire \ram[43][6] ;
   wire \ram[43][5] ;
   wire \ram[43][4] ;
   wire \ram[43][3] ;
   wire \ram[43][2] ;
   wire \ram[43][1] ;
   wire \ram[43][0] ;
   wire \ram[42][15] ;
   wire \ram[42][14] ;
   wire \ram[42][13] ;
   wire \ram[42][12] ;
   wire \ram[42][11] ;
   wire \ram[42][10] ;
   wire \ram[42][9] ;
   wire \ram[42][8] ;
   wire \ram[42][7] ;
   wire \ram[42][6] ;
   wire \ram[42][5] ;
   wire \ram[42][4] ;
   wire \ram[42][3] ;
   wire \ram[42][2] ;
   wire \ram[42][1] ;
   wire \ram[42][0] ;
   wire \ram[41][15] ;
   wire \ram[41][14] ;
   wire \ram[41][13] ;
   wire \ram[41][12] ;
   wire \ram[41][11] ;
   wire \ram[41][10] ;
   wire \ram[41][9] ;
   wire \ram[41][8] ;
   wire \ram[41][7] ;
   wire \ram[41][6] ;
   wire \ram[41][5] ;
   wire \ram[41][4] ;
   wire \ram[41][3] ;
   wire \ram[41][2] ;
   wire \ram[41][1] ;
   wire \ram[41][0] ;
   wire \ram[40][15] ;
   wire \ram[40][14] ;
   wire \ram[40][13] ;
   wire \ram[40][12] ;
   wire \ram[40][11] ;
   wire \ram[40][10] ;
   wire \ram[40][9] ;
   wire \ram[40][8] ;
   wire \ram[40][7] ;
   wire \ram[40][6] ;
   wire \ram[40][5] ;
   wire \ram[40][4] ;
   wire \ram[40][3] ;
   wire \ram[40][2] ;
   wire \ram[40][1] ;
   wire \ram[40][0] ;
   wire \ram[39][15] ;
   wire \ram[39][14] ;
   wire \ram[39][13] ;
   wire \ram[39][12] ;
   wire \ram[39][11] ;
   wire \ram[39][10] ;
   wire \ram[39][9] ;
   wire \ram[39][8] ;
   wire \ram[39][7] ;
   wire \ram[39][6] ;
   wire \ram[39][5] ;
   wire \ram[39][4] ;
   wire \ram[39][3] ;
   wire \ram[39][2] ;
   wire \ram[39][1] ;
   wire \ram[39][0] ;
   wire \ram[38][15] ;
   wire \ram[38][14] ;
   wire \ram[38][13] ;
   wire \ram[38][12] ;
   wire \ram[38][11] ;
   wire \ram[38][10] ;
   wire \ram[38][9] ;
   wire \ram[38][8] ;
   wire \ram[38][7] ;
   wire \ram[38][6] ;
   wire \ram[38][5] ;
   wire \ram[38][4] ;
   wire \ram[38][3] ;
   wire \ram[38][2] ;
   wire \ram[38][1] ;
   wire \ram[38][0] ;
   wire \ram[37][15] ;
   wire \ram[37][14] ;
   wire \ram[37][13] ;
   wire \ram[37][12] ;
   wire \ram[37][11] ;
   wire \ram[37][10] ;
   wire \ram[37][9] ;
   wire \ram[37][8] ;
   wire \ram[37][7] ;
   wire \ram[37][6] ;
   wire \ram[37][5] ;
   wire \ram[37][4] ;
   wire \ram[37][3] ;
   wire \ram[37][2] ;
   wire \ram[37][1] ;
   wire \ram[37][0] ;
   wire \ram[36][15] ;
   wire \ram[36][14] ;
   wire \ram[36][13] ;
   wire \ram[36][12] ;
   wire \ram[36][11] ;
   wire \ram[36][10] ;
   wire \ram[36][9] ;
   wire \ram[36][8] ;
   wire \ram[36][7] ;
   wire \ram[36][6] ;
   wire \ram[36][5] ;
   wire \ram[36][4] ;
   wire \ram[36][3] ;
   wire \ram[36][2] ;
   wire \ram[36][1] ;
   wire \ram[36][0] ;
   wire \ram[35][15] ;
   wire \ram[35][14] ;
   wire \ram[35][13] ;
   wire \ram[35][12] ;
   wire \ram[35][11] ;
   wire \ram[35][10] ;
   wire \ram[35][9] ;
   wire \ram[35][8] ;
   wire \ram[35][7] ;
   wire \ram[35][6] ;
   wire \ram[35][5] ;
   wire \ram[35][4] ;
   wire \ram[35][3] ;
   wire \ram[35][2] ;
   wire \ram[35][1] ;
   wire \ram[35][0] ;
   wire \ram[34][15] ;
   wire \ram[34][14] ;
   wire \ram[34][13] ;
   wire \ram[34][12] ;
   wire \ram[34][11] ;
   wire \ram[34][10] ;
   wire \ram[34][9] ;
   wire \ram[34][8] ;
   wire \ram[34][7] ;
   wire \ram[34][6] ;
   wire \ram[34][5] ;
   wire \ram[34][4] ;
   wire \ram[34][3] ;
   wire \ram[34][2] ;
   wire \ram[34][1] ;
   wire \ram[34][0] ;
   wire \ram[33][15] ;
   wire \ram[33][14] ;
   wire \ram[33][13] ;
   wire \ram[33][12] ;
   wire \ram[33][11] ;
   wire \ram[33][10] ;
   wire \ram[33][9] ;
   wire \ram[33][8] ;
   wire \ram[33][7] ;
   wire \ram[33][6] ;
   wire \ram[33][5] ;
   wire \ram[33][4] ;
   wire \ram[33][3] ;
   wire \ram[33][2] ;
   wire \ram[33][1] ;
   wire \ram[33][0] ;
   wire \ram[32][15] ;
   wire \ram[32][14] ;
   wire \ram[32][13] ;
   wire \ram[32][12] ;
   wire \ram[32][11] ;
   wire \ram[32][10] ;
   wire \ram[32][9] ;
   wire \ram[32][8] ;
   wire \ram[32][7] ;
   wire \ram[32][6] ;
   wire \ram[32][5] ;
   wire \ram[32][4] ;
   wire \ram[32][3] ;
   wire \ram[32][2] ;
   wire \ram[32][1] ;
   wire \ram[32][0] ;
   wire \ram[31][15] ;
   wire \ram[31][14] ;
   wire \ram[31][13] ;
   wire \ram[31][12] ;
   wire \ram[31][11] ;
   wire \ram[31][10] ;
   wire \ram[31][9] ;
   wire \ram[31][8] ;
   wire \ram[31][7] ;
   wire \ram[31][6] ;
   wire \ram[31][5] ;
   wire \ram[31][4] ;
   wire \ram[31][3] ;
   wire \ram[31][2] ;
   wire \ram[31][1] ;
   wire \ram[31][0] ;
   wire \ram[30][15] ;
   wire \ram[30][14] ;
   wire \ram[30][13] ;
   wire \ram[30][12] ;
   wire \ram[30][11] ;
   wire \ram[30][10] ;
   wire \ram[30][9] ;
   wire \ram[30][8] ;
   wire \ram[30][7] ;
   wire \ram[30][6] ;
   wire \ram[30][5] ;
   wire \ram[30][4] ;
   wire \ram[30][3] ;
   wire \ram[30][2] ;
   wire \ram[30][1] ;
   wire \ram[30][0] ;
   wire \ram[29][15] ;
   wire \ram[29][14] ;
   wire \ram[29][13] ;
   wire \ram[29][12] ;
   wire \ram[29][11] ;
   wire \ram[29][10] ;
   wire \ram[29][9] ;
   wire \ram[29][8] ;
   wire \ram[29][7] ;
   wire \ram[29][6] ;
   wire \ram[29][5] ;
   wire \ram[29][4] ;
   wire \ram[29][3] ;
   wire \ram[29][2] ;
   wire \ram[29][1] ;
   wire \ram[29][0] ;
   wire \ram[28][15] ;
   wire \ram[28][14] ;
   wire \ram[28][13] ;
   wire \ram[28][12] ;
   wire \ram[28][11] ;
   wire \ram[28][10] ;
   wire \ram[28][9] ;
   wire \ram[28][8] ;
   wire \ram[28][7] ;
   wire \ram[28][6] ;
   wire \ram[28][5] ;
   wire \ram[28][4] ;
   wire \ram[28][3] ;
   wire \ram[28][2] ;
   wire \ram[28][1] ;
   wire \ram[28][0] ;
   wire \ram[27][15] ;
   wire \ram[27][14] ;
   wire \ram[27][13] ;
   wire \ram[27][12] ;
   wire \ram[27][11] ;
   wire \ram[27][10] ;
   wire \ram[27][9] ;
   wire \ram[27][8] ;
   wire \ram[27][7] ;
   wire \ram[27][6] ;
   wire \ram[27][5] ;
   wire \ram[27][4] ;
   wire \ram[27][3] ;
   wire \ram[27][2] ;
   wire \ram[27][1] ;
   wire \ram[27][0] ;
   wire \ram[26][15] ;
   wire \ram[26][14] ;
   wire \ram[26][13] ;
   wire \ram[26][12] ;
   wire \ram[26][11] ;
   wire \ram[26][10] ;
   wire \ram[26][9] ;
   wire \ram[26][8] ;
   wire \ram[26][7] ;
   wire \ram[26][6] ;
   wire \ram[26][5] ;
   wire \ram[26][4] ;
   wire \ram[26][3] ;
   wire \ram[26][2] ;
   wire \ram[26][1] ;
   wire \ram[26][0] ;
   wire \ram[25][15] ;
   wire \ram[25][14] ;
   wire \ram[25][13] ;
   wire \ram[25][12] ;
   wire \ram[25][11] ;
   wire \ram[25][10] ;
   wire \ram[25][9] ;
   wire \ram[25][8] ;
   wire \ram[25][7] ;
   wire \ram[25][6] ;
   wire \ram[25][5] ;
   wire \ram[25][4] ;
   wire \ram[25][3] ;
   wire \ram[25][2] ;
   wire \ram[25][1] ;
   wire \ram[25][0] ;
   wire \ram[24][15] ;
   wire \ram[24][14] ;
   wire \ram[24][13] ;
   wire \ram[24][12] ;
   wire \ram[24][11] ;
   wire \ram[24][10] ;
   wire \ram[24][9] ;
   wire \ram[24][8] ;
   wire \ram[24][7] ;
   wire \ram[24][6] ;
   wire \ram[24][5] ;
   wire \ram[24][4] ;
   wire \ram[24][3] ;
   wire \ram[24][2] ;
   wire \ram[24][1] ;
   wire \ram[24][0] ;
   wire \ram[23][15] ;
   wire \ram[23][14] ;
   wire \ram[23][13] ;
   wire \ram[23][12] ;
   wire \ram[23][11] ;
   wire \ram[23][10] ;
   wire \ram[23][9] ;
   wire \ram[23][8] ;
   wire \ram[23][7] ;
   wire \ram[23][6] ;
   wire \ram[23][5] ;
   wire \ram[23][4] ;
   wire \ram[23][3] ;
   wire \ram[23][2] ;
   wire \ram[23][1] ;
   wire \ram[23][0] ;
   wire \ram[22][15] ;
   wire \ram[22][14] ;
   wire \ram[22][13] ;
   wire \ram[22][12] ;
   wire \ram[22][11] ;
   wire \ram[22][10] ;
   wire \ram[22][9] ;
   wire \ram[22][8] ;
   wire \ram[22][7] ;
   wire \ram[22][6] ;
   wire \ram[22][5] ;
   wire \ram[22][4] ;
   wire \ram[22][3] ;
   wire \ram[22][2] ;
   wire \ram[22][1] ;
   wire \ram[22][0] ;
   wire \ram[21][15] ;
   wire \ram[21][14] ;
   wire \ram[21][13] ;
   wire \ram[21][12] ;
   wire \ram[21][11] ;
   wire \ram[21][10] ;
   wire \ram[21][9] ;
   wire \ram[21][8] ;
   wire \ram[21][7] ;
   wire \ram[21][6] ;
   wire \ram[21][5] ;
   wire \ram[21][4] ;
   wire \ram[21][3] ;
   wire \ram[21][2] ;
   wire \ram[21][1] ;
   wire \ram[21][0] ;
   wire \ram[20][15] ;
   wire \ram[20][14] ;
   wire \ram[20][13] ;
   wire \ram[20][12] ;
   wire \ram[20][11] ;
   wire \ram[20][10] ;
   wire \ram[20][9] ;
   wire \ram[20][8] ;
   wire \ram[20][7] ;
   wire \ram[20][6] ;
   wire \ram[20][5] ;
   wire \ram[20][4] ;
   wire \ram[20][3] ;
   wire \ram[20][2] ;
   wire \ram[20][1] ;
   wire \ram[20][0] ;
   wire \ram[19][15] ;
   wire \ram[19][14] ;
   wire \ram[19][13] ;
   wire \ram[19][12] ;
   wire \ram[19][11] ;
   wire \ram[19][10] ;
   wire \ram[19][9] ;
   wire \ram[19][8] ;
   wire \ram[19][7] ;
   wire \ram[19][6] ;
   wire \ram[19][5] ;
   wire \ram[19][4] ;
   wire \ram[19][3] ;
   wire \ram[19][2] ;
   wire \ram[19][1] ;
   wire \ram[19][0] ;
   wire \ram[18][15] ;
   wire \ram[18][14] ;
   wire \ram[18][13] ;
   wire \ram[18][12] ;
   wire \ram[18][11] ;
   wire \ram[18][10] ;
   wire \ram[18][9] ;
   wire \ram[18][8] ;
   wire \ram[18][7] ;
   wire \ram[18][6] ;
   wire \ram[18][5] ;
   wire \ram[18][4] ;
   wire \ram[18][3] ;
   wire \ram[18][2] ;
   wire \ram[18][1] ;
   wire \ram[18][0] ;
   wire \ram[17][15] ;
   wire \ram[17][14] ;
   wire \ram[17][13] ;
   wire \ram[17][12] ;
   wire \ram[17][11] ;
   wire \ram[17][10] ;
   wire \ram[17][9] ;
   wire \ram[17][8] ;
   wire \ram[17][7] ;
   wire \ram[17][6] ;
   wire \ram[17][5] ;
   wire \ram[17][4] ;
   wire \ram[17][3] ;
   wire \ram[17][2] ;
   wire \ram[17][1] ;
   wire \ram[17][0] ;
   wire \ram[16][15] ;
   wire \ram[16][14] ;
   wire \ram[16][13] ;
   wire \ram[16][12] ;
   wire \ram[16][11] ;
   wire \ram[16][10] ;
   wire \ram[16][9] ;
   wire \ram[16][8] ;
   wire \ram[16][7] ;
   wire \ram[16][6] ;
   wire \ram[16][5] ;
   wire \ram[16][4] ;
   wire \ram[16][3] ;
   wire \ram[16][2] ;
   wire \ram[16][1] ;
   wire \ram[16][0] ;
   wire \ram[15][15] ;
   wire \ram[15][14] ;
   wire \ram[15][13] ;
   wire \ram[15][12] ;
   wire \ram[15][11] ;
   wire \ram[15][10] ;
   wire \ram[15][9] ;
   wire \ram[15][8] ;
   wire \ram[15][7] ;
   wire \ram[15][6] ;
   wire \ram[15][5] ;
   wire \ram[15][4] ;
   wire \ram[15][3] ;
   wire \ram[15][2] ;
   wire \ram[15][1] ;
   wire \ram[15][0] ;
   wire \ram[14][15] ;
   wire \ram[14][14] ;
   wire \ram[14][13] ;
   wire \ram[14][12] ;
   wire \ram[14][11] ;
   wire \ram[14][10] ;
   wire \ram[14][9] ;
   wire \ram[14][8] ;
   wire \ram[14][7] ;
   wire \ram[14][6] ;
   wire \ram[14][5] ;
   wire \ram[14][4] ;
   wire \ram[14][3] ;
   wire \ram[14][2] ;
   wire \ram[14][1] ;
   wire \ram[14][0] ;
   wire \ram[13][15] ;
   wire \ram[13][14] ;
   wire \ram[13][13] ;
   wire \ram[13][12] ;
   wire \ram[13][11] ;
   wire \ram[13][10] ;
   wire \ram[13][9] ;
   wire \ram[13][8] ;
   wire \ram[13][7] ;
   wire \ram[13][6] ;
   wire \ram[13][5] ;
   wire \ram[13][4] ;
   wire \ram[13][3] ;
   wire \ram[13][2] ;
   wire \ram[13][1] ;
   wire \ram[13][0] ;
   wire \ram[12][15] ;
   wire \ram[12][14] ;
   wire \ram[12][13] ;
   wire \ram[12][12] ;
   wire \ram[12][11] ;
   wire \ram[12][10] ;
   wire \ram[12][9] ;
   wire \ram[12][8] ;
   wire \ram[12][7] ;
   wire \ram[12][6] ;
   wire \ram[12][5] ;
   wire \ram[12][4] ;
   wire \ram[12][3] ;
   wire \ram[12][2] ;
   wire \ram[12][1] ;
   wire \ram[12][0] ;
   wire \ram[11][15] ;
   wire \ram[11][14] ;
   wire \ram[11][13] ;
   wire \ram[11][12] ;
   wire \ram[11][11] ;
   wire \ram[11][10] ;
   wire \ram[11][9] ;
   wire \ram[11][8] ;
   wire \ram[11][7] ;
   wire \ram[11][6] ;
   wire \ram[11][5] ;
   wire \ram[11][4] ;
   wire \ram[11][3] ;
   wire \ram[11][2] ;
   wire \ram[11][1] ;
   wire \ram[11][0] ;
   wire \ram[10][15] ;
   wire \ram[10][14] ;
   wire \ram[10][13] ;
   wire \ram[10][12] ;
   wire \ram[10][11] ;
   wire \ram[10][10] ;
   wire \ram[10][9] ;
   wire \ram[10][8] ;
   wire \ram[10][7] ;
   wire \ram[10][6] ;
   wire \ram[10][5] ;
   wire \ram[10][4] ;
   wire \ram[10][3] ;
   wire \ram[10][2] ;
   wire \ram[10][1] ;
   wire \ram[10][0] ;
   wire \ram[9][15] ;
   wire \ram[9][14] ;
   wire \ram[9][13] ;
   wire \ram[9][12] ;
   wire \ram[9][11] ;
   wire \ram[9][10] ;
   wire \ram[9][9] ;
   wire \ram[9][8] ;
   wire \ram[9][7] ;
   wire \ram[9][6] ;
   wire \ram[9][5] ;
   wire \ram[9][4] ;
   wire \ram[9][3] ;
   wire \ram[9][2] ;
   wire \ram[9][1] ;
   wire \ram[9][0] ;
   wire \ram[8][15] ;
   wire \ram[8][14] ;
   wire \ram[8][13] ;
   wire \ram[8][12] ;
   wire \ram[8][11] ;
   wire \ram[8][10] ;
   wire \ram[8][9] ;
   wire \ram[8][8] ;
   wire \ram[8][7] ;
   wire \ram[8][6] ;
   wire \ram[8][5] ;
   wire \ram[8][4] ;
   wire \ram[8][3] ;
   wire \ram[8][2] ;
   wire \ram[8][1] ;
   wire \ram[8][0] ;
   wire \ram[7][15] ;
   wire \ram[7][14] ;
   wire \ram[7][13] ;
   wire \ram[7][12] ;
   wire \ram[7][11] ;
   wire \ram[7][10] ;
   wire \ram[7][9] ;
   wire \ram[7][8] ;
   wire \ram[7][7] ;
   wire \ram[7][6] ;
   wire \ram[7][5] ;
   wire \ram[7][4] ;
   wire \ram[7][3] ;
   wire \ram[7][2] ;
   wire \ram[7][1] ;
   wire \ram[7][0] ;
   wire \ram[6][15] ;
   wire \ram[6][14] ;
   wire \ram[6][13] ;
   wire \ram[6][12] ;
   wire \ram[6][11] ;
   wire \ram[6][10] ;
   wire \ram[6][9] ;
   wire \ram[6][8] ;
   wire \ram[6][7] ;
   wire \ram[6][6] ;
   wire \ram[6][5] ;
   wire \ram[6][4] ;
   wire \ram[6][3] ;
   wire \ram[6][2] ;
   wire \ram[6][1] ;
   wire \ram[6][0] ;
   wire \ram[5][15] ;
   wire \ram[5][14] ;
   wire \ram[5][13] ;
   wire \ram[5][12] ;
   wire \ram[5][11] ;
   wire \ram[5][10] ;
   wire \ram[5][9] ;
   wire \ram[5][8] ;
   wire \ram[5][7] ;
   wire \ram[5][6] ;
   wire \ram[5][5] ;
   wire \ram[5][4] ;
   wire \ram[5][3] ;
   wire \ram[5][2] ;
   wire \ram[5][1] ;
   wire \ram[5][0] ;
   wire \ram[4][15] ;
   wire \ram[4][14] ;
   wire \ram[4][13] ;
   wire \ram[4][12] ;
   wire \ram[4][11] ;
   wire \ram[4][10] ;
   wire \ram[4][9] ;
   wire \ram[4][8] ;
   wire \ram[4][7] ;
   wire \ram[4][6] ;
   wire \ram[4][5] ;
   wire \ram[4][4] ;
   wire \ram[4][3] ;
   wire \ram[4][2] ;
   wire \ram[4][1] ;
   wire \ram[4][0] ;
   wire \ram[3][15] ;
   wire \ram[3][14] ;
   wire \ram[3][13] ;
   wire \ram[3][12] ;
   wire \ram[3][11] ;
   wire \ram[3][10] ;
   wire \ram[3][9] ;
   wire \ram[3][8] ;
   wire \ram[3][7] ;
   wire \ram[3][6] ;
   wire \ram[3][5] ;
   wire \ram[3][4] ;
   wire \ram[3][3] ;
   wire \ram[3][2] ;
   wire \ram[3][1] ;
   wire \ram[3][0] ;
   wire \ram[2][15] ;
   wire \ram[2][14] ;
   wire \ram[2][13] ;
   wire \ram[2][12] ;
   wire \ram[2][11] ;
   wire \ram[2][10] ;
   wire \ram[2][9] ;
   wire \ram[2][8] ;
   wire \ram[2][7] ;
   wire \ram[2][6] ;
   wire \ram[2][5] ;
   wire \ram[2][4] ;
   wire \ram[2][3] ;
   wire \ram[2][2] ;
   wire \ram[2][1] ;
   wire \ram[2][0] ;
   wire \ram[1][15] ;
   wire \ram[1][14] ;
   wire \ram[1][13] ;
   wire \ram[1][12] ;
   wire \ram[1][11] ;
   wire \ram[1][10] ;
   wire \ram[1][9] ;
   wire \ram[1][8] ;
   wire \ram[1][7] ;
   wire \ram[1][6] ;
   wire \ram[1][5] ;
   wire \ram[1][4] ;
   wire \ram[1][3] ;
   wire \ram[1][2] ;
   wire \ram[1][1] ;
   wire \ram[1][0] ;
   wire \ram[0][15] ;
   wire \ram[0][14] ;
   wire \ram[0][13] ;
   wire \ram[0][12] ;
   wire \ram[0][11] ;
   wire \ram[0][10] ;
   wire \ram[0][9] ;
   wire \ram[0][8] ;
   wire \ram[0][7] ;
   wire \ram[0][6] ;
   wire \ram[0][5] ;
   wire \ram[0][4] ;
   wire \ram[0][3] ;
   wire \ram[0][2] ;
   wire \ram[0][1] ;
   wire \ram[0][0] ;
   wire N4126;
   wire N4127;
   wire N4128;
   wire N4129;
   wire N4130;
   wire N4131;
   wire N4132;
   wire N4133;
   wire N4134;
   wire N4135;
   wire N4136;
   wire N4137;
   wire N4138;
   wire N4139;
   wire N4140;
   wire N4141;
   wire n6;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n27;
   wire n30;
   wire n33;
   wire n36;
   wire n39;
   wire n42;
   wire n45;
   wire n48;
   wire n51;
   wire n54;
   wire n57;
   wire n60;
   wire n63;
   wire n66;
   wire n69;
   wire n71;
   wire n72;
   wire n74;
   wire n77;
   wire n79;
   wire n81;
   wire n83;
   wire n85;
   wire n87;
   wire n89;
   wire n91;
   wire n93;
   wire n95;
   wire n97;
   wire n99;
   wire n101;
   wire n103;
   wire n105;
   wire n106;
   wire n108;
   wire n111;
   wire n113;
   wire n115;
   wire n117;
   wire n119;
   wire n121;
   wire n123;
   wire n125;
   wire n127;
   wire n129;
   wire n131;
   wire n133;
   wire n135;
   wire n137;
   wire n139;
   wire n140;
   wire n142;
   wire n145;
   wire n147;
   wire n149;
   wire n151;
   wire n153;
   wire n155;
   wire n157;
   wire n159;
   wire n161;
   wire n163;
   wire n165;
   wire n167;
   wire n169;
   wire n171;
   wire n173;
   wire n174;
   wire n176;
   wire n179;
   wire n181;
   wire n183;
   wire n185;
   wire n187;
   wire n189;
   wire n191;
   wire n193;
   wire n195;
   wire n197;
   wire n199;
   wire n201;
   wire n203;
   wire n205;
   wire n207;
   wire n208;
   wire n210;
   wire n213;
   wire n215;
   wire n217;
   wire n219;
   wire n221;
   wire n223;
   wire n225;
   wire n227;
   wire n229;
   wire n231;
   wire n233;
   wire n235;
   wire n237;
   wire n239;
   wire n241;
   wire n243;
   wire n246;
   wire n248;
   wire n250;
   wire n252;
   wire n254;
   wire n256;
   wire n258;
   wire n260;
   wire n262;
   wire n264;
   wire n266;
   wire n268;
   wire n270;
   wire n272;
   wire n274;
   wire n276;
   wire n279;
   wire n281;
   wire n283;
   wire n285;
   wire n287;
   wire n289;
   wire n291;
   wire n293;
   wire n295;
   wire n297;
   wire n299;
   wire n301;
   wire n303;
   wire n305;
   wire n307;
   wire n309;
   wire n312;
   wire n314;
   wire n316;
   wire n318;
   wire n320;
   wire n322;
   wire n324;
   wire n326;
   wire n328;
   wire n330;
   wire n332;
   wire n334;
   wire n336;
   wire n338;
   wire n340;
   wire n341;
   wire n343;
   wire n346;
   wire n348;
   wire n350;
   wire n352;
   wire n354;
   wire n356;
   wire n358;
   wire n360;
   wire n362;
   wire n364;
   wire n366;
   wire n368;
   wire n370;
   wire n372;
   wire n374;
   wire n376;
   wire n379;
   wire n381;
   wire n383;
   wire n385;
   wire n387;
   wire n389;
   wire n391;
   wire n393;
   wire n395;
   wire n397;
   wire n399;
   wire n401;
   wire n403;
   wire n405;
   wire n407;
   wire n409;
   wire n412;
   wire n414;
   wire n416;
   wire n418;
   wire n420;
   wire n422;
   wire n424;
   wire n426;
   wire n428;
   wire n430;
   wire n432;
   wire n434;
   wire n436;
   wire n438;
   wire n440;
   wire n442;
   wire n445;
   wire n447;
   wire n449;
   wire n451;
   wire n453;
   wire n455;
   wire n457;
   wire n459;
   wire n461;
   wire n463;
   wire n465;
   wire n467;
   wire n469;
   wire n471;
   wire n473;
   wire n474;
   wire n476;
   wire n479;
   wire n481;
   wire n483;
   wire n485;
   wire n487;
   wire n489;
   wire n491;
   wire n493;
   wire n495;
   wire n497;
   wire n499;
   wire n501;
   wire n503;
   wire n505;
   wire n507;
   wire n509;
   wire n512;
   wire n514;
   wire n516;
   wire n518;
   wire n520;
   wire n522;
   wire n524;
   wire n526;
   wire n528;
   wire n530;
   wire n532;
   wire n534;
   wire n536;
   wire n538;
   wire n540;
   wire n542;
   wire n544;
   wire n545;
   wire n547;
   wire n548;
   wire n550;
   wire n551;
   wire n553;
   wire n554;
   wire n556;
   wire n557;
   wire n559;
   wire n561;
   wire n563;
   wire n565;
   wire n566;
   wire n568;
   wire n570;
   wire n572;
   wire n574;
   wire n575;
   wire n577;
   wire n579;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3297;
   wire n3298;
   wire n3299;
   wire n3300;
   wire n3301;
   wire n3302;
   wire n3303;
   wire n3304;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire n3330;
   wire n3331;
   wire n3332;
   wire n3333;
   wire n3334;
   wire n3335;
   wire n3336;
   wire n3337;
   wire n3338;
   wire n3339;
   wire n3340;
   wire n3341;
   wire n3342;
   wire n3343;
   wire n3344;
   wire n3345;
   wire n3346;
   wire n3347;
   wire n3348;
   wire n3349;
   wire n3350;
   wire n3351;
   wire n3352;
   wire n3353;
   wire n3354;
   wire n3355;
   wire n3356;
   wire n3357;
   wire n3358;
   wire n3359;
   wire n3360;
   wire n3361;
   wire n3362;
   wire n3363;
   wire n3364;
   wire n3365;
   wire n3366;
   wire n3367;
   wire n3368;
   wire n3369;
   wire n3370;
   wire n3371;
   wire n3372;
   wire n3373;
   wire n3374;
   wire n3375;
   wire n3376;
   wire n3377;
   wire n3378;
   wire n3379;
   wire n3380;
   wire n3381;
   wire n3382;
   wire n3383;
   wire n3384;
   wire n3385;
   wire n3386;
   wire n3387;
   wire n3388;
   wire n3389;
   wire n3390;
   wire n3391;
   wire n3392;
   wire n3393;
   wire n3394;
   wire n3395;
   wire n3396;
   wire n3397;
   wire n3398;
   wire n3399;
   wire n3400;
   wire n3401;
   wire n3402;
   wire n3403;
   wire n3404;
   wire n3405;
   wire n3406;
   wire n3407;
   wire n3408;
   wire n3409;
   wire n3410;
   wire n3411;
   wire n3412;
   wire n3413;
   wire n3414;
   wire n3415;
   wire n3416;
   wire n3417;
   wire n3418;
   wire n3419;
   wire n3420;
   wire n3421;
   wire n3422;
   wire n3423;
   wire n3424;
   wire n3425;
   wire n3426;
   wire n3427;
   wire n3428;
   wire n3429;
   wire n3430;
   wire n3431;
   wire n3432;
   wire n3433;
   wire n3434;
   wire n3435;
   wire n3436;
   wire n3437;
   wire n3438;
   wire n3439;
   wire n3440;
   wire n3441;
   wire n3442;
   wire n3443;
   wire n3444;
   wire n3445;
   wire n3446;
   wire n3447;
   wire n3448;
   wire n3449;
   wire n3450;
   wire n3451;
   wire n3452;
   wire n3453;
   wire n3454;
   wire n3455;
   wire n3456;
   wire n3457;
   wire n3458;
   wire n3459;
   wire n3460;
   wire n3461;
   wire n3462;
   wire n3463;
   wire n3464;
   wire n3465;
   wire n3466;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3475;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3485;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3589;
   wire n3590;
   wire n3591;
   wire n3592;
   wire n3593;
   wire n3594;
   wire n3595;
   wire n3596;
   wire n3597;
   wire n3598;
   wire n3599;
   wire n3600;
   wire n3601;
   wire n3602;
   wire n3603;
   wire n3604;
   wire n3605;
   wire n3606;
   wire n3607;
   wire n3608;
   wire n3609;
   wire n3610;
   wire n3611;
   wire n3612;
   wire n3613;
   wire n3614;
   wire n3615;
   wire n3616;
   wire n3617;
   wire n3618;
   wire n3619;
   wire n3620;
   wire n3621;
   wire n3622;
   wire n3623;
   wire n3624;
   wire n3625;
   wire n3626;
   wire n3627;
   wire n3628;
   wire n3629;
   wire n3630;
   wire n3631;
   wire n3632;
   wire n3633;
   wire n3634;
   wire n3635;
   wire n3636;
   wire n3637;
   wire n3638;
   wire n3639;
   wire n3640;
   wire n3641;
   wire n3642;
   wire n3643;
   wire n3644;
   wire n3645;
   wire n3646;
   wire n3647;
   wire n3648;
   wire n3649;
   wire n3650;
   wire n3651;
   wire n3652;
   wire n3653;
   wire n3654;
   wire n3655;
   wire n3656;
   wire n3657;
   wire n3658;
   wire n3659;
   wire n3660;
   wire n3661;
   wire n3662;
   wire n3663;
   wire n3664;
   wire n3665;
   wire n3666;
   wire n3667;
   wire n3668;
   wire n3669;
   wire n3670;
   wire n3671;
   wire n3672;
   wire n3673;
   wire n3674;
   wire n3675;
   wire n3676;
   wire n3677;
   wire n3678;
   wire n3679;
   wire n3680;
   wire n3681;
   wire n3682;
   wire n3683;
   wire n3684;
   wire n3685;
   wire n3686;
   wire n3687;
   wire n3688;
   wire n3689;
   wire n3690;
   wire n3691;
   wire n3692;
   wire n3693;
   wire n3694;
   wire n3695;
   wire n3696;
   wire n3697;
   wire n3698;
   wire n3699;
   wire n3700;
   wire n3701;
   wire n3702;
   wire n3703;
   wire n3704;
   wire n3705;
   wire n3706;
   wire n3707;
   wire n3708;
   wire n3709;
   wire n3710;
   wire n3711;
   wire n3712;
   wire n3713;
   wire n3714;
   wire n3715;
   wire n3716;
   wire n3717;
   wire n3718;
   wire n3719;
   wire n3720;
   wire n3721;
   wire n3722;
   wire n3723;
   wire n3724;
   wire n3725;
   wire n3726;
   wire n3727;
   wire n3728;
   wire n3729;
   wire n3730;
   wire n3731;
   wire n3732;
   wire n3733;
   wire n3734;
   wire n3735;
   wire n3736;
   wire n3737;
   wire n3738;
   wire n3739;
   wire n3740;
   wire n3741;
   wire n3742;
   wire n3743;
   wire n3744;
   wire n3745;
   wire n3746;
   wire n3747;
   wire n3748;
   wire n3749;
   wire n3750;
   wire n3751;
   wire n3752;
   wire n3753;
   wire n3754;
   wire n3755;
   wire n3756;
   wire n3757;
   wire n3758;
   wire n3759;
   wire n3760;
   wire n3761;
   wire n3762;
   wire n3763;
   wire n3764;
   wire n3765;
   wire n3766;
   wire n3767;
   wire n3768;
   wire n3769;
   wire n3770;
   wire n3771;
   wire n3772;
   wire n3773;
   wire n3774;
   wire n3775;
   wire n3776;
   wire n3777;
   wire n3778;
   wire n3779;
   wire n3780;
   wire n3781;
   wire n3782;
   wire n3783;
   wire n3784;
   wire n3785;
   wire n3786;
   wire n3787;
   wire n3788;
   wire n3789;
   wire n3790;
   wire n3791;
   wire n3792;
   wire n3793;
   wire n3794;
   wire n3795;
   wire n3796;
   wire n3797;
   wire n3798;
   wire n3799;
   wire n3800;
   wire n3801;
   wire n3802;
   wire n3803;
   wire n3804;
   wire n3805;
   wire n3806;
   wire n3807;
   wire n3808;
   wire n3809;
   wire n3810;
   wire n3811;
   wire n3812;
   wire n3813;
   wire n3814;
   wire n3815;
   wire n3816;
   wire n3817;
   wire n3818;
   wire n3819;
   wire n3820;
   wire n3821;
   wire n3822;
   wire n3823;
   wire n3824;
   wire n3825;
   wire n3826;
   wire n3827;
   wire n3828;
   wire n3829;
   wire n3830;
   wire n3831;
   wire n3832;
   wire n3833;
   wire n3834;
   wire n3835;
   wire n3836;
   wire n3837;
   wire n3838;
   wire n3839;
   wire n3840;
   wire n3841;
   wire n3842;
   wire n3843;
   wire n3844;
   wire n3845;
   wire n3846;
   wire n3847;
   wire n3848;
   wire n3849;
   wire n3850;
   wire n3851;
   wire n3852;
   wire n3853;
   wire n3854;
   wire n3855;
   wire n3856;
   wire n3857;
   wire n3858;
   wire n3859;
   wire n3860;
   wire n3861;
   wire n3862;
   wire n3863;
   wire n3864;
   wire n3865;
   wire n3866;
   wire n3867;
   wire n3868;
   wire n3869;
   wire n3870;
   wire n3871;
   wire n3872;
   wire n3873;
   wire n3874;
   wire n3875;
   wire n3876;
   wire n3877;
   wire n3878;
   wire n3879;
   wire n3880;
   wire n3881;
   wire n3882;
   wire n3883;
   wire n3884;
   wire n3885;
   wire n3886;
   wire n3887;
   wire n3888;
   wire n3889;
   wire n3890;
   wire n3891;
   wire n3892;
   wire n3893;
   wire n3894;
   wire n3895;
   wire n3896;
   wire n3897;
   wire n3898;
   wire n3899;
   wire n3900;
   wire n3901;
   wire n3902;
   wire n3903;
   wire n3904;
   wire n3905;
   wire n3906;
   wire n3907;
   wire n3908;
   wire n3909;
   wire n3910;
   wire n3911;
   wire n3912;
   wire n3913;
   wire n3914;
   wire n3915;
   wire n3916;
   wire n3917;
   wire n3918;
   wire n3919;
   wire n3920;
   wire n3921;
   wire n3922;
   wire n3923;
   wire n3924;
   wire n3925;
   wire n3926;
   wire n3927;
   wire n3928;
   wire n3929;
   wire n3930;
   wire n3931;
   wire n3932;
   wire n3933;
   wire n3934;
   wire n3935;
   wire n3936;
   wire n3937;
   wire n3938;
   wire n3939;
   wire n3940;
   wire n3941;
   wire n3942;
   wire n3943;
   wire n3944;
   wire n3945;
   wire n3946;
   wire n3947;
   wire n3948;
   wire n3949;
   wire n3950;
   wire n3951;
   wire n3952;
   wire n3953;
   wire n3954;
   wire n3955;
   wire n3956;
   wire n3957;
   wire n3958;
   wire n3959;
   wire n3960;
   wire n3961;
   wire n3962;
   wire n3963;
   wire n3964;
   wire n3965;
   wire n3966;
   wire n3967;
   wire n3968;
   wire n3969;
   wire n3970;
   wire n3971;
   wire n3972;
   wire n3973;
   wire n3974;
   wire n3975;
   wire n3976;
   wire n3977;
   wire n3978;
   wire n3979;
   wire n3980;
   wire n3981;
   wire n3982;
   wire n3983;
   wire n3984;
   wire n3985;
   wire n3986;
   wire n3987;
   wire n3988;
   wire n3989;
   wire n3990;
   wire n3991;
   wire n3992;
   wire n3993;
   wire n3994;
   wire n3995;
   wire n3996;
   wire n3997;
   wire n3998;
   wire n3999;
   wire n4000;
   wire n4001;
   wire n4002;
   wire n4003;
   wire n4004;
   wire n4005;
   wire n4006;
   wire n4007;
   wire n4008;
   wire n4009;
   wire n4010;
   wire n4011;
   wire n4012;
   wire n4013;
   wire n4014;
   wire n4015;
   wire n4016;
   wire n4017;
   wire n4018;
   wire n4019;
   wire n4020;
   wire n4021;
   wire n4022;
   wire n4023;
   wire n4024;
   wire n4025;
   wire n4026;
   wire n4027;
   wire n4028;
   wire n4029;
   wire n4030;
   wire n4031;
   wire n4032;
   wire n4033;
   wire n4034;
   wire n4035;
   wire n4036;
   wire n4037;
   wire n4038;
   wire n4039;
   wire n4040;
   wire n4041;
   wire n4042;
   wire n4043;
   wire n4044;
   wire n4045;
   wire n4046;
   wire n4047;
   wire n4048;
   wire n4049;
   wire n4050;
   wire n4051;
   wire n4052;
   wire n4053;
   wire n4054;
   wire n4055;
   wire n4056;
   wire n4057;
   wire n4058;
   wire n4059;
   wire n4060;
   wire n4061;
   wire n4062;
   wire n4063;
   wire n4064;
   wire n4065;
   wire n4066;
   wire n4067;
   wire n4068;
   wire n4069;
   wire n4070;
   wire n4071;
   wire n4072;
   wire n4073;
   wire n4074;
   wire n4075;
   wire n4076;
   wire n4077;
   wire n4078;
   wire n4079;
   wire n4080;
   wire n4081;
   wire n4082;
   wire n4083;
   wire n4084;
   wire n4085;
   wire n4086;
   wire n4087;
   wire n4088;
   wire n4089;
   wire n4090;
   wire n4091;
   wire n4092;
   wire n4093;
   wire n4094;
   wire n4095;
   wire n4096;
   wire n4097;
   wire n4098;
   wire n4099;
   wire n4100;
   wire n4101;
   wire n4102;
   wire n4103;
   wire n4104;
   wire n4105;
   wire n4106;
   wire n4107;
   wire n4108;
   wire n4109;
   wire n4110;
   wire n4111;
   wire n4112;
   wire n4113;
   wire n4114;
   wire n4115;
   wire n4116;
   wire n4117;
   wire n4118;
   wire n4119;
   wire n4120;
   wire n4121;
   wire n4122;
   wire n4123;
   wire n4124;
   wire n4125;
   wire n4126;
   wire n4127;
   wire n4128;
   wire n4129;
   wire n4130;
   wire n4131;
   wire n4132;
   wire n4133;
   wire n4134;
   wire n4135;
   wire n4136;
   wire n4137;
   wire n4138;
   wire n4139;
   wire n4140;
   wire n4141;
   wire n4142;
   wire n4143;
   wire n4144;
   wire n4145;
   wire n4146;
   wire n4147;
   wire n4148;
   wire n4149;
   wire n4150;
   wire n4151;
   wire n4152;
   wire n4153;
   wire n4154;
   wire n4155;
   wire n4156;
   wire n4157;
   wire n4158;
   wire n4159;
   wire n4160;
   wire n4161;
   wire n4162;
   wire n4163;
   wire n4164;
   wire n4165;
   wire n4166;
   wire n4167;
   wire n4168;
   wire n4169;
   wire n4170;
   wire n4171;
   wire n4172;
   wire n4173;
   wire n4174;
   wire n4175;
   wire n4176;
   wire n4177;
   wire n4178;
   wire n4179;
   wire n4180;
   wire n4181;
   wire n4182;
   wire n4183;
   wire n4184;
   wire n4185;
   wire n4186;
   wire n4187;
   wire n4188;
   wire n4189;
   wire n4190;
   wire n4191;
   wire n4192;
   wire n4193;
   wire n4194;
   wire n4195;
   wire n4196;
   wire n4197;
   wire n4198;
   wire n4199;
   wire n4200;
   wire n4201;
   wire n4202;
   wire n4203;
   wire n4204;
   wire n4205;
   wire n4206;
   wire n4207;
   wire n4208;
   wire n4209;
   wire n4210;
   wire n4211;
   wire n4212;
   wire n4213;
   wire n4214;
   wire n4215;
   wire n4216;
   wire n4217;
   wire n4218;
   wire n4219;
   wire n4220;
   wire n4221;
   wire n4222;
   wire n4223;
   wire n4224;
   wire n4225;
   wire n4226;
   wire n4227;
   wire n4228;
   wire n4229;
   wire n4230;
   wire n4231;
   wire n4232;
   wire n4233;
   wire n4234;
   wire n4235;
   wire n4236;
   wire n4237;
   wire n4238;
   wire n4239;
   wire n4240;
   wire n4241;
   wire n4242;
   wire n4243;
   wire n4244;
   wire n4245;
   wire n4246;
   wire n4247;
   wire n4248;
   wire n4249;
   wire n4250;
   wire n4251;
   wire n4252;
   wire n4253;
   wire n4254;
   wire n4255;
   wire n4256;
   wire n4257;
   wire n4258;
   wire n4259;
   wire n4260;
   wire n4261;
   wire n4262;
   wire n4263;
   wire n4264;
   wire n4265;
   wire n4266;
   wire n4267;
   wire n4268;
   wire n4269;
   wire n4270;
   wire n4271;
   wire n4272;
   wire n4273;
   wire n4274;
   wire n4275;
   wire n4276;
   wire n4277;
   wire n4278;
   wire n4279;
   wire n4280;
   wire n4281;
   wire n4282;
   wire n4283;
   wire n4284;
   wire n4285;
   wire n4286;
   wire n4287;
   wire n4288;
   wire n4289;
   wire n4290;
   wire n4291;
   wire n4292;
   wire n4293;
   wire n4294;
   wire n4295;
   wire n4296;
   wire n4297;
   wire n4298;
   wire n4299;
   wire n4300;
   wire n4301;
   wire n4302;
   wire n4303;
   wire n4304;
   wire n4305;
   wire n4306;
   wire n4307;
   wire n4308;
   wire n4309;
   wire n4310;
   wire n4311;
   wire n4312;
   wire n4313;
   wire n4314;
   wire n4315;
   wire n4316;
   wire n4317;
   wire n4318;
   wire n4319;
   wire n4320;
   wire n4321;
   wire n4322;
   wire n4323;
   wire n4324;
   wire n4325;
   wire n4326;
   wire n4327;
   wire n4328;
   wire n4329;
   wire n4330;
   wire n4331;
   wire n4332;
   wire n4333;
   wire n4334;
   wire n4335;
   wire n4336;
   wire n4337;
   wire n4338;
   wire n4339;
   wire n4340;
   wire n4341;
   wire n4342;
   wire n4343;
   wire n4344;
   wire n4345;
   wire n4346;
   wire n4347;
   wire n4348;
   wire n4349;
   wire n4350;
   wire n4351;
   wire n4352;
   wire n4353;
   wire n4354;
   wire n4355;
   wire n4356;
   wire n4357;
   wire n4358;
   wire n4359;
   wire n4360;
   wire n4361;
   wire n4362;
   wire n4363;
   wire n4364;
   wire n4365;
   wire n4366;
   wire n4367;
   wire n4368;
   wire n4369;
   wire n4370;
   wire n4371;
   wire n4372;
   wire n4373;
   wire n4374;
   wire n4375;
   wire n4376;
   wire n4377;
   wire n4378;
   wire n4379;
   wire n4380;
   wire n4381;
   wire n4382;
   wire n4383;
   wire n4384;
   wire n4385;
   wire n4386;
   wire n4387;
   wire n4388;
   wire n4389;
   wire n4390;
   wire n4391;
   wire n4392;
   wire n4393;
   wire n4394;
   wire n4395;
   wire n4396;
   wire n4397;
   wire n4398;
   wire n4399;
   wire n4400;
   wire n4401;
   wire n4402;
   wire n4403;
   wire n4404;
   wire n4405;
   wire n4406;
   wire n4407;
   wire n4408;
   wire n4409;
   wire n4410;
   wire n4411;
   wire n4412;
   wire n4413;
   wire n4414;
   wire n4415;
   wire n4416;
   wire n4417;
   wire n4418;
   wire n4419;
   wire n4420;
   wire n4421;
   wire n4422;
   wire n4423;
   wire n4424;
   wire n4425;
   wire n4426;
   wire n4427;
   wire n4428;
   wire n4429;
   wire n4430;
   wire n4431;
   wire n4432;
   wire n4433;
   wire n4434;
   wire n4435;
   wire n4436;
   wire n4437;
   wire n4438;
   wire n4439;
   wire n4440;
   wire n4441;
   wire n4442;
   wire n4443;
   wire n4444;
   wire n4445;
   wire n4446;
   wire n4447;
   wire n4448;
   wire n4449;
   wire n4450;
   wire n4451;
   wire n4452;
   wire n4453;
   wire n4454;
   wire n4455;
   wire n4456;
   wire n4457;
   wire n4458;
   wire n4459;
   wire n4460;
   wire n4461;
   wire n4462;
   wire n4463;
   wire n4464;
   wire n4465;
   wire n4466;
   wire n4467;
   wire n4468;
   wire n4469;
   wire n4470;
   wire n4471;
   wire n4472;
   wire n4473;
   wire n4474;
   wire n4475;
   wire n4476;
   wire n4477;
   wire n4478;
   wire n4479;
   wire n4480;
   wire n4481;
   wire n4482;
   wire n4483;
   wire n4484;
   wire n4485;
   wire n4486;
   wire n4487;
   wire n4488;
   wire n4489;
   wire n4490;
   wire n4491;
   wire n4492;
   wire n4493;
   wire n4494;
   wire n4495;
   wire n4496;
   wire n4497;
   wire n4498;
   wire n4499;
   wire n4500;
   wire n4501;
   wire n4502;
   wire n4503;
   wire n4504;
   wire n4505;
   wire n4506;
   wire n4507;
   wire n4508;
   wire n4509;
   wire n4510;
   wire n4511;
   wire n4512;
   wire n4513;
   wire n4514;
   wire n4515;
   wire n4516;
   wire n4517;
   wire n4518;
   wire n4519;
   wire n4520;
   wire n4521;
   wire n4522;
   wire n4523;
   wire n4524;
   wire n4525;
   wire n4526;
   wire n4527;
   wire n4528;
   wire n4529;
   wire n4530;
   wire n4531;
   wire n4532;
   wire n4533;
   wire n4534;
   wire n4535;
   wire n4536;
   wire n4537;
   wire n4538;
   wire n4539;
   wire n4540;
   wire n4541;
   wire n4542;
   wire n4543;
   wire n4544;
   wire n4545;
   wire n4546;
   wire n4547;
   wire n4548;
   wire n4549;
   wire n4550;
   wire n4551;
   wire n4552;
   wire n4553;
   wire n4554;
   wire n4555;
   wire n4556;
   wire n4557;
   wire n4558;
   wire n4559;
   wire n4560;
   wire n4561;
   wire n4562;
   wire n4563;
   wire n4564;
   wire n4565;
   wire n4566;
   wire n4567;
   wire n4568;
   wire n4569;
   wire n4570;
   wire n4571;
   wire n4572;
   wire n4573;
   wire n4574;
   wire n4575;
   wire n4576;
   wire n4577;
   wire n4578;
   wire n4579;
   wire n4580;
   wire n4581;
   wire n4582;
   wire n4583;
   wire n4584;
   wire n4585;
   wire n4586;
   wire n4587;
   wire n4588;
   wire n4589;
   wire n4590;
   wire n4591;
   wire n4592;
   wire n4593;
   wire n4594;
   wire n4595;
   wire n4596;
   wire n4597;
   wire n4598;
   wire n4599;
   wire n4600;
   wire n4601;
   wire n4602;
   wire n4603;
   wire n4604;
   wire n4605;
   wire n4606;
   wire n4607;
   wire n4608;
   wire n4609;
   wire n4610;
   wire n4611;
   wire n4612;
   wire n4613;
   wire n4614;
   wire n4615;
   wire n4616;
   wire n4617;
   wire n4618;
   wire n4619;
   wire n4620;
   wire n4621;
   wire n4622;
   wire n4623;
   wire n4624;
   wire n4625;
   wire n4626;
   wire n4627;
   wire n4628;
   wire n4629;
   wire n4630;
   wire n4631;
   wire n4632;
   wire n4633;
   wire n4634;
   wire n4635;
   wire n4636;
   wire n4637;
   wire n4638;
   wire n4639;
   wire n4640;
   wire n4641;
   wire n4642;
   wire n4643;
   wire n4644;
   wire n4645;
   wire n4646;
   wire n4647;
   wire n4648;
   wire n4649;
   wire n4650;
   wire n4651;
   wire n4652;
   wire n4653;
   wire n4654;
   wire n4655;
   wire n4656;
   wire n4657;
   wire n4658;
   wire n4659;
   wire n4660;
   wire n4661;
   wire n4662;
   wire n4663;
   wire n4664;
   wire n4665;
   wire n4666;
   wire n4667;
   wire n4668;
   wire n4669;
   wire n4670;
   wire n4671;
   wire n4672;
   wire n4673;
   wire n4674;
   wire n4675;
   wire n4676;
   wire n4677;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n7;
   wire n24;
   wire n25;
   wire n26;
   wire n28;
   wire n29;
   wire n31;
   wire n32;
   wire n34;
   wire n35;
   wire n37;
   wire n38;
   wire n40;
   wire n41;
   wire n43;
   wire n44;
   wire n46;
   wire n47;
   wire n49;
   wire n50;
   wire n52;
   wire n53;
   wire n55;
   wire n56;
   wire n58;
   wire n59;
   wire n61;
   wire n62;
   wire n64;
   wire n65;
   wire n67;
   wire n68;
   wire n70;
   wire n73;
   wire n75;
   wire n76;
   wire n78;
   wire n80;
   wire n82;
   wire n84;
   wire n86;
   wire n88;
   wire n90;
   wire n92;
   wire n94;
   wire n96;
   wire n98;
   wire n100;
   wire n102;
   wire n104;
   wire n107;
   wire n109;
   wire n110;
   wire n112;
   wire n114;
   wire n116;
   wire n118;
   wire n120;
   wire n122;
   wire n124;
   wire n126;
   wire n128;
   wire n130;
   wire n132;
   wire n134;
   wire n136;
   wire n138;
   wire n141;
   wire n143;
   wire n144;
   wire n146;
   wire n148;
   wire n150;
   wire n152;
   wire n154;
   wire n156;
   wire n158;
   wire n160;
   wire n162;
   wire n164;
   wire n166;
   wire n168;
   wire n170;
   wire n172;
   wire n175;
   wire n177;
   wire n178;
   wire n180;
   wire n182;
   wire n184;
   wire n186;
   wire n188;
   wire n190;
   wire n192;
   wire n194;
   wire n196;
   wire n198;
   wire n200;
   wire n202;
   wire n204;
   wire n206;
   wire n209;
   wire n211;
   wire n212;
   wire n214;
   wire n216;
   wire n218;
   wire n220;
   wire n222;
   wire n224;
   wire n226;
   wire n228;
   wire n230;
   wire n232;
   wire n234;
   wire n236;
   wire n238;
   wire n240;
   wire n242;
   wire n244;
   wire n245;
   wire n247;
   wire n249;
   wire n251;
   wire n253;
   wire n255;
   wire n257;
   wire n259;
   wire n261;
   wire n263;
   wire n265;
   wire n267;
   wire n269;
   wire n271;
   wire n273;
   wire n275;
   wire n277;
   wire n278;
   wire n280;
   wire n282;
   wire n284;
   wire n286;
   wire n288;
   wire n290;
   wire n292;
   wire n294;
   wire n296;
   wire n298;
   wire n300;
   wire n302;
   wire n304;
   wire n306;
   wire n308;
   wire n310;
   wire n311;
   wire n313;
   wire n315;
   wire n317;
   wire n319;
   wire n321;
   wire n323;
   wire n325;
   wire n327;
   wire n329;
   wire n331;
   wire n333;
   wire n335;
   wire n337;
   wire n339;
   wire n342;
   wire n344;
   wire n345;
   wire n347;
   wire n349;
   wire n351;
   wire n353;
   wire n355;
   wire n357;
   wire n359;
   wire n361;
   wire n363;
   wire n365;
   wire n367;
   wire n369;
   wire n371;
   wire n373;
   wire n375;
   wire n377;
   wire n378;
   wire n380;
   wire n382;
   wire n384;
   wire n386;
   wire n388;
   wire n390;
   wire n392;
   wire n394;
   wire n396;
   wire n398;
   wire n400;
   wire n402;
   wire n404;
   wire n406;
   wire n408;
   wire n410;
   wire n411;
   wire n413;
   wire n415;
   wire n417;
   wire n419;
   wire n421;
   wire n423;
   wire n425;
   wire n427;
   wire n429;
   wire n431;
   wire n433;
   wire n435;
   wire n437;
   wire n439;
   wire n441;
   wire n443;
   wire n444;
   wire n446;
   wire n448;
   wire n450;
   wire n452;
   wire n454;
   wire n456;
   wire n458;
   wire n460;
   wire n462;
   wire n464;
   wire n466;
   wire n468;
   wire n470;
   wire n472;
   wire n475;
   wire n477;
   wire n478;
   wire n480;
   wire n482;
   wire n484;
   wire n486;
   wire n488;
   wire n490;
   wire n492;
   wire n494;
   wire n496;
   wire n498;
   wire n500;
   wire n502;
   wire n504;
   wire n506;
   wire n508;
   wire n510;
   wire n511;
   wire n513;
   wire n515;
   wire n517;
   wire n519;
   wire n521;
   wire n523;
   wire n525;
   wire n527;
   wire n529;
   wire n531;
   wire n533;
   wire n535;
   wire n537;
   wire n539;
   wire n541;
   wire n543;
   wire n546;
   wire n549;
   wire n552;
   wire n555;
   wire n558;
   wire n560;
   wire n562;
   wire n564;
   wire n567;
   wire n569;
   wire n571;
   wire n573;
   wire n576;
   wire n578;
   wire n580;
   wire n4678;
   wire n4679;
   wire n4680;
   wire n4681;
   wire n4682;
   wire n4683;
   wire n4684;
   wire n4685;
   wire n4686;
   wire n4687;
   wire n4688;
   wire n4689;
   wire n4690;
   wire n4691;
   wire n4692;
   wire n4693;
   wire n4694;
   wire n4695;
   wire n4696;
   wire n4697;
   wire n4698;
   wire n4699;
   wire n4700;
   wire n4701;
   wire n4702;
   wire n4703;
   wire n4704;
   wire n4705;
   wire n4706;
   wire n4707;
   wire n4708;
   wire n4709;
   wire n4710;
   wire n4711;
   wire n4712;
   wire n4713;
   wire n4714;
   wire n4715;
   wire n4716;
   wire n4717;
   wire n4718;
   wire n4719;
   wire n4720;
   wire n4721;
   wire n4722;
   wire n4723;
   wire n4724;
   wire n4725;
   wire n4726;
   wire n4727;
   wire n4728;
   wire n4729;
   wire n4730;
   wire n4731;
   wire n4732;
   wire n4733;
   wire n4734;
   wire n4735;
   wire n4736;
   wire n4737;
   wire n4738;
   wire n4739;
   wire n4740;
   wire n4741;
   wire n4742;
   wire n4743;
   wire n4744;
   wire n4745;
   wire n4746;
   wire n4747;
   wire n4748;
   wire n4749;
   wire n4750;
   wire n4751;
   wire n4752;
   wire n4753;
   wire n4754;
   wire n4755;
   wire n4756;
   wire n4757;
   wire n4758;
   wire n4759;
   wire n4760;
   wire n4761;
   wire n4762;
   wire n4763;
   wire n4764;
   wire n4765;
   wire n4766;
   wire n4767;
   wire n4768;
   wire n4769;
   wire n4770;
   wire n4771;
   wire n4772;
   wire n4773;
   wire n4774;
   wire n4775;
   wire n4776;
   wire n4777;
   wire n4778;
   wire n4779;
   wire n4780;
   wire n4781;
   wire n4782;
   wire n4783;
   wire n4784;
   wire n4785;
   wire n4786;
   wire n4787;
   wire n4788;
   wire n4789;
   wire n4790;
   wire n4791;
   wire n4792;
   wire n4793;
   wire n4794;
   wire n4795;
   wire n4796;
   wire n4797;
   wire n4798;
   wire n4799;
   wire n4800;
   wire n4801;
   wire n4802;
   wire n4803;
   wire n4804;
   wire n4805;
   wire n4806;
   wire n4807;
   wire n4808;
   wire n4809;
   wire n4810;
   wire n4811;
   wire n4812;
   wire n4813;
   wire n4814;
   wire n4815;
   wire n4816;
   wire n4817;
   wire n4818;
   wire n4819;
   wire n4820;
   wire n4821;
   wire n4822;
   wire n4823;
   wire n4824;
   wire n4825;
   wire n4826;
   wire n4827;
   wire n4828;
   wire n4829;
   wire n4830;
   wire n4831;
   wire n4832;
   wire n4833;
   wire n4834;
   wire n4835;
   wire n4836;
   wire n4837;
   wire n4838;
   wire n4839;
   wire n4840;
   wire n4841;
   wire n4842;
   wire n4843;
   wire n4844;
   wire n4845;
   wire n4846;
   wire n4847;
   wire n4848;
   wire n4849;
   wire n4850;
   wire n4851;
   wire n4852;
   wire n4853;
   wire n4854;
   wire n4855;
   wire n4856;
   wire n4857;
   wire n4858;
   wire n4859;
   wire n4860;
   wire n4861;
   wire n4862;
   wire n4863;
   wire n4864;
   wire n4865;
   wire n4866;
   wire n4867;
   wire n4868;
   wire n4869;
   wire n4870;
   wire n4871;
   wire n4872;
   wire n4873;
   wire n4874;
   wire n4875;
   wire n4876;
   wire n4877;
   wire n4878;
   wire n4879;
   wire n4880;
   wire n4881;
   wire n4882;
   wire n4883;
   wire n4884;
   wire n4885;
   wire n4886;
   wire n4887;
   wire n4888;
   wire n4889;
   wire n4890;
   wire n4891;
   wire n4892;
   wire n4893;
   wire n4894;
   wire n4895;
   wire n4896;
   wire n4897;
   wire n4898;
   wire n4899;
   wire n4900;
   wire n4901;
   wire n4902;
   wire n4903;
   wire n4904;
   wire n4905;
   wire n4906;
   wire n4907;
   wire n4908;
   wire n4909;
   wire n4910;
   wire n4911;
   wire n4912;
   wire n4913;
   wire n4914;
   wire n4915;
   wire n4916;
   wire n4917;
   wire n4918;
   wire n4919;
   wire n4920;
   wire n4921;
   wire n4922;
   wire n4923;
   wire n4924;
   wire n4925;
   wire n4926;
   wire n4927;
   wire n4928;
   wire n4929;
   wire n4930;
   wire n4931;
   wire n4932;
   wire n4933;
   wire n4934;
   wire n4935;
   wire n4936;
   wire n4937;
   wire n4938;
   wire n4939;
   wire n4940;
   wire n4941;
   wire n4942;
   wire n4943;
   wire n4944;
   wire n4945;
   wire n4946;
   wire n4947;
   wire n4948;
   wire n4949;
   wire n4950;
   wire n4951;
   wire n4952;
   wire n4953;
   wire n4954;
   wire n4955;
   wire n4956;
   wire n4957;
   wire n4958;
   wire n4959;
   wire n4960;
   wire n4961;
   wire n4962;
   wire n4963;
   wire n4964;
   wire n4965;
   wire n4966;
   wire n4967;
   wire n4968;
   wire n4969;
   wire n4970;
   wire n4971;
   wire n4972;
   wire n4973;
   wire n4974;
   wire n4975;
   wire n4976;
   wire n4977;
   wire n4978;
   wire n4979;
   wire n4980;
   wire n4981;
   wire n4982;
   wire n4983;
   wire n4984;
   wire n4985;
   wire n4986;
   wire n4987;
   wire n4988;
   wire n4989;
   wire n4990;
   wire n4991;
   wire n4992;
   wire n4993;
   wire n4994;
   wire n4995;
   wire n4996;
   wire n4997;
   wire n4998;
   wire n4999;
   wire n5000;
   wire n5001;
   wire n5002;
   wire n5003;
   wire n5004;
   wire n5005;
   wire n5006;
   wire n5007;
   wire n5008;
   wire n5009;
   wire n5010;
   wire n5011;
   wire n5012;
   wire n5013;
   wire n5014;
   wire n5015;
   wire n5016;
   wire n5017;
   wire n5018;
   wire n5019;
   wire n5020;
   wire n5021;
   wire n5022;
   wire n5023;
   wire n5024;
   wire n5025;
   wire n5026;
   wire n5027;
   wire n5028;
   wire n5029;
   wire n5030;
   wire n5031;
   wire n5032;
   wire n5033;
   wire n5034;
   wire n5035;
   wire n5036;
   wire n5037;
   wire n5038;
   wire n5039;
   wire n5040;
   wire n5041;
   wire n5042;
   wire n5043;
   wire n5044;
   wire n5045;
   wire n5046;
   wire n5047;
   wire n5048;
   wire n5049;
   wire n5050;
   wire n5051;
   wire n5052;
   wire n5053;
   wire n5054;
   wire n5055;
   wire n5056;
   wire n5057;
   wire n5058;
   wire n5059;
   wire n5060;
   wire n5061;
   wire n5062;
   wire n5063;
   wire n5064;
   wire n5065;
   wire n5066;
   wire n5067;
   wire n5068;
   wire n5069;
   wire n5070;
   wire n5071;
   wire n5072;
   wire n5073;
   wire n5074;
   wire n5075;
   wire n5076;
   wire n5077;
   wire n5078;
   wire n5079;
   wire n5080;
   wire n5081;
   wire n5082;
   wire n5083;
   wire n5084;
   wire n5085;
   wire n5086;
   wire n5087;
   wire n5088;
   wire n5089;
   wire n5090;
   wire n5091;
   wire n5092;
   wire n5093;
   wire n5094;
   wire n5095;
   wire n5096;
   wire n5097;
   wire n5098;
   wire n5099;
   wire n5100;
   wire n5101;
   wire n5102;
   wire n5103;
   wire n5104;
   wire n5105;
   wire n5106;
   wire n5107;
   wire n5108;
   wire n5109;
   wire n5110;
   wire n5111;
   wire n5112;
   wire n5113;
   wire n5114;
   wire n5115;
   wire n5116;
   wire n5117;
   wire n5118;
   wire n5119;
   wire n5120;
   wire n5121;
   wire n5122;
   wire n5123;
   wire n5124;
   wire n5125;
   wire n5126;
   wire n5127;
   wire n5128;
   wire n5129;
   wire n5130;
   wire n5131;
   wire n5132;
   wire n5133;
   wire n5134;
   wire n5135;
   wire n5136;
   wire n5137;
   wire n5138;
   wire n5139;
   wire n5140;
   wire n5141;
   wire n5142;
   wire n5143;
   wire n5144;
   wire n5145;
   wire n5146;
   wire n5147;
   wire n5148;
   wire n5149;
   wire n5150;
   wire n5151;
   wire n5152;
   wire n5153;
   wire n5154;
   wire n5155;
   wire n5156;
   wire n5157;
   wire n5158;
   wire n5159;
   wire n5160;
   wire n5161;
   wire n5162;
   wire n5163;
   wire n5164;
   wire n5165;
   wire n5166;
   wire n5167;
   wire n5168;
   wire n5169;
   wire n5170;
   wire n5171;
   wire n5172;
   wire n5173;
   wire n5174;
   wire n5175;
   wire n5176;
   wire n5177;
   wire n5178;
   wire n5179;
   wire n5180;
   wire n5181;
   wire n5182;
   wire n5183;
   wire n5184;
   wire n5185;
   wire n5186;
   wire n5187;
   wire n5188;
   wire n5189;
   wire n5190;
   wire n5191;
   wire n5192;
   wire n5193;
   wire n5194;
   wire n5195;
   wire n5196;
   wire n5197;
   wire n5198;
   wire n5199;
   wire n5200;
   wire n5201;
   wire n5202;
   wire n5203;
   wire n5204;
   wire n5205;
   wire n5206;
   wire n5207;
   wire n5208;
   wire n5209;
   wire n5210;
   wire n5211;
   wire n5212;
   wire n5213;
   wire n5214;
   wire n5215;
   wire n5216;
   wire n5217;
   wire n5218;
   wire n5219;
   wire n5220;
   wire n5221;
   wire n5222;
   wire n5223;
   wire n5224;
   wire n5225;
   wire n5226;
   wire n5227;
   wire n5228;
   wire n5229;
   wire n5230;
   wire n5231;
   wire n5232;
   wire n5233;
   wire n5234;
   wire n5235;
   wire n5236;
   wire n5237;
   wire n5238;
   wire n5239;
   wire n5240;
   wire n5241;
   wire n5242;
   wire n5243;
   wire n5244;
   wire n5245;
   wire n5246;
   wire n5247;
   wire n5248;
   wire n5249;
   wire n5250;
   wire n5251;
   wire n5252;
   wire n5253;
   wire n5254;
   wire n5255;
   wire n5256;
   wire n5257;
   wire n5258;
   wire n5259;
   wire n5260;
   wire n5261;
   wire n5262;
   wire n5263;
   wire n5264;
   wire n5265;
   wire n5266;
   wire n5267;
   wire n5268;
   wire n5269;
   wire n5270;
   wire n5271;
   wire n5272;
   wire n5273;
   wire n5274;
   wire n5275;
   wire n5276;
   wire n5277;
   wire n5278;
   wire n5279;
   wire n5280;
   wire n5281;
   wire n5282;
   wire n5283;
   wire n5284;
   wire n5285;
   wire n5286;
   wire n5287;
   wire n5288;
   wire n5289;
   wire n5290;
   wire n5291;
   wire n5292;
   wire n5293;
   wire n5294;
   wire n5295;
   wire n5296;
   wire n5297;
   wire n5298;
   wire n5299;
   wire n5300;
   wire n5301;
   wire n5302;
   wire n5303;
   wire n5304;
   wire n5305;
   wire n5306;
   wire n5307;
   wire n5308;
   wire n5309;
   wire n5310;
   wire n5311;
   wire n5312;
   wire n5313;
   wire n5314;
   wire n5315;
   wire n5316;
   wire n5317;
   wire n5318;
   wire n5319;
   wire n5320;
   wire n5321;
   wire n5322;
   wire n5323;
   wire n5324;
   wire n5325;
   wire n5326;
   wire n5327;
   wire n5328;
   wire n5329;
   wire n5330;
   wire n5331;
   wire n5332;
   wire n5333;
   wire n5334;
   wire n5335;
   wire n5336;
   wire n5337;
   wire n5338;
   wire n5339;
   wire n5340;
   wire n5341;
   wire n5342;
   wire n5343;
   wire n5344;
   wire n5345;
   wire n5346;
   wire n5347;
   wire n5348;
   wire n5349;
   wire n5350;
   wire n5351;
   wire n5352;
   wire n5353;
   wire n5354;
   wire n5355;
   wire n5356;
   wire n5357;
   wire n5358;
   wire n5359;
   wire n5360;
   wire n5361;
   wire n5362;
   wire n5363;
   wire n5364;
   wire n5365;
   wire n5366;
   wire n5367;
   wire n5368;
   wire n5369;
   wire n5370;
   wire n5371;
   wire n5372;
   wire n5373;
   wire n5374;
   wire n5375;
   wire n5376;
   wire n5377;
   wire n5378;
   wire n5379;
   wire n5380;
   wire n5381;
   wire n5382;
   wire n5383;
   wire n5384;
   wire n5385;
   wire n5386;
   wire n5387;
   wire n5388;
   wire n5389;
   wire n5390;
   wire n5391;
   wire n5392;
   wire n5393;
   wire n5394;
   wire n5395;
   wire n5396;
   wire n5397;
   wire n5398;
   wire n5399;
   wire n5400;
   wire n5401;
   wire n5402;
   wire n5403;
   wire n5404;
   wire n5405;
   wire n5406;
   wire n5407;
   wire n5408;
   wire n5409;
   wire n5410;
   wire n5411;
   wire n5412;
   wire n5413;
   wire n5414;
   wire n5415;
   wire n5416;
   wire n5417;
   wire n5418;
   wire n5419;
   wire n5420;
   wire n5421;
   wire n5422;
   wire n5423;
   wire n5424;
   wire n5425;
   wire n5426;
   wire n5427;
   wire n5428;
   wire n5429;
   wire n5430;
   wire n5431;
   wire n5432;
   wire n5433;
   wire n5434;
   wire n5435;
   wire n5436;
   wire n5437;
   wire n5438;
   wire n5439;
   wire n5440;
   wire n5441;
   wire n5442;
   wire n5443;
   wire n5444;
   wire n5445;
   wire n5446;
   wire n5447;
   wire n5448;
   wire n5449;
   wire n5450;
   wire n5451;
   wire n5452;
   wire n5453;
   wire n5454;
   wire n5455;
   wire n5456;
   wire n5457;
   wire n5458;
   wire n5459;
   wire n5460;
   wire n5461;
   wire n5462;
   wire n5463;
   wire n5464;
   wire n5465;
   wire n5466;
   wire n5467;
   wire n5468;
   wire n5469;
   wire n5470;
   wire n5471;
   wire n5472;
   wire n5473;
   wire n5474;
   wire n5475;
   wire n5476;
   wire n5477;
   wire n5478;
   wire n5479;
   wire n5480;
   wire n5481;
   wire n5482;
   wire n5483;
   wire n5484;
   wire n5485;
   wire n5486;
   wire n5487;
   wire n5488;
   wire n5489;
   wire n5490;
   wire n5491;
   wire n5492;
   wire n5493;
   wire n5494;
   wire n5495;
   wire n5496;
   wire n5497;
   wire n5498;
   wire n5499;
   wire n5500;
   wire n5501;
   wire n5502;
   wire n5503;
   wire n5504;
   wire n5505;
   wire n5506;
   wire n5507;
   wire n5508;
   wire n5509;
   wire n5510;
   wire n5511;
   wire n5512;
   wire n5513;
   wire n5514;
   wire n5515;
   wire n5516;
   wire n5517;
   wire n5518;
   wire n5519;
   wire n5520;
   wire n5521;
   wire n5522;
   wire n5523;
   wire n5524;
   wire n5525;
   wire n5526;
   wire n5527;
   wire n5528;
   wire n5529;
   wire n5530;
   wire n5531;
   wire n5532;
   wire n5533;
   wire n5534;
   wire n5535;
   wire n5536;
   wire n5537;
   wire n5538;
   wire n5539;
   wire n5540;
   wire n5541;
   wire n5542;
   wire n5543;
   wire n5544;
   wire n5545;
   wire n5546;
   wire n5547;
   wire n5548;
   wire n5549;
   wire n5550;
   wire n5551;
   wire n5552;
   wire n5553;
   wire n5554;
   wire n5555;
   wire n5556;
   wire n5557;
   wire n5558;
   wire n5559;
   wire n5560;
   wire n5561;
   wire n5562;
   wire n5563;
   wire n5564;
   wire n5565;
   wire n5566;
   wire n5567;
   wire n5568;
   wire n5569;
   wire n5570;
   wire n5571;
   wire n5572;
   wire n5573;
   wire n5574;
   wire n5575;
   wire n5576;
   wire n5577;
   wire n5578;
   wire n5579;
   wire n5580;
   wire n5581;
   wire n5582;
   wire n5583;
   wire n5584;
   wire n5585;
   wire n5586;
   wire n5587;
   wire n5588;
   wire n5589;
   wire n5590;
   wire n5591;
   wire n5592;
   wire n5593;
   wire n5594;
   wire n5595;
   wire n5596;
   wire n5597;
   wire n5598;
   wire n5599;
   wire n5600;
   wire n5601;
   wire n5602;
   wire n5603;
   wire n5604;
   wire n5605;
   wire n5606;
   wire n5607;
   wire n5608;
   wire n5609;
   wire n5610;
   wire n5611;
   wire n5612;
   wire n5613;
   wire n5614;
   wire n5615;
   wire n5616;
   wire n5617;
   wire n5618;
   wire n5619;
   wire n5620;
   wire n5621;
   wire n5622;
   wire n5623;
   wire n5624;
   wire n5625;
   wire n5626;
   wire n5627;
   wire n5628;
   wire n5629;
   wire n5630;
   wire n5631;
   wire n5632;
   wire n5633;
   wire n5634;
   wire n5635;
   wire n5636;
   wire n5637;
   wire n5638;
   wire n5639;
   wire n5640;
   wire n5641;
   wire n5642;
   wire n5643;
   wire n5644;
   wire n5645;
   wire n5646;
   wire n5647;
   wire n5648;
   wire n5649;
   wire n5650;
   wire n5651;
   wire n5652;
   wire n5653;
   wire n5654;
   wire n5655;
   wire n5656;
   wire n5657;
   wire n5658;
   wire n5659;
   wire n5660;
   wire n5661;
   wire n5662;
   wire n5663;
   wire n5664;
   wire n5665;
   wire n5666;
   wire n5667;
   wire n5668;
   wire n5669;
   wire n5670;
   wire n5671;
   wire n5672;
   wire n5673;
   wire n5674;
   wire n5675;
   wire n5676;
   wire n5677;
   wire n5678;
   wire n5679;
   wire n5680;
   wire n5681;
   wire n5682;
   wire n5683;
   wire n5684;
   wire n5685;
   wire n5686;
   wire n5687;
   wire n5688;
   wire n5689;
   wire n5690;
   wire n5691;
   wire n5692;
   wire n5693;
   wire n5694;
   wire n5695;
   wire n5696;
   wire n5697;
   wire n5698;
   wire n5699;
   wire n5700;
   wire n5701;
   wire n5702;
   wire n5703;
   wire n5704;
   wire n5705;
   wire n5706;
   wire n5707;
   wire n5708;
   wire n5709;
   wire n5710;
   wire n5711;
   wire n5712;
   wire n5713;
   wire n5714;
   wire n5715;
   wire n5716;
   wire n5717;
   wire n5718;
   wire n5719;
   wire n5720;
   wire n5721;
   wire n5722;
   wire n5723;
   wire n5724;
   wire n5725;
   wire n5726;
   wire n5727;
   wire n5728;
   wire n5729;
   wire n5730;
   wire n5731;
   wire n5732;
   wire n5733;
   wire n5734;
   wire n5735;
   wire n5736;
   wire n5737;
   wire n5738;
   wire n5739;
   wire n5740;
   wire n5741;
   wire n5742;
   wire n5743;
   wire n5744;
   wire n5745;
   wire n5746;
   wire n5747;
   wire n5748;
   wire n5749;
   wire n5750;
   wire n5751;
   wire n5752;
   wire n5753;
   wire n5754;
   wire n5755;
   wire n5756;
   wire n5757;
   wire n5758;
   wire n5759;
   wire n5760;
   wire n5761;
   wire n5762;
   wire n5763;
   wire n5764;
   wire n5765;
   wire n5766;
   wire n5767;
   wire n5768;
   wire n5769;
   wire n5770;
   wire n5771;
   wire n5772;
   wire n5773;
   wire n5774;
   wire n5775;
   wire n5776;
   wire n5777;
   wire n5778;
   wire n5779;
   wire n5780;
   wire n5781;
   wire n5782;
   wire n5783;
   wire n5784;
   wire n5785;
   wire n5786;
   wire n5787;
   wire n5788;
   wire n5789;
   wire n5790;
   wire n5791;
   wire n5792;
   wire n5793;
   wire n5794;
   wire n5795;
   wire n5796;
   wire n5797;
   wire n5798;
   wire n5799;
   wire n5800;
   wire n5801;
   wire n5802;
   wire n5803;
   wire n5804;
   wire n5805;
   wire n5806;
   wire n5807;
   wire n5808;
   wire n5809;
   wire n5810;
   wire n5811;
   wire n5812;
   wire n5813;
   wire n5814;
   wire n5815;
   wire n5816;
   wire n5817;
   wire n5818;
   wire n5819;
   wire n5820;
   wire n5821;
   wire n5822;
   wire n5823;
   wire n5824;
   wire n5825;
   wire n5826;
   wire n5827;
   wire n5828;
   wire n5829;
   wire n5830;
   wire n5831;
   wire n5832;
   wire n5833;
   wire n5834;
   wire n5835;
   wire n5836;
   wire n5837;
   wire n5838;
   wire n5839;
   wire n5840;
   wire n5841;
   wire n5842;
   wire n5843;
   wire n5844;
   wire n5845;
   wire n5846;
   wire n5847;
   wire n5848;
   wire n5849;
   wire n5850;
   wire n5851;
   wire n5852;
   wire n5853;
   wire n5854;
   wire n5855;
   wire n5856;
   wire n5857;
   wire n5858;
   wire n5859;
   wire n5860;
   wire n5861;
   wire n5862;
   wire n5863;
   wire n5864;
   wire n5865;
   wire n5866;
   wire n5867;
   wire n5868;
   wire n5869;
   wire n5870;
   wire n5871;
   wire n5872;
   wire n5873;
   wire n5874;
   wire n5875;
   wire n5876;
   wire n5877;
   wire n5878;
   wire n5879;
   wire n5880;
   wire n5881;
   wire n5882;
   wire n5883;
   wire n5884;
   wire n5885;
   wire n5886;
   wire n5887;
   wire n5888;
   wire n5889;
   wire n5890;
   wire n5891;
   wire n5892;
   wire n5893;
   wire n5894;
   wire n5895;
   wire n5896;
   wire n5897;
   wire n5898;
   wire n5899;
   wire n5900;
   wire n5901;
   wire n5902;
   wire n5903;
   wire n5904;
   wire n5905;
   wire n5906;
   wire n5907;
   wire n5908;
   wire n5909;
   wire n5910;
   wire n5911;
   wire n5912;
   wire n5913;
   wire n5914;
   wire n5915;
   wire n5916;
   wire n5917;
   wire n5918;
   wire n5919;
   wire n5920;
   wire n5921;
   wire n5922;
   wire n5923;
   wire n5924;
   wire n5925;
   wire n5926;
   wire n5927;
   wire n5928;
   wire n5929;
   wire n5930;
   wire n5931;
   wire n5932;
   wire n5933;
   wire n5934;
   wire n5935;
   wire n5936;
   wire n5937;
   wire n5938;
   wire n5939;
   wire n5940;
   wire n5941;
   wire n5942;
   wire n5943;
   wire n5944;
   wire n5945;
   wire n5946;
   wire n5947;
   wire n5948;
   wire n5949;
   wire n5950;
   wire n5951;
   wire n5952;
   wire n5953;
   wire n5954;
   wire n5955;
   wire n5956;
   wire n5957;
   wire n5958;
   wire n5959;
   wire n5960;
   wire n5961;
   wire n5962;
   wire n5963;
   wire n5964;
   wire n5965;
   wire n5966;
   wire n5967;
   wire n5968;
   wire n5969;
   wire n5970;
   wire n5971;
   wire n5972;
   wire n5973;
   wire n5974;
   wire n5975;
   wire n5976;
   wire n5977;
   wire n5978;
   wire n5979;
   wire n5980;
   wire n5981;
   wire n5982;
   wire n5983;
   wire n5984;
   wire n5985;
   wire n5986;
   wire n5987;
   wire n5988;
   wire n5989;
   wire n5990;
   wire n5991;
   wire n5992;
   wire n5993;
   wire n5994;
   wire n5995;
   wire n5996;
   wire n5997;
   wire n5998;
   wire n5999;
   wire n6000;
   wire n6001;
   wire n6002;
   wire n6003;
   wire n6004;
   wire n6005;
   wire n6006;
   wire n6007;
   wire n6008;
   wire n6009;
   wire n6010;
   wire n6011;
   wire n6012;
   wire n6013;
   wire n6014;
   wire n6015;
   wire n6016;
   wire n6038;
   wire n6136;
   wire n6459;
   wire n6469;
   wire n6470;
   wire n6471;
   wire n7439;
   wire n7440;
   wire n7441;
   wire n7442;
   wire n7443;
   wire n7444;
   wire n7445;

   assign N20 = mem_access_addr[2] ;
   assign N21 = mem_access_addr[3] ;
   assign N22 = mem_access_addr[4] ;
   assign N23 = mem_access_addr[5] ;
   assign N24 = mem_access_addr[6] ;
   assign N25 = mem_access_addr[7] ;
   assign N26 = mem_access_addr[8] ;
   assign N27 = mem_access_addr[9] ;

   BUFCKEHD FE_PHC7506_n2582 (.O(FE_PHN7506_n2582), 
	.I(n2582));
   BUFCHD FE_PHC7505_n2417 (.O(FE_PHN7505_n2417), 
	.I(n2417));
   BUFCKEHD FE_PHC7504_n2582 (.O(FE_PHN7504_n2582), 
	.I(FE_PHN7506_n2582));
   BUFCHD FE_PHC7503_n1001 (.O(FE_PHN7503_n1001), 
	.I(FE_PHN7457_n1001));
   BUFCHD FE_PHC7502_n1014 (.O(FE_PHN7502_n1014), 
	.I(FE_PHN7490_n1014));
   BUFCHD FE_PHC7501_n2890 (.O(FE_PHN7501_n2890), 
	.I(n2890));
   BUFCKEHD FE_PHC7500_n2180 (.O(FE_PHN7500_n2180), 
	.I(FE_PHN7230_n2180));
   BUFCKEHD FE_PHC7499_n4102 (.O(FE_PHN7499_n4102), 
	.I(FE_PHN4942_n4102));
   BUFCKEHD FE_PHC7498_n2395 (.O(FE_PHN7498_n2395), 
	.I(FE_PHN4778_n2395));
   BUFCHD FE_PHC7497_n2417 (.O(FE_PHN7497_n2417), 
	.I(FE_PHN7505_n2417));
   BUFCHD FE_PHC7496_n2582 (.O(FE_PHN7496_n2582), 
	.I(FE_PHN7504_n2582));
   BUFCKEHD FE_PHC7495_n1013 (.O(n1013), 
	.I(FE_PHN7495_n1013));
   BUFCHD FE_PHC7494_n1001 (.O(FE_PHN7494_n1001), 
	.I(FE_PHN7503_n1001));
   BUFCKEHD FE_PHC7493_n3964 (.O(FE_PHN7493_n3964), 
	.I(n3964));
   BUFCKEHD FE_PHC7492_n1017 (.O(FE_PHN7492_n1017), 
	.I(n1017));
   BUFCHD FE_PHC7491_n974 (.O(FE_PHN7491_n974), 
	.I(n974));
   BUFCKEHD FE_PHC7490_n1014 (.O(FE_PHN7490_n1014), 
	.I(n1014));
   BUFCKEHD FE_PHC7489_n2394 (.O(FE_PHN7489_n2394), 
	.I(FE_PHN4792_n2394));
   BUFCKEHD FE_PHC7488_n3953 (.O(FE_PHN7488_n3953), 
	.I(FE_PHN3941_n3953));
   BUFCKEHD FE_PHC7487_n3934 (.O(FE_PHN7487_n3934), 
	.I(n3934));
   BUFDHD FE_PHC7486_n2132 (.O(FE_PHN7486_n2132), 
	.I(FE_PHN4845_n2132));
   BUFCHD FE_PHC7485_n2168 (.O(FE_PHN7485_n2168), 
	.I(FE_PHN4775_n2168));
   BUFCKEHD FE_PHC7484_n3960 (.O(FE_PHN7484_n3960), 
	.I(FE_PHN3944_n3960));
   BUFCKEHD FE_PHC7483_n2571 (.O(FE_PHN7483_n2571), 
	.I(FE_PHN4819_n2571));
   BUFCKEHD FE_PHC7482_n3923 (.O(FE_PHN7482_n3923), 
	.I(FE_PHN3501_n3923));
   BUFCKEHD FE_PHC7481_n2892 (.O(FE_PHN7481_n2892), 
	.I(FE_PHN4868_n2892));
   BUFCKEHD FE_PHC7480_n2155 (.O(FE_PHN7480_n2155), 
	.I(FE_PHN6691_n2155));
   BUFCHD FE_PHC7479_n2175 (.O(FE_PHN7479_n2175), 
	.I(FE_PHN4921_n2175));
   BUFCKEHD FE_PHC7478_n3968 (.O(FE_PHN7478_n3968), 
	.I(FE_PHN3798_n3968));
   BUFCHD FE_PHC7477_n2628 (.O(FE_PHN7477_n2628), 
	.I(FE_PHN4859_n2628));
   BUFCKEHD FE_PHC7476_n2159 (.O(FE_PHN7476_n2159), 
	.I(FE_PHN4886_n2159));
   BUFCHD FE_PHC7475_n2592 (.O(FE_PHN7475_n2592), 
	.I(FE_PHN6688_n2592));
   BUFCKEHD FE_PHC7474_n4155 (.O(FE_PHN7474_n4155), 
	.I(FE_PHN4846_n4155));
   BUFCHD FE_PHC7473_n2170 (.O(FE_PHN7473_n2170), 
	.I(FE_PHN4809_n2170));
   BUFCHD FE_PHC7472_n4137 (.O(FE_PHN7472_n4137), 
	.I(FE_PHN7409_n4137));
   BUFCHD FE_PHC7471_n4147 (.O(FE_PHN7471_n4147), 
	.I(FE_PHN4903_n4147));
   BUFCHD FE_PHC7470_n2166 (.O(FE_PHN7470_n2166), 
	.I(FE_PHN4860_n2166));
   BUFCHD FE_PHC7469_n3230 (.O(FE_PHN7469_n3230), 
	.I(FE_PHN4873_n3230));
   BUFCHD FE_PHC7468_n2614 (.O(FE_PHN7468_n2614), 
	.I(FE_PHN4889_n2614));
   BUFCKEHD FE_PHC7467_n2395 (.O(FE_PHN7467_n2395), 
	.I(FE_PHN7498_n2395));
   BUFCHD FE_PHC7466_n2130 (.O(FE_PHN7466_n2130), 
	.I(FE_PHN6658_n2130));
   BUFCHD FE_PHC7465_n2890 (.O(FE_PHN7465_n2890), 
	.I(FE_PHN7501_n2890));
   BUFCHD FE_PHC7464_n4102 (.O(FE_PHN7464_n4102), 
	.I(FE_PHN7499_n4102));
   BUFCHD FE_PHC7463_n2180 (.O(FE_PHN7463_n2180), 
	.I(FE_PHN7500_n2180));
   BUFCKEHD FE_PHC7462_n2417 (.O(n2417), 
	.I(FE_PHN7462_n2417));
   BUFCKEHD FE_PHC7461_n2582 (.O(n2582), 
	.I(FE_PHN7461_n2582));
   BUFCKEHD FE_PHC7460_n979 (.O(FE_PHN7460_n979), 
	.I(FE_PHN4898_n979));
   BUFCKEHD FE_PHC7459_n1154 (.O(FE_PHN7459_n1154), 
	.I(FE_PHN4863_n1154));
   BUFCKEHD FE_PHC7458_n938 (.O(FE_PHN7458_n938), 
	.I(n938));
   BUFIHD FE_PHC7457_n1001 (.O(FE_PHN7457_n1001), 
	.I(n1001));
   BUFCKEHD FE_PHC7456_n4215 (.O(n4215), 
	.I(FE_PHN7456_n4215));
   BUFCHD FE_PHC7455_n3129 (.O(FE_PHN7455_n3129), 
	.I(n3129));
   BUFCKEHD FE_PHC7454_n4229 (.O(n4229), 
	.I(FE_PHN7454_n4229));
   BUFCKEHD FE_PHC7453_n3964 (.O(n3964), 
	.I(FE_PHN7453_n3964));
   BUFCKEHD FE_PHC7452_n3028 (.O(FE_PHN7452_n3028), 
	.I(n3028));
   BUFCKEHD FE_PHC7451_n974 (.O(n974), 
	.I(FE_PHN7451_n974));
   BUFCHD FE_PHC7450_n1017 (.O(FE_PHN7450_n1017), 
	.I(FE_PHN7492_n1017));
   BUFCKEHD FE_PHC7449_n1014 (.O(n1014), 
	.I(FE_PHN7449_n1014));
   BUFCHD FE_PHC7448_n2426 (.O(FE_PHN7448_n2426), 
	.I(FE_PHN4839_n2426));
   BUFCKEHD FE_PHC7447_n4013 (.O(FE_PHN7447_n4013), 
	.I(n4013));
   BUFCKEHD FE_PHC7446_n2119 (.O(FE_PHN7446_n2119), 
	.I(FE_PHN4909_n2119));
   BUFCHD FE_PHC7445_n2393 (.O(FE_PHN7445_n2393), 
	.I(FE_PHN4802_n2393));
   BUFCHD FE_PHC7444_n2133 (.O(FE_PHN7444_n2133), 
	.I(FE_PHN4938_n2133));
   BUFCHD FE_PHC7443_n2604 (.O(FE_PHN7443_n2604), 
	.I(FE_PHN6683_n2604));
   BUFCKEHD FE_PHC7442_n3068 (.O(FE_PHN7442_n3068), 
	.I(n3068));
   BUFCHD FE_PHC7441_n2164 (.O(FE_PHN7441_n2164), 
	.I(FE_PHN4789_n2164));
   BUFCKEHD FE_PHC7440_n2126 (.O(FE_PHN7440_n2126), 
	.I(FE_PHN4950_n2126));
   BUFCHD FE_PHC7439_n2378 (.O(FE_PHN7439_n2378), 
	.I(FE_PHN4908_n2378));
   BUFCKEHD FE_PHC7438_n2151 (.O(FE_PHN7438_n2151), 
	.I(FE_PHN4791_n2151));
   BUFCHD FE_PHC7437_n2610 (.O(FE_PHN7437_n2610), 
	.I(FE_PHN6710_n2610));
   BUFCKEHD FE_PHC7436_n2165 (.O(FE_PHN7436_n2165), 
	.I(FE_PHN4840_n2165));
   BUFCKEHD FE_PHC7435_n2379 (.O(FE_PHN7435_n2379), 
	.I(FE_PHN4850_n2379));
   BUFCHD FE_PHC7434_n2118 (.O(FE_PHN7434_n2118), 
	.I(FE_PHN6656_n2118));
   BUFCHD FE_PHC7433_n2167 (.O(FE_PHN7433_n2167), 
	.I(FE_PHN4795_n2167));
   BUFCHD FE_PHC7432_n2603 (.O(FE_PHN7432_n2603), 
	.I(FE_PHN6677_n2603));
   BUFCKEHD FE_PHC7431_n2135 (.O(FE_PHN7431_n2135), 
	.I(FE_PHN4816_n2135));
   BUFCHD FE_PHC7430_n2887 (.O(FE_PHN7430_n2887), 
	.I(FE_PHN7280_n2887));
   BUFCHD FE_PHC7429_n2169 (.O(FE_PHN7429_n2169), 
	.I(FE_PHN4874_n2169));
   BUFCKEHD FE_PHC7428_n3953 (.O(FE_PHN7428_n3953), 
	.I(FE_PHN7488_n3953));
   BUFCHD FE_PHC7427_n2179 (.O(FE_PHN7427_n2179), 
	.I(n2179));
   BUFCKEHD FE_PHC7426_n3934 (.O(FE_PHN7426_n3934), 
	.I(FE_PHN7487_n3934));
   BUFCHD FE_PHC7425_n2154 (.O(FE_PHN7425_n2154), 
	.I(FE_PHN4955_n2154));
   BUFCHD FE_PHC7424_n2168 (.O(FE_PHN7424_n2168), 
	.I(FE_PHN7485_n2168));
   BUFCHD FE_PHC7423_n2892 (.O(FE_PHN7423_n2892), 
	.I(FE_PHN7481_n2892));
   BUFCKEHD FE_PHC7422_n2570 (.O(FE_PHN7422_n2570), 
	.I(FE_PHN4880_n2570));
   BUFCHD FE_PHC7421_n2434 (.O(FE_PHN7421_n2434), 
	.I(FE_PHN4895_n2434));
   BUFEHD FE_PHC7420_n3968 (.O(FE_PHN7420_n3968), 
	.I(FE_PHN7478_n3968));
   BUFCKEHD FE_PHC7419_n4155 (.O(FE_PHN7419_n4155), 
	.I(FE_PHN7474_n4155));
   BUFCHD FE_PHC7418_n2410 (.O(FE_PHN7418_n2410), 
	.I(FE_PHN6645_n2410));
   BUFCKEHD FE_PHC7417_n2152 (.O(FE_PHN7417_n2152), 
	.I(FE_PHN4824_n2152));
   BUFCHD FE_PHC7416_n2132 (.O(FE_PHN7416_n2132), 
	.I(FE_PHN7486_n2132));
   BUFCKEHD FE_PHC7415_n2175 (.O(FE_PHN7415_n2175), 
	.I(FE_PHN7479_n2175));
   BUFCHD FE_PHC7414_n2394 (.O(FE_PHN7414_n2394), 
	.I(FE_PHN7489_n2394));
   BUFCHD FE_PHC7413_n2170 (.O(FE_PHN7413_n2170), 
	.I(FE_PHN7473_n2170));
   BUFCKEHD FE_PHC7412_n2120 (.O(FE_PHN7412_n2120), 
	.I(FE_PHN4851_n2120));
   BUFEHD FE_PHC7411_n2628 (.O(FE_PHN7411_n2628), 
	.I(FE_PHN7477_n2628));
   BUFCHD FE_PHC7410_n4121 (.O(FE_PHN7410_n4121), 
	.I(FE_PHN4777_n4121));
   BUFHHD FE_PHC7409_n4137 (.O(FE_PHN7409_n4137), 
	.I(n4137));
   BUFCHD FE_PHC7408_n2402 (.O(FE_PHN7408_n2402), 
	.I(FE_PHN4853_n2402));
   BUFCHD FE_PHC7407_n2571 (.O(FE_PHN7407_n2571), 
	.I(FE_PHN7483_n2571));
   BUFCHD FE_PHC7406_n3960 (.O(FE_PHN7406_n3960), 
	.I(FE_PHN7484_n3960));
   BUFCHD FE_PHC7405_n2155 (.O(FE_PHN7405_n2155), 
	.I(FE_PHN7480_n2155));
   BUFCHD FE_PHC7404_n3923 (.O(FE_PHN7404_n3923), 
	.I(FE_PHN7482_n3923));
   BUFCHD FE_PHC7403_n2625 (.O(FE_PHN7403_n2625), 
	.I(FE_PHN4927_n2625));
   BUFCHD FE_PHC7402_n2578 (.O(FE_PHN7402_n2578), 
	.I(FE_PHN4843_n2578));
   BUFCKEHD FE_PHC7401_n1863 (.O(FE_PHN7401_n1863), 
	.I(FE_PHN4919_n1863));
   BUFDHD FE_PHC7400_n2159 (.O(FE_PHN7400_n2159), 
	.I(FE_PHN7476_n2159));
   BUFCHD FE_PHC7399_n4139 (.O(FE_PHN7399_n4139), 
	.I(FE_PHN7223_n4139));
   BUFCHD FE_PHC7398_n2166 (.O(FE_PHN7398_n2166), 
	.I(FE_PHN7470_n2166));
   BUFCKEHD FE_PHC7397_n2395 (.O(FE_PHN7397_n2395), 
	.I(FE_PHN7467_n2395));
   BUFEHD FE_PHC7396_n2592 (.O(FE_PHN7396_n2592), 
	.I(FE_PHN7475_n2592));
   BUFCHD FE_PHC7395_n3230 (.O(FE_PHN7395_n3230), 
	.I(FE_PHN7469_n3230));
   BUFCHD FE_PHC7394_n4163 (.O(FE_PHN7394_n4163), 
	.I(FE_PHN4782_n4163));
   BUFCHD FE_PHC7393_n2614 (.O(FE_PHN7393_n2614), 
	.I(FE_PHN7468_n2614));
   BUFCHD FE_PHC7392_n4147 (.O(FE_PHN7392_n4147), 
	.I(FE_PHN7471_n4147));
   BUFCHD FE_PHC7391_n2130 (.O(FE_PHN7391_n2130), 
	.I(FE_PHN7466_n2130));
   BUFCHD FE_PHC7390_n2890 (.O(FE_PHN7390_n2890), 
	.I(FE_PHN7465_n2890));
   BUFCHD FE_PHC7389_n4102 (.O(FE_PHN7389_n4102), 
	.I(FE_PHN7464_n4102));
   BUFCHD FE_PHC7388_n2180 (.O(FE_PHN7388_n2180), 
	.I(FE_PHN7463_n2180));
   BUFCKGHD FE_PHC7387_n2417 (.O(FE_PHN7387_n2417), 
	.I(FE_PHN7497_n2417));
   BUFCHD FE_PHC7386_n2582 (.O(FE_PHN7386_n2582), 
	.I(FE_PHN7496_n2582));
   BUFCHD FE_PHC7385_n914 (.O(FE_PHN7385_n914), 
	.I(FE_PHN3504_n914));
   BUFCKEHD FE_PHC7384_n2857 (.O(FE_PHN7384_n2857), 
	.I(FE_PHN4911_n2857));
   BUFCKEHD FE_PHC7383_n901 (.O(FE_PHN7383_n901), 
	.I(FE_PHN3579_n901));
   BUFCHD FE_PHC7382_n1007 (.O(FE_PHN7382_n1007), 
	.I(n1007));
   BUFCHD FE_PHC7381_n2594 (.O(FE_PHN7381_n2594), 
	.I(FE_PHN4892_n2594));
   BUFCHD FE_PHC7380_n996 (.O(FE_PHN7380_n996), 
	.I(FE_PHN5716_n996));
   BUFCHD FE_PHC7379_n2380 (.O(FE_PHN7379_n2380), 
	.I(FE_PHN4797_n2380));
   BUFCHD FE_PHC7378_n2398 (.O(FE_PHN7378_n2398), 
	.I(FE_PHN4811_n2398));
   BUFCHD FE_PHC7377_n4027 (.O(FE_PHN7377_n4027), 
	.I(FE_PHN4391_n4027));
   BUFCKEHD FE_PHC7376_n4210 (.O(FE_PHN7376_n4210), 
	.I(n4210));
   BUFCHD FE_PHC7375_n1054 (.O(FE_PHN7375_n1054), 
	.I(FE_PHN4893_n1054));
   BUFCHD FE_PHC7374_n2696 (.O(FE_PHN7374_n2696), 
	.I(FE_PHN5718_n2696));
   BUFCHD FE_PHC7373_n2172 (.O(FE_PHN7373_n2172), 
	.I(FE_PHN4948_n2172));
   BUFCHD FE_PHC7372_n3965 (.O(FE_PHN7372_n3965), 
	.I(n3965));
   BUFCHD FE_PHC7371_n3212 (.O(FE_PHN7371_n3212), 
	.I(FE_PHN3390_n3212));
   BUFCHD FE_PHC7370_n1922 (.O(FE_PHN7370_n1922), 
	.I(FE_PHN4614_n1922));
   BUFCHD FE_PHC7369_n4308 (.O(FE_PHN7369_n4308), 
	.I(FE_PHN3683_n4308));
   BUFCKEHD FE_PHC7368_n4274 (.O(FE_PHN7368_n4274), 
	.I(FE_PHN3628_n4274));
   BUFCKEHD FE_PHC7367_n1880 (.O(FE_PHN7367_n1880), 
	.I(FE_PHN3833_n1880));
   BUFCHD FE_PHC7366_n985 (.O(FE_PHN7366_n985), 
	.I(n985));
   BUFCHD FE_PHC7365_n2587 (.O(FE_PHN7365_n2587), 
	.I(FE_PHN4820_n2587));
   BUFCHD FE_PHC7364_n2619 (.O(FE_PHN7364_n2619), 
	.I(n2619));
   BUFCKEHD FE_PHC7363_n2181 (.O(FE_PHN7363_n2181), 
	.I(FE_PHN4932_n2181));
   BUFCHD FE_PHC7362_n933 (.O(FE_PHN7362_n933), 
	.I(FE_PHN3463_n933));
   BUFCKEHD FE_PHC7361_n2163 (.O(FE_PHN7361_n2163), 
	.I(FE_PHN3883_n2163));
   BUFCKEHD FE_PHC7360_n4142 (.O(FE_PHN7360_n4142), 
	.I(FE_PHN3465_n4142));
   BUFCHD FE_PHC7359_n1918 (.O(FE_PHN7359_n1918), 
	.I(FE_PHN3893_n1918));
   BUFCHD FE_PHC7358_n2876 (.O(FE_PHN7358_n2876), 
	.I(FE_PHN4916_n2876));
   BUFCHD FE_PHC7357_n1094 (.O(FE_PHN7357_n1094), 
	.I(FE_PHN4844_n1094));
   BUFCHD FE_PHC7356_n1031 (.O(FE_PHN7356_n1031), 
	.I(FE_PHN4902_n1031));
   BUFCHD FE_PHC7355_n3955 (.O(FE_PHN7355_n3955), 
	.I(FE_PHN3780_n3955));
   BUFCHD FE_PHC7354_n3971 (.O(FE_PHN7354_n3971), 
	.I(FE_PHN3587_n3971));
   BUFCHD FE_PHC7353_n2566 (.O(FE_PHN7353_n2566), 
	.I(FE_PHN5692_n2566));
   BUFCKEHD FE_PHC7352_n3932 (.O(FE_PHN7352_n3932), 
	.I(n3932));
   BUFCHD FE_PHC7351_n4110 (.O(FE_PHN7351_n4110), 
	.I(FE_PHN3467_n4110));
   BUFCHD FE_PHC7350_n4018 (.O(FE_PHN7350_n4018), 
	.I(FE_PHN4776_n4018));
   BUFCHD FE_PHC7349_n2428 (.O(FE_PHN7349_n2428), 
	.I(FE_PHN4774_n2428));
   BUFCHD FE_PHC7348_n2388 (.O(FE_PHN7348_n2388), 
	.I(FE_PHN3992_n2388));
   BUFCKEHD FE_PHC7347_n4273 (.O(FE_PHN7347_n4273), 
	.I(FE_PHN3947_n4273));
   BUFCKEHD FE_PHC7346_n3970 (.O(FE_PHN7346_n3970), 
	.I(n3970));
   BUFCHD FE_PHC7345_n1874 (.O(FE_PHN7345_n1874), 
	.I(FE_PHN6495_n1874));
   BUFCHD FE_PHC7344_n2747 (.O(FE_PHN7344_n2747), 
	.I(FE_PHN4941_n2747));
   BUFCHD FE_PHC7343_n2618 (.O(FE_PHN7343_n2618), 
	.I(FE_PHN4815_n2618));
   BUFCHD FE_PHC7342_n2432 (.O(FE_PHN7342_n2432), 
	.I(FE_PHN3607_n2432));
   BUFCHD FE_PHC7341_n2695 (.O(FE_PHN7341_n2695), 
	.I(FE_PHN4865_n2695));
   BUFCHD FE_PHC7340_n4116 (.O(FE_PHN7340_n4116), 
	.I(FE_PHN3606_n4116));
   BUFCHD FE_PHC7339_n2121 (.O(FE_PHN7339_n2121), 
	.I(FE_PHN4822_n2121));
   BUFCHD FE_PHC7338_n2149 (.O(FE_PHN7338_n2149), 
	.I(FE_PHN4788_n2149));
   BUFCHD FE_PHC7337_n1015 (.O(FE_PHN7337_n1015), 
	.I(FE_PHN4876_n1015));
   BUFCHD FE_PHC7336_n4294 (.O(FE_PHN7336_n4294), 
	.I(FE_PHN3574_n4294));
   BUFCHD FE_PHC7335_n2611 (.O(FE_PHN7335_n2611), 
	.I(FE_PHN4912_n2611));
   BUFCKEHD FE_PHC7334_n953 (.O(FE_PHN7334_n953), 
	.I(FE_PHN4838_n953));
   BUFCHD FE_PHC7333_n1190 (.O(FE_PHN7333_n1190), 
	.I(FE_PHN4934_n1190));
   BUFCHD FE_PHC7332_n2412 (.O(FE_PHN7332_n2412), 
	.I(FE_PHN4781_n2412));
   BUFCHD FE_PHC7331_n2750 (.O(FE_PHN7331_n2750), 
	.I(FE_PHN4918_n2750));
   BUFCKEHD FE_PHC7330_n1919 (.O(FE_PHN7330_n1919), 
	.I(FE_PHN3792_n1919));
   BUFCHD FE_PHC7329_n1872 (.O(FE_PHN7329_n1872), 
	.I(FE_PHN3469_n1872));
   BUFCHD FE_PHC7328_n1906 (.O(FE_PHN7328_n1906), 
	.I(FE_PHN3831_n1906));
   BUFCKEHD FE_PHC7327_n2602 (.O(FE_PHN7327_n2602), 
	.I(FE_PHN4793_n2602));
   BUFCKEHD FE_PHC7326_n950 (.O(FE_PHN7326_n950), 
	.I(FE_PHN4233_n950));
   BUFCHD FE_PHC7325_n2576 (.O(FE_PHN7325_n2576), 
	.I(FE_PHN4883_n2576));
   BUFCHD FE_PHC7324_n1178 (.O(FE_PHN7324_n1178), 
	.I(FE_PHN4939_n1178));
   BUFCKEHD FE_PHC7323_n2124 (.O(FE_PHN7323_n2124), 
	.I(FE_PHN4828_n2124));
   BUFCHD FE_PHC7322_n4148 (.O(FE_PHN7322_n4148), 
	.I(FE_PHN3689_n4148));
   BUFCHD FE_PHC7321_n906 (.O(FE_PHN7321_n906), 
	.I(FE_PHN3836_n906));
   BUFCHD FE_PHC7320_n964 (.O(FE_PHN7320_n964), 
	.I(FE_PHN3585_n964));
   BUFCKEHD FE_PHC7319_n979 (.O(FE_PHN7319_n979), 
	.I(FE_PHN7460_n979));
   BUFCHD FE_PHC7318_n2622 (.O(FE_PHN7318_n2622), 
	.I(FE_PHN4931_n2622));
   BUFCHD FE_PHC7317_n2572 (.O(FE_PHN7317_n2572), 
	.I(FE_PHN4885_n2572));
   BUFCKEHD FE_PHC7316_n2138 (.O(FE_PHN7316_n2138), 
	.I(FE_PHN4825_n2138));
   BUFCHD FE_PHC7315_n2612 (.O(FE_PHN7315_n2612), 
	.I(FE_PHN4852_n2612));
   BUFCHD FE_PHC7314_n4114 (.O(FE_PHN7314_n4114), 
	.I(FE_PHN6506_n4114));
   BUFCHD FE_PHC7313_n1154 (.O(FE_PHN7313_n1154), 
	.I(FE_PHN7459_n1154));
   BUFCHD FE_PHC7312_n2251 (.O(FE_PHN7312_n2251), 
	.I(FE_PHN4945_n2251));
   BUFCHD FE_PHC7311_n938 (.O(FE_PHN7311_n938), 
	.I(FE_PHN7458_n938));
   BUFCHD FE_PHC7310_n1001 (.O(FE_PHN7310_n1001), 
	.I(FE_PHN7494_n1001));
   BUFCKEHD FE_PHC7309_n4046 (.O(FE_PHN7309_n4046), 
	.I(FE_PHN3927_n4046));
   BUFCHD FE_PHC7308_n3072 (.O(FE_PHN7308_n3072), 
	.I(n3072));
   BUFCKEHD FE_PHC7307_n3052 (.O(n3052), 
	.I(FE_PHN7307_n3052));
   BUFCHD FE_PHC7306_n2564 (.O(FE_PHN7306_n2564), 
	.I(FE_PHN3949_n2564));
   BUFCHD FE_PHC7305_n4180 (.O(FE_PHN7305_n4180), 
	.I(FE_PHN5908_n4180));
   BUFCHD FE_PHC7304_n928 (.O(FE_PHN7304_n928), 
	.I(FE_PHN3744_n928));
   BUFCHD FE_PHC7303_n905 (.O(FE_PHN7303_n905), 
	.I(FE_PHN3861_n905));
   BUFCHD FE_PHC7302_n3919 (.O(FE_PHN7302_n3919), 
	.I(FE_PHN4432_n3919));
   BUFCHD FE_PHC7301_n4215 (.O(FE_PHN7301_n4215), 
	.I(n4215));
   BUFCKEHD FE_PHC7300_n4219 (.O(FE_PHN7300_n4219), 
	.I(FE_PHN5955_n4219));
   BUFCHD FE_PHC7299_n2574 (.O(FE_PHN7299_n2574), 
	.I(FE_PHN3821_n2574));
   BUFCHD FE_PHC7298_n4174 (.O(FE_PHN7298_n4174), 
	.I(n4174));
   BUFCKEHD FE_PHC7297_n975 (.O(FE_PHN7297_n975), 
	.I(n975));
   BUFCHD FE_PHC7296_n2599 (.O(FE_PHN7296_n2599), 
	.I(FE_PHN3700_n2599));
   BUFCHD FE_PHC7295_n1082 (.O(FE_PHN7295_n1082), 
	.I(n1082));
   BUFCHD FE_PHC7294_n948 (.O(FE_PHN7294_n948), 
	.I(FE_PHN3471_n948));
   BUFCKEHD FE_PHC7293_n3129 (.O(n3129), 
	.I(FE_PHN7293_n3129));
   BUFCHD FE_PHC7292_n2580 (.O(FE_PHN7292_n2580), 
	.I(FE_PHN3920_n2580));
   BUFCHD FE_PHC7291_n3028 (.O(FE_PHN7291_n3028), 
	.I(FE_PHN7452_n3028));
   BUFCHD FE_PHC7290_n1017 (.O(FE_PHN7290_n1017), 
	.I(FE_PHN7450_n1017));
   BUFCHD FE_PHC7289_n4229 (.O(FE_PHN7289_n4229), 
	.I(n4229));
   BUFCKEHD FE_PHC7288_n1014 (.O(FE_PHN7288_n1014), 
	.I(FE_PHN7502_n1014));
   BUFCHD FE_PHC7287_n3964 (.O(FE_PHN7287_n3964), 
	.I(FE_PHN7493_n3964));
   BUFCHD FE_PHC7286_n974 (.O(FE_PHN7286_n974), 
	.I(FE_PHN7491_n974));
   BUFCKEHD FE_PHC7285_n1013 (.O(FE_PHN7285_n1013), 
	.I(n1013));
   BUFCHD FE_PHC7284_n4365 (.O(FE_PHN7284_n4365), 
	.I(FE_PHN3667_n4365));
   BUFCKEHD FE_PHC7283_n2972 (.O(FE_PHN7283_n2972), 
	.I(n2972));
   BUFEHD FE_PHC7282_n4409 (.O(FE_PHN7282_n4409), 
	.I(FE_PHN3770_n4409));
   BUFEHD FE_PHC7281_n3068 (.O(FE_PHN7281_n3068), 
	.I(FE_PHN7442_n3068));
   BUFEHD FE_PHC7280_n2887 (.O(FE_PHN7280_n2887), 
	.I(n2887));
   BUFCKEHD FE_PHC7279_n2426 (.O(FE_PHN7279_n2426), 
	.I(FE_PHN7448_n2426));
   BUFEHD FE_PHC7278_n4013 (.O(FE_PHN7278_n4013), 
	.I(FE_PHN7447_n4013));
   BUFCKIHD FE_PHC7277_n2133 (.O(FE_PHN7277_n2133), 
	.I(FE_PHN7444_n2133));
   BUFEHD FE_PHC7276_n2892 (.O(FE_PHN7276_n2892), 
	.I(FE_PHN7423_n2892));
   BUFCKEHD FE_PHC7275_n2425 (.O(FE_PHN7275_n2425), 
	.I(FE_PHN4790_n2425));
   BUFCKEHD FE_PHC7274_n2379 (.O(FE_PHN7274_n2379), 
	.I(FE_PHN7435_n2379));
   BUFCKEHD FE_PHC7273_n2377 (.O(FE_PHN7273_n2377), 
	.I(FE_PHN4827_n2377));
   BUFCKEHD FE_PHC7272_n4011 (.O(FE_PHN7272_n4011), 
	.I(FE_PHN4787_n4011));
   BUFCHD FE_PHC7271_n2119 (.O(FE_PHN7271_n2119), 
	.I(FE_PHN7446_n2119));
   BUFCHD FE_PHC7270_n2151 (.O(FE_PHN7270_n2151), 
	.I(FE_PHN7438_n2151));
   BUFCKEHD FE_PHC7269_n2427 (.O(FE_PHN7269_n2427), 
	.I(FE_PHN4829_n2427));
   BUFCKEHD FE_PHC7268_n2126 (.O(FE_PHN7268_n2126), 
	.I(FE_PHN7440_n2126));
   BUFCKEHD FE_PHC7267_n2395 (.O(FE_PHN7267_n2395), 
	.I(FE_PHN7397_n2395));
   BUFEHD FE_PHC7266_n4002 (.O(FE_PHN7266_n4002), 
	.I(FE_PHN4958_n4002));
   BUFCKEHD FE_PHC7265_n2603 (.O(FE_PHN7265_n2603), 
	.I(FE_PHN7432_n2603));
   BUFCKEHD FE_PHC7264_n2434 (.O(FE_PHN7264_n2434), 
	.I(FE_PHN7421_n2434));
   BUFCKEHD FE_PHC7263_n2610 (.O(FE_PHN7263_n2610), 
	.I(FE_PHN7437_n2610));
   BUFCHD FE_PHC7262_n3953 (.O(FE_PHN7262_n3953), 
	.I(FE_PHN7428_n3953));
   BUFCKEHD FE_PHC7261_n2570 (.O(FE_PHN7261_n2570), 
	.I(FE_PHN7422_n2570));
   BUFCKEHD FE_PHC7260_n2135 (.O(FE_PHN7260_n2135), 
	.I(FE_PHN7431_n2135));
   BUFEHD FE_PHC7259_n2179 (.O(FE_PHN7259_n2179), 
	.I(FE_PHN7427_n2179));
   BUFCKEHD FE_PHC7258_n2378 (.O(FE_PHN7258_n2378), 
	.I(FE_PHN7439_n2378));
   BUFCHD FE_PHC7257_n2165 (.O(FE_PHN7257_n2165), 
	.I(FE_PHN7436_n2165));
   BUFCHD FE_PHC7256_n2168 (.O(FE_PHN7256_n2168), 
	.I(FE_PHN7424_n2168));
   BUFCHD FE_PHC7255_n2175 (.O(FE_PHN7255_n2175), 
	.I(FE_PHN7415_n2175));
   BUFCHD FE_PHC7254_n2118 (.O(FE_PHN7254_n2118), 
	.I(FE_PHN7434_n2118));
   BUFCKEHD FE_PHC7253_n2393 (.O(FE_PHN7253_n2393), 
	.I(FE_PHN7445_n2393));
   BUFCHD FE_PHC7252_n2169 (.O(FE_PHN7252_n2169), 
	.I(FE_PHN7429_n2169));
   BUFCKEHD FE_PHC7251_n2152 (.O(FE_PHN7251_n2152), 
	.I(FE_PHN7417_n2152));
   BUFCKLHD FE_PHC7250_n2164 (.O(FE_PHN7250_n2164), 
	.I(FE_PHN7441_n2164));
   BUFCKEHD FE_PHC7249_n2890 (.O(n2890), 
	.I(FE_PHN7249_n2890));
   BUFEHD FE_PHC7248_n2120 (.O(FE_PHN7248_n2120), 
	.I(FE_PHN7412_n2120));
   BUFCHD FE_PHC7247_n3934 (.O(FE_PHN7247_n3934), 
	.I(FE_PHN7426_n3934));
   BUFCKEHD FE_PHC7246_n2571 (.O(FE_PHN7246_n2571), 
	.I(FE_PHN7407_n2571));
   BUFCKEHD FE_PHC7245_n4153 (.O(FE_PHN7245_n4153), 
	.I(FE_PHN4780_n4153));
   BUFCHD FE_PHC7244_n2410 (.O(FE_PHN7244_n2410), 
	.I(FE_PHN7418_n2410));
   BUFCHD FE_PHC7243_n3960 (.O(FE_PHN7243_n3960), 
	.I(FE_PHN7406_n3960));
   BUFCHD FE_PHC7242_n4137 (.O(FE_PHN7242_n4137), 
	.I(FE_PHN7472_n4137));
   BUFCKEHD FE_PHC7241_n2578 (.O(FE_PHN7241_n2578), 
	.I(FE_PHN7402_n2578));
   BUFCHD FE_PHC7240_n3923 (.O(FE_PHN7240_n3923), 
	.I(FE_PHN7404_n3923));
   BUFEHD FE_PHC7239_n2132 (.O(FE_PHN7239_n2132), 
	.I(FE_PHN7416_n2132));
   BUFCHD FE_PHC7238_n3230 (.O(FE_PHN7238_n3230), 
	.I(FE_PHN7395_n3230));
   BUFEHD FE_PHC7237_n3968 (.O(FE_PHN7237_n3968), 
	.I(FE_PHN7420_n3968));
   BUFCKEHD FE_PHC7236_n2417 (.O(FE_PHN7236_n2417), 
	.I(FE_PHN7387_n2417));
   BUFCHD FE_PHC7235_n4155 (.O(FE_PHN7235_n4155), 
	.I(FE_PHN7419_n4155));
   BUFCHD FE_PHC7234_n2167 (.O(FE_PHN7234_n2167), 
	.I(FE_PHN7433_n2167));
   BUFCKIHD FE_PHC7233_n4121 (.O(FE_PHN7233_n4121), 
	.I(FE_PHN7410_n4121));
   BUFCHD FE_PHC7232_n2155 (.O(FE_PHN7232_n2155), 
	.I(FE_PHN7405_n2155));
   BUFCHD FE_PHC7231_n2154 (.O(FE_PHN7231_n2154), 
	.I(FE_PHN7425_n2154));
   BUFLHD FE_PHC7230_n2180 (.O(FE_PHN7230_n2180), 
	.I(n2180));
   BUFCHD FE_PHC7229_n2394 (.O(FE_PHN7229_n2394), 
	.I(FE_PHN7414_n2394));
   BUFEHD FE_PHC7228_n2402 (.O(FE_PHN7228_n2402), 
	.I(FE_PHN7408_n2402));
   BUFCHD FE_PHC7227_n2625 (.O(FE_PHN7227_n2625), 
	.I(FE_PHN7403_n2625));
   BUFCHD FE_PHC7226_n2159 (.O(FE_PHN7226_n2159), 
	.I(FE_PHN7400_n2159));
   BUFCHD FE_PHC7225_n2170 (.O(FE_PHN7225_n2170), 
	.I(FE_PHN7413_n2170));
   BUFCKEHD FE_PHC7224_n2582 (.O(FE_PHN7224_n2582), 
	.I(FE_PHN7386_n2582));
   BUFMHD FE_PHC7223_n4139 (.O(FE_PHN7223_n4139), 
	.I(FE_PHN4861_n4139));
   BUFCHD FE_PHC7222_n4147 (.O(FE_PHN7222_n4147), 
	.I(FE_PHN7392_n4147));
   BUFCKGHD FE_PHC7221_n2166 (.O(FE_PHN7221_n2166), 
	.I(FE_PHN7398_n2166));
   BUFCHD FE_PHC7220_n2592 (.O(FE_PHN7220_n2592), 
	.I(FE_PHN7396_n2592));
   BUFCHD FE_PHC7219_n2628 (.O(FE_PHN7219_n2628), 
	.I(FE_PHN7411_n2628));
   BUFCKLHD FE_PHC7218_n1863 (.O(FE_PHN7218_n1863), 
	.I(FE_PHN7401_n1863));
   BUFCKGHD FE_PHC7217_n2614 (.O(FE_PHN7217_n2614), 
	.I(FE_PHN7393_n2614));
   BUFCKGHD FE_PHC7216_n4102 (.O(FE_PHN7216_n4102), 
	.I(FE_PHN7389_n4102));
   BUFCHD FE_PHC7215_n4163 (.O(FE_PHN7215_n4163), 
	.I(FE_PHN7394_n4163));
   BUFCHD FE_PHC7214_n2130 (.O(FE_PHN7214_n2130), 
	.I(FE_PHN7391_n2130));
   BUFCKMHD FE_PHC7213_n2604 (.O(FE_PHN7213_n2604), 
	.I(FE_PHN7443_n2604));
   BUFCHD FE_PHC7212_n3150 (.O(FE_PHN7212_n3150), 
	.I(FE_PHN4960_n3150));
   BUFCKEHD FE_PHC7211_n4135 (.O(FE_PHN7211_n4135), 
	.I(FE_PHN4835_n4135));
   BUFCKEHD FE_PHC7210_n880 (.O(FE_PHN7210_n880), 
	.I(FE_PHN3771_n880));
   BUFCHD FE_PHC7209_n1913 (.O(FE_PHN7209_n1913), 
	.I(FE_PHN4959_n1913));
   BUFCHD FE_PHC7208_n2422 (.O(FE_PHN7208_n2422), 
	.I(n2422));
   BUFCKEHD FE_PHC7207_n4107 (.O(FE_PHN7207_n4107), 
	.I(FE_PHN4878_n4107));
   BUFCKEHD FE_PHC7206_n3017 (.O(FE_PHN7206_n3017), 
	.I(n3017));
   BUFCKEHD FE_PHC7205_n1086 (.O(FE_PHN7205_n1086), 
	.I(FE_PHN4951_n1086));
   BUFCHD FE_PHC7204_n4016 (.O(FE_PHN7204_n4016), 
	.I(FE_PHN3680_n4016));
   BUFCHD FE_PHC7203_n2697 (.O(FE_PHN7203_n2697), 
	.I(FE_PHN4879_n2697));
   BUFCHD FE_PHC7202_n3944 (.O(FE_PHN7202_n3944), 
	.I(FE_PHN3450_n3944));
   BUFCKEHD FE_PHC7201_n3962 (.O(FE_PHN7201_n3962), 
	.I(FE_PHN3966_n3962));
   BUFCHD FE_PHC7200_n921 (.O(FE_PHN7200_n921), 
	.I(FE_PHN4946_n921));
   BUFCKEHD FE_PHC7199_n2609 (.O(FE_PHN7199_n2609), 
	.I(FE_PHN4855_n2609));
   BUFCKEHD FE_PHC7198_n2123 (.O(FE_PHN7198_n2123), 
	.I(FE_PHN4900_n2123));
   BUFCHD FE_PHC7197_n2177 (.O(FE_PHN7197_n2177), 
	.I(FE_PHN4926_n2177));
   BUFCKEHD FE_PHC7196_n2589 (.O(FE_PHN7196_n2589), 
	.I(FE_PHN4887_n2589));
   BUFCKEHD FE_PHC7195_n2743 (.O(FE_PHN7195_n2743), 
	.I(FE_PHN4924_n2743));
   BUFCHD FE_PHC7194_n2873 (.O(FE_PHN7194_n2873), 
	.I(FE_PHN5685_n2873));
   BUFCHD FE_PHC7193_n1028 (.O(FE_PHN7193_n1028), 
	.I(FE_PHN4929_n1028));
   BUFCHD FE_PHC7192_n973 (.O(FE_PHN7192_n973), 
	.I(FE_PHN4935_n973));
   BUFCKEHD FE_PHC7191_n2749 (.O(FE_PHN7191_n2749), 
	.I(FE_PHN4896_n2749));
   BUFCKEHD FE_PHC7190_n3047 (.O(FE_PHN7190_n3047), 
	.I(n3047));
   BUFCKEHD FE_PHC7189_n3021 (.O(FE_PHN7189_n3021), 
	.I(FE_PHN5735_n3021));
   BUFCHD FE_PHC7188_n2171 (.O(FE_PHN7188_n2171), 
	.I(FE_PHN4813_n2171));
   BUFCHD FE_PHC7187_n1908 (.O(FE_PHN7187_n1908), 
	.I(FE_PHN4933_n1908));
   BUFCKEHD FE_PHC7186_n2590 (.O(FE_PHN7186_n2590), 
	.I(FE_PHN4910_n2590));
   BUFCKEHD FE_PHC7185_n2381 (.O(FE_PHN7185_n2381), 
	.I(FE_PHN4905_n2381));
   BUFCHD FE_PHC7184_n2122 (.O(FE_PHN7184_n2122), 
	.I(FE_PHN4826_n2122));
   BUFCKEHD FE_PHC7183_n2935 (.O(FE_PHN7183_n2935), 
	.I(FE_PHN4359_n2935));
   BUFCHD FE_PHC7182_n4151 (.O(FE_PHN7182_n4151), 
	.I(FE_PHN4805_n4151));
   BUFCKEHD FE_PHC7181_n1375 (.O(FE_PHN7181_n1375), 
	.I(FE_PHN6618_n1375));
   BUFCKEHD FE_PHC7180_n2616 (.O(FE_PHN7180_n2616), 
	.I(FE_PHN4858_n2616));
   BUFCKEHD FE_PHC7179_n1012 (.O(FE_PHN7179_n1012), 
	.I(FE_PHN4943_n1012));
   BUFCKEHD FE_PHC7178_n967 (.O(FE_PHN7178_n967), 
	.I(FE_PHN4928_n967));
   BUFCHD FE_PHC7177_n981 (.O(FE_PHN7177_n981), 
	.I(FE_PHN5740_n981));
   BUFCHD FE_PHC7176_n2624 (.O(FE_PHN7176_n2624), 
	.I(FE_PHN4906_n2624));
   BUFCHD FE_PHC7175_n2919 (.O(FE_PHN7175_n2919), 
	.I(FE_PHN4897_n2919));
   BUFCKEHD FE_PHC7174_n4008 (.O(FE_PHN7174_n4008), 
	.I(FE_PHN3237_n4008));
   BUFCKEHD FE_PHC7173_n4158 (.O(FE_PHN7173_n4158), 
	.I(FE_PHN3786_n4158));
   BUFCHD FE_PHC7172_n2176 (.O(FE_PHN7172_n2176), 
	.I(FE_PHN4796_n2176));
   BUFCKEHD FE_PHC7171_n2904 (.O(FE_PHN7171_n2904), 
	.I(FE_PHN4314_n2904));
   BUFCKEHD FE_PHC7170_n2701 (.O(FE_PHN7170_n2701), 
	.I(FE_PHN4856_n2701));
   BUFDHD FE_PHC7169_n4404 (.O(FE_PHN7169_n4404), 
	.I(FE_PHN3597_n4404));
   BUFCHD FE_PHC7168_n4331 (.O(FE_PHN7168_n4331), 
	.I(FE_PHN3483_n4331));
   BUFCKEHD FE_PHC7167_n1865 (.O(FE_PHN7167_n1865), 
	.I(FE_PHN6613_n1865));
   BUFCKEHD FE_PHC7166_n2908 (.O(FE_PHN7166_n2908), 
	.I(FE_PHN6617_n2908));
   BUFCKEHD FE_PHC7165_n3033 (.O(FE_PHN7165_n3033), 
	.I(n3033));
   BUFCKEHD FE_PHC7164_n2889 (.O(FE_PHN7164_n2889), 
	.I(n2889));
   BUFCKEHD FE_PHC7163_n4259 (.O(FE_PHN7163_n4259), 
	.I(FE_PHN3925_n4259));
   BUFCHD FE_PHC7162_n3965 (.O(FE_PHN7162_n3965), 
	.I(FE_PHN7372_n3965));
   BUFCHD FE_PHC7161_n4358 (.O(FE_PHN7161_n4358), 
	.I(FE_PHN3319_n4358));
   BUFCKEHD FE_PHC7160_n1158 (.O(FE_PHN7160_n1158), 
	.I(FE_PHN6564_n1158));
   BUFCKEHD FE_PHC7159_n4035 (.O(FE_PHN7159_n4035), 
	.I(FE_PHN3750_n4035));
   BUFCHD FE_PHC7158_n4150 (.O(FE_PHN7158_n4150), 
	.I(FE_PHN4818_n4150));
   BUFCKEHD FE_PHC7157_n4062 (.O(FE_PHN7157_n4062), 
	.I(FE_PHN3748_n4062));
   BUFCKEHD FE_PHC7156_n2386 (.O(FE_PHN7156_n2386), 
	.I(FE_PHN6612_n2386));
   BUFCHD FE_PHC7155_n3945 (.O(FE_PHN7155_n3945), 
	.I(FE_PHN3498_n3945));
   BUFCHD FE_PHC7154_n2922 (.O(FE_PHN7154_n2922), 
	.I(FE_PHN3754_n2922));
   BUFCKEHD FE_PHC7153_n3212 (.O(FE_PHN7153_n3212), 
	.I(FE_PHN7371_n3212));
   BUFCKEHD FE_PHC7152_n2390 (.O(FE_PHN7152_n2390), 
	.I(FE_PHN6609_n2390));
   BUFEHD FE_PHC7151_n1007 (.O(FE_PHN7151_n1007), 
	.I(FE_PHN7382_n1007));
   BUFCHD FE_PHC7150_n2893 (.O(FE_PHN7150_n2893), 
	.I(FE_PHN4841_n2893));
   BUFCHD FE_PHC7149_n1286 (.O(FE_PHN7149_n1286), 
	.I(FE_PHN4925_n1286));
   BUFCHD FE_PHC7148_n2907 (.O(FE_PHN7148_n2907), 
	.I(FE_PHN4799_n2907));
   BUFCHD FE_PHC7147_n1019 (.O(FE_PHN7147_n1019), 
	.I(FE_PHN4957_n1019));
   BUFCHD FE_PHC7146_n2626 (.O(FE_PHN7146_n2626), 
	.I(FE_PHN4849_n2626));
   BUFCHD FE_PHC7145_n1003 (.O(FE_PHN7145_n1003), 
	.I(FE_PHN4907_n1003));
   BUFCKEHD FE_PHC7144_n888 (.O(FE_PHN7144_n888), 
	.I(FE_PHN3813_n888));
   BUFCKEHD FE_PHC7143_n4308 (.O(FE_PHN7143_n4308), 
	.I(FE_PHN7369_n4308));
   BUFCHD FE_PHC7142_n2161 (.O(FE_PHN7142_n2161), 
	.I(FE_PHN4884_n2161));
   BUFCHD FE_PHC7141_n4034 (.O(FE_PHN7141_n4034), 
	.I(FE_PHN3516_n4034));
   BUFCHD FE_PHC7140_n2925 (.O(FE_PHN7140_n2925), 
	.I(FE_PHN4783_n2925));
   BUFCHD FE_PHC7139_n2144 (.O(FE_PHN7139_n2144), 
	.I(FE_PHN5655_n2144));
   BUFCKEHD FE_PHC7138_n2432 (.O(FE_PHN7138_n2432), 
	.I(FE_PHN7342_n2432));
   BUFCKEHD FE_PHC7137_n3979 (.O(FE_PHN7137_n3979), 
	.I(FE_PHN3442_n3979));
   BUFEHD FE_PHC7136_n4210 (.O(FE_PHN7136_n4210), 
	.I(FE_PHN7376_n4210));
   BUFCKEHD FE_PHC7135_n4032 (.O(FE_PHN7135_n4032), 
	.I(FE_PHN4449_n4032));
   BUFEHD FE_PHC7134_n2938 (.O(FE_PHN7134_n2938), 
	.I(n2938));
   BUFCHD FE_PHC7133_n4012 (.O(FE_PHN7133_n4012), 
	.I(FE_PHN4784_n4012));
   BUFCKEHD FE_PHC7132_n2403 (.O(FE_PHN7132_n2403), 
	.I(FE_PHN4418_n2403));
   BUFCHD FE_PHC7131_n2941 (.O(FE_PHN7131_n2941), 
	.I(FE_PHN4786_n2941));
   BUFEHD FE_PHC7130_n901 (.O(FE_PHN7130_n901), 
	.I(FE_PHN7383_n901));
   BUFCHD FE_PHC7129_n985 (.O(FE_PHN7129_n985), 
	.I(FE_PHN7366_n985));
   BUFCHD FE_PHC7128_n2375 (.O(FE_PHN7128_n2375), 
	.I(FE_PHN4837_n2375));
   BUFCHD FE_PHC7127_n983 (.O(FE_PHN7127_n983), 
	.I(FE_PHN4794_n983));
   BUFEHD FE_PHC7126_n996 (.O(FE_PHN7126_n996), 
	.I(FE_PHN7380_n996));
   BUFCHD FE_PHC7125_n2125 (.O(FE_PHN7125_n2125), 
	.I(FE_PHN4914_n2125));
   BUFCHD FE_PHC7124_n4242 (.O(FE_PHN7124_n4242), 
	.I(FE_PHN3910_n4242));
   BUFCHD FE_PHC7123_n2696 (.O(FE_PHN7123_n2696), 
	.I(FE_PHN7374_n2696));
   BUFEHD FE_PHC7122_n4274 (.O(FE_PHN7122_n4274), 
	.I(FE_PHN7368_n4274));
   BUFCHD FE_PHC7121_n2857 (.O(FE_PHN7121_n2857), 
	.I(FE_PHN7384_n2857));
   BUFCHD FE_PHC7120_n3983 (.O(FE_PHN7120_n3983), 
	.I(FE_PHN3342_n3983));
   BUFCHD FE_PHC7119_n2587 (.O(FE_PHN7119_n2587), 
	.I(FE_PHN7365_n2587));
   BUFCHD FE_PHC7118_n917 (.O(FE_PHN7118_n917), 
	.I(FE_PHN3432_n917));
   BUFCKEHD FE_PHC7117_n3260 (.O(FE_PHN7117_n3260), 
	.I(FE_PHN3388_n3260));
   BUFCHD FE_PHC7116_n2257 (.O(FE_PHN7116_n2257), 
	.I(FE_PHN4954_n2257));
   BUFCHD FE_PHC7115_n3980 (.O(FE_PHN7115_n3980), 
	.I(FE_PHN3741_n3980));
   BUFCKEHD FE_PHC7114_n1906 (.O(FE_PHN7114_n1906), 
	.I(FE_PHN7328_n1906));
   BUFCKEHD FE_PHC7113_n4031 (.O(FE_PHN7113_n4031), 
	.I(FE_PHN3406_n4031));
   BUFCHD FE_PHC7112_n2398 (.O(FE_PHN7112_n2398), 
	.I(FE_PHN7378_n2398));
   BUFCKEHD FE_PHC7111_n2876 (.O(FE_PHN7111_n2876), 
	.I(FE_PHN7358_n2876));
   BUFEHD FE_PHC7110_n962 (.O(FE_PHN7110_n962), 
	.I(FE_PHN3803_n962));
   BUFCHD FE_PHC7109_n930 (.O(FE_PHN7109_n930), 
	.I(FE_PHN3401_n930));
   BUFCHD FE_PHC7108_n933 (.O(FE_PHN7108_n933), 
	.I(FE_PHN7362_n933));
   BUFCHD FE_PHC7107_n914 (.O(FE_PHN7107_n914), 
	.I(FE_PHN7385_n914));
   BUFEHD FE_PHC7106_n2577 (.O(FE_PHN7106_n2577), 
	.I(n2577));
   BUFCHD FE_PHC7105_n2424 (.O(FE_PHN7105_n2424), 
	.I(FE_PHN4833_n2424));
   BUFCHD FE_PHC7104_n949 (.O(FE_PHN7104_n949), 
	.I(FE_PHN3832_n949));
   BUFCHD FE_PHC7103_n2407 (.O(FE_PHN7103_n2407), 
	.I(FE_PHN4807_n2407));
   BUFCHD FE_PHC7102_n2148 (.O(FE_PHN7102_n2148), 
	.I(FE_PHN4806_n2148));
   BUFCHD FE_PHC7101_n2695 (.O(FE_PHN7101_n2695), 
	.I(FE_PHN7341_n2695));
   BUFCHD FE_PHC7100_n1054 (.O(FE_PHN7100_n1054), 
	.I(FE_PHN7375_n1054));
   BUFEHD FE_PHC7099_n2566 (.O(FE_PHN7099_n2566), 
	.I(FE_PHN7353_n2566));
   BUFEHD FE_PHC7098_n4273 (.O(FE_PHN7098_n4273), 
	.I(FE_PHN7347_n4273));
   BUFCKGHD FE_PHC7097_n1031 (.O(FE_PHN7097_n1031), 
	.I(FE_PHN7356_n1031));
   BUFCKEHD FE_PHC7096_n2419 (.O(FE_PHN7096_n2419), 
	.I(FE_PHN3921_n2419));
   BUFCHD FE_PHC7095_n2181 (.O(FE_PHN7095_n2181), 
	.I(FE_PHN7363_n2181));
   BUFCHD FE_PHC7094_n980 (.O(FE_PHN7094_n980), 
	.I(FE_PHN4834_n980));
   BUFCKEHD FE_PHC7093_n2615 (.O(FE_PHN7093_n2615), 
	.I(FE_PHN4940_n2615));
   BUFCHD FE_PHC7092_n3981 (.O(FE_PHN7092_n3981), 
	.I(FE_PHN4831_n3981));
   BUFCHD FE_PHC7091_n2747 (.O(FE_PHN7091_n2747), 
	.I(FE_PHN7344_n2747));
   BUFCKEHD FE_PHC7090_n4027 (.O(FE_PHN7090_n4027), 
	.I(FE_PHN7377_n4027));
   BUFCHD FE_PHC7089_n3971 (.O(FE_PHN7089_n3971), 
	.I(FE_PHN7354_n3971));
   BUFCKEHD FE_PHC7088_n2163 (.O(FE_PHN7088_n2163), 
	.I(FE_PHN7361_n2163));
   BUFCHD FE_PHC7087_n3966 (.O(FE_PHN7087_n3966), 
	.I(FE_PHN3720_n3966));
   BUFEHD FE_PHC7086_n2750 (.O(FE_PHN7086_n2750), 
	.I(FE_PHN7331_n2750));
   BUFCHD FE_PHC7085_n4294 (.O(FE_PHN7085_n4294), 
	.I(FE_PHN7336_n4294));
   BUFCHD FE_PHC7084_n2406 (.O(FE_PHN7084_n2406), 
	.I(n2406));
   BUFCHD FE_PHC7083_n2429 (.O(FE_PHN7083_n2429), 
	.I(FE_PHN5648_n2429));
   BUFCKEHD FE_PHC7082_n2382 (.O(FE_PHN7082_n2382), 
	.I(FE_PHN4830_n2382));
   BUFCHD FE_PHC7081_n2172 (.O(FE_PHN7081_n2172), 
	.I(FE_PHN7373_n2172));
   BUFEHD FE_PHC7080_n3970 (.O(FE_PHN7080_n3970), 
	.I(FE_PHN7346_n3970));
   BUFCHD FE_PHC7079_n2121 (.O(FE_PHN7079_n2121), 
	.I(FE_PHN7339_n2121));
   BUFCKEHD FE_PHC7078_n2131 (.O(FE_PHN7078_n2131), 
	.I(FE_PHN3452_n2131));
   BUFEHD FE_PHC7077_n3955 (.O(FE_PHN7077_n3955), 
	.I(FE_PHN7355_n3955));
   BUFCHD FE_PHC7076_n2619 (.O(FE_PHN7076_n2619), 
	.I(FE_PHN7364_n2619));
   BUFCKEHD FE_PHC7075_n4018 (.O(FE_PHN7075_n4018), 
	.I(FE_PHN7350_n4018));
   BUFCKGHD FE_PHC7074_n979 (.O(FE_PHN7074_n979), 
	.I(FE_PHN7319_n979));
   BUFCKEHD FE_PHC7073_n2401 (.O(FE_PHN7073_n2401), 
	.I(FE_PHN4798_n2401));
   BUFCKEHD FE_PHC7072_n2156 (.O(FE_PHN7072_n2156), 
	.I(FE_PHN4821_n2156));
   BUFCHD FE_PHC7071_n1015 (.O(FE_PHN7071_n1015), 
	.I(FE_PHN7337_n1015));
   BUFCHD FE_PHC7070_n2376 (.O(FE_PHN7070_n2376), 
	.I(FE_PHN4854_n2376));
   BUFCKEHD FE_PHC7069_n1190 (.O(FE_PHN7069_n1190), 
	.I(FE_PHN7333_n1190));
   BUFCHD FE_PHC7068_n2380 (.O(FE_PHN7068_n2380), 
	.I(FE_PHN7379_n2380));
   BUFCHD FE_PHC7067_n927 (.O(FE_PHN7067_n927), 
	.I(FE_PHN3566_n927));
   BUFCHD FE_PHC7066_n2428 (.O(FE_PHN7066_n2428), 
	.I(FE_PHN7349_n2428));
   BUFCKKHD FE_PHC7065_n944 (.O(FE_PHN7065_n944), 
	.I(FE_PHN3976_n944));
   BUFCHD FE_PHC7064_n1094 (.O(FE_PHN7064_n1094), 
	.I(FE_PHN7357_n1094));
   BUFCHD FE_PHC7063_n1874 (.O(FE_PHN7063_n1874), 
	.I(FE_PHN7345_n1874));
   BUFGHD FE_PHC7062_n2611 (.O(FE_PHN7062_n2611), 
	.I(FE_PHN7335_n2611));
   BUFCHD FE_PHC7061_n1178 (.O(FE_PHN7061_n1178), 
	.I(FE_PHN7324_n1178));
   BUFCHD FE_PHC7060_n1872 (.O(FE_PHN7060_n1872), 
	.I(FE_PHN7329_n1872));
   BUFCHD FE_PHC7059_n4116 (.O(FE_PHN7059_n4116), 
	.I(FE_PHN7340_n4116));
   BUFCHD FE_PHC7058_n2411 (.O(FE_PHN7058_n2411), 
	.I(FE_PHN4800_n2411));
   BUFEHD FE_PHC7057_n4148 (.O(FE_PHN7057_n4148), 
	.I(FE_PHN7322_n4148));
   BUFCHD FE_PHC7056_n1918 (.O(FE_PHN7056_n1918), 
	.I(FE_PHN7359_n1918));
   BUFCHD FE_PHC7055_n964 (.O(FE_PHN7055_n964), 
	.I(FE_PHN7320_n964));
   BUFCHD FE_PHC7054_n2423 (.O(FE_PHN7054_n2423), 
	.I(FE_PHN4881_n2423));
   BUFCKEHD FE_PHC7053_n3932 (.O(FE_PHN7053_n3932), 
	.I(FE_PHN7352_n3932));
   BUFCHD FE_PHC7052_n950 (.O(FE_PHN7052_n950), 
	.I(FE_PHN7326_n950));
   BUFCHD FE_PHC7051_n2594 (.O(FE_PHN7051_n2594), 
	.I(FE_PHN7381_n2594));
   BUFCHD FE_PHC7050_n906 (.O(FE_PHN7050_n906), 
	.I(FE_PHN7321_n906));
   BUFCHD FE_PHC7049_n2137 (.O(FE_PHN7049_n2137), 
	.I(FE_PHN4823_n2137));
   BUFCHD FE_PHC7048_n2138 (.O(FE_PHN7048_n2138), 
	.I(FE_PHN7316_n2138));
   BUFCHD FE_PHC7047_n2149 (.O(FE_PHN7047_n2149), 
	.I(FE_PHN7338_n2149));
   BUFCHD FE_PHC7046_n2618 (.O(FE_PHN7046_n2618), 
	.I(FE_PHN7343_n2618));
   BUFCHD FE_PHC7045_n2124 (.O(FE_PHN7045_n2124), 
	.I(FE_PHN7323_n2124));
   BUFCHD FE_PHC7044_n4142 (.O(FE_PHN7044_n4142), 
	.I(FE_PHN7360_n4142));
   BUFCKKHD FE_PHC7043_n1880 (.O(FE_PHN7043_n1880), 
	.I(FE_PHN7367_n1880));
   BUFCHD FE_PHC7042_n1154 (.O(FE_PHN7042_n1154), 
	.I(FE_PHN7313_n1154));
   BUFCHD FE_PHC7041_n2622 (.O(FE_PHN7041_n2622), 
	.I(FE_PHN7318_n2622));
   BUFCKMHD FE_PHC7040_n953 (.O(FE_PHN7040_n953), 
	.I(FE_PHN7334_n953));
   BUFCHD FE_PHC7039_n2598 (.O(FE_PHN7039_n2598), 
	.I(FE_PHN4438_n2598));
   BUFCKLHD FE_PHC7038_n1922 (.O(FE_PHN7038_n1922), 
	.I(FE_PHN7370_n1922));
   BUFCHD FE_PHC7037_n2602 (.O(FE_PHN7037_n2602), 
	.I(FE_PHN7327_n2602));
   BUFCHD FE_PHC7036_n1919 (.O(FE_PHN7036_n1919), 
	.I(FE_PHN7330_n1919));
   BUFCHD FE_PHC7035_n2576 (.O(FE_PHN7035_n2576), 
	.I(FE_PHN7325_n2576));
   BUFCKEHD FE_PHC7034_n938 (.O(FE_PHN7034_n938), 
	.I(FE_PHN7311_n938));
   BUFCKLHD FE_PHC7033_n4110 (.O(FE_PHN7033_n4110), 
	.I(FE_PHN7351_n4110));
   BUFCHD FE_PHC7032_n2388 (.O(FE_PHN7032_n2388), 
	.I(FE_PHN7348_n2388));
   BUFCHD FE_PHC7031_n1001 (.O(FE_PHN7031_n1001), 
	.I(FE_PHN7310_n1001));
   BUFCHD FE_PHC7030_n2412 (.O(FE_PHN7030_n2412), 
	.I(FE_PHN7332_n2412));
   BUFCHD FE_PHC7029_n4114 (.O(FE_PHN7029_n4114), 
	.I(FE_PHN7314_n4114));
   BUFCHD FE_PHC7028_n2572 (.O(FE_PHN7028_n2572), 
	.I(FE_PHN7317_n2572));
   BUFCHD FE_PHC7027_n2251 (.O(FE_PHN7027_n2251), 
	.I(FE_PHN7312_n2251));
   BUFCHD FE_PHC7026_n2612 (.O(FE_PHN7026_n2612), 
	.I(FE_PHN7315_n2612));
   BUFCHD FE_PHC7025_n844 (.O(FE_PHN7025_n844), 
	.I(FE_PHN4520_n844));
   BUFCKEHD FE_PHC7024_n3131 (.O(FE_PHN7024_n3131), 
	.I(FE_PHN3453_n3131));
   BUFCHD FE_PHC7023_n3924 (.O(FE_PHN7023_n3924), 
	.I(FE_PHN3449_n3924));
   BUFCKEHD FE_PHC7022_n4204 (.O(FE_PHN7022_n4204), 
	.I(FE_PHN4032_n4204));
   BUFCHD FE_PHC7021_n2995 (.O(FE_PHN7021_n2995), 
	.I(n2995));
   BUFCHD FE_PHC7020_n1021 (.O(FE_PHN7020_n1021), 
	.I(FE_PHN3829_n1021));
   BUFCKEHD FE_PHC7019_n3112 (.O(FE_PHN7019_n3112), 
	.I(FE_PHN4045_n3112));
   BUFCHD FE_PHC7018_ram_229__12_ (.O(FE_PHN7018_ram_229__12_), 
	.I(FE_PHN3531_ram_229__12_));
   BUFCHD FE_PHC7017_n882 (.O(FE_PHN7017_n882), 
	.I(FE_PHN3492_n882));
   BUFCHD FE_PHC7016_n2928 (.O(FE_PHN7016_n2928), 
	.I(FE_PHN3718_n2928));
   BUFCHD FE_PHC7015_n1030 (.O(FE_PHN7015_n1030), 
	.I(FE_PHN3820_n1030));
   BUFCHD FE_PHC7014_n3078 (.O(FE_PHN7014_n3078), 
	.I(FE_PHN4177_n3078));
   BUFCHD FE_PHC7013_n2970 (.O(FE_PHN7013_n2970), 
	.I(FE_PHN3867_n2970));
   BUFCHD FE_PHC7012_n4243 (.O(FE_PHN7012_n4243), 
	.I(FE_PHN3268_n4243));
   BUFCKEHD FE_PHC7011_n2980 (.O(FE_PHN7011_n2980), 
	.I(FE_PHN4238_n2980));
   BUFCKEHD FE_PHC7010_n3087 (.O(FE_PHN7010_n3087), 
	.I(FE_PHN3282_n3087));
   BUFCHD FE_PHC7009_n2896 (.O(FE_PHN7009_n2896), 
	.I(FE_PHN4528_n2896));
   BUFCHD FE_PHC7008_n4245 (.O(FE_PHN7008_n4245), 
	.I(FE_PHN4136_n4245));
   BUFCHD FE_PHC7007_n4238 (.O(FE_PHN7007_n4238), 
	.I(FE_PHN3599_n4238));
   BUFCHD FE_PHC7006_n870 (.O(FE_PHN7006_n870), 
	.I(FE_PHN3990_n870));
   BUFCKEHD FE_PHC7005_ram_145__7_ (.O(FE_PHN7005_ram_145__7_), 
	.I(FE_PHN4123_ram_145__7_));
   BUFCHD FE_PHC7004_n4359 (.O(FE_PHN7004_n4359), 
	.I(FE_PHN3581_n4359));
   BUFCHD FE_PHC7003_n4094 (.O(FE_PHN7003_n4094), 
	.I(FE_PHN5611_n4094));
   BUFCHD FE_PHC7002_n4196 (.O(FE_PHN7002_n4196), 
	.I(FE_PHN3396_n4196));
   BUFCHD FE_PHC7001_n4262 (.O(FE_PHN7001_n4262), 
	.I(FE_PHN3521_n4262));
   BUFCHD FE_PHC7000_n3921 (.O(FE_PHN7000_n3921), 
	.I(FE_PHN3710_n3921));
   BUFCKEHD FE_PHC6999_n999 (.O(FE_PHN6999_n999), 
	.I(FE_PHN3877_n999));
   BUFCHD FE_PHC6998_n2906 (.O(FE_PHN6998_n2906), 
	.I(FE_PHN4442_n2906));
   BUFCHD FE_PHC6997_n891 (.O(FE_PHN6997_n891), 
	.I(FE_PHN3971_n891));
   BUFCKEHD FE_PHC6996_n4281 (.O(FE_PHN6996_n4281), 
	.I(FE_PHN3370_n4281));
   BUFCHD FE_PHC6995_n3075 (.O(FE_PHN6995_n3075), 
	.I(FE_PHN3868_n3075));
   BUFCHD FE_PHC6994_n4251 (.O(FE_PHN6994_n4251), 
	.I(FE_PHN4060_n4251));
   BUFCKEHD FE_PHC6993_n3926 (.O(FE_PHN6993_n3926), 
	.I(FE_PHN3724_n3926));
   BUFCHD FE_PHC6992_n3056 (.O(FE_PHN6992_n3056), 
	.I(FE_PHN3648_n3056));
   BUFCHD FE_PHC6991_n4134 (.O(FE_PHN6991_n4134), 
	.I(FE_PHN4398_n4134));
   BUFCHD FE_PHC6990_n3099 (.O(FE_PHN6990_n3099), 
	.I(FE_PHN4108_n3099));
   BUFCHD FE_PHC6989_n2997 (.O(FE_PHN6989_n2997), 
	.I(FE_PHN3736_n2997));
   BUFCHD FE_PHC6988_n969 (.O(FE_PHN6988_n969), 
	.I(FE_PHN3957_n969));
   BUFCHD FE_PHC6987_n3918 (.O(FE_PHN6987_n3918), 
	.I(FE_PHN4555_n3918));
   BUFCHD FE_PHC6986_n1068 (.O(FE_PHN6986_n1068), 
	.I(n1068));
   BUFCHD FE_PHC6985_n3969 (.O(FE_PHN6985_n3969), 
	.I(FE_PHN3289_n3969));
   BUFCHD FE_PHC6984_n3265 (.O(FE_PHN6984_n3265), 
	.I(FE_PHN4135_n3265));
   BUFCKEHD FE_PHC6983_n3940 (.O(FE_PHN6983_n3940), 
	.I(FE_PHN3795_n3940));
   BUFCHD FE_PHC6982_n884 (.O(FE_PHN6982_n884), 
	.I(FE_PHN3318_n884));
   BUFCKEHD FE_PHC6981_n4201 (.O(FE_PHN6981_n4201), 
	.I(n4201));
   BUFCKEHD FE_PHC6980_n951 (.O(FE_PHN6980_n951), 
	.I(FE_PHN4291_n951));
   BUFCHD FE_PHC6979_n890 (.O(FE_PHN6979_n890), 
	.I(FE_PHN3570_n890));
   BUFCHD FE_PHC6978_n4333 (.O(FE_PHN6978_n4333), 
	.I(FE_PHN3936_n4333));
   BUFCHD FE_PHC6977_n3108 (.O(FE_PHN6977_n3108), 
	.I(FE_PHN3386_n3108));
   BUFCKEHD FE_PHC6976_ram_214__13_ (.O(FE_PHN6976_ram_214__13_), 
	.I(FE_PHN4441_ram_214__13_));
   BUFCKEHD FE_PHC6975_n4266 (.O(FE_PHN6975_n4266), 
	.I(FE_PHN3480_n4266));
   BUFCKEHD FE_PHC6974_n1006 (.O(FE_PHN6974_n1006), 
	.I(FE_PHN4336_n1006));
   BUFCHD FE_PHC6973_n2926 (.O(FE_PHN6973_n2926), 
	.I(n2926));
   BUFCHD FE_PHC6972_n4269 (.O(FE_PHN6972_n4269), 
	.I(FE_PHN4171_n4269));
   BUFCKEHD FE_PHC6971_n2994 (.O(FE_PHN6971_n2994), 
	.I(FE_PHN3584_n2994));
   BUFCHD FE_PHC6970_n3098 (.O(FE_PHN6970_n3098), 
	.I(FE_PHN3616_n3098));
   BUFCHD FE_PHC6969_n2897 (.O(FE_PHN6969_n2897), 
	.I(FE_PHN4436_n2897));
   BUFCKEHD FE_PHC6968_n3024 (.O(FE_PHN6968_n3024), 
	.I(FE_PHN4550_n3024));
   BUFCHD FE_PHC6967_n2933 (.O(FE_PHN6967_n2933), 
	.I(FE_PHN3979_n2933));
   BUFCHD FE_PHC6966_n3076 (.O(FE_PHN6966_n3076), 
	.I(FE_PHN3959_n3076));
   BUFCKEHD FE_PHC6965_n3084 (.O(FE_PHN6965_n3084), 
	.I(FE_PHN4098_n3084));
   BUFCKEHD FE_PHC6964_n3958 (.O(FE_PHN6964_n3958), 
	.I(FE_PHN3524_n3958));
   BUFCHD FE_PHC6963_n4271 (.O(FE_PHN6963_n4271), 
	.I(FE_PHN3652_n4271));
   BUFCKEHD FE_PHC6962_n4339 (.O(FE_PHN6962_n4339), 
	.I(FE_PHN4066_n4339));
   BUFCHD FE_PHC6961_n3994 (.O(FE_PHN6961_n3994), 
	.I(FE_PHN3819_n3994));
   BUFCHD FE_PHC6960_n1110 (.O(FE_PHN6960_n1110), 
	.I(FE_PHN5172_n1110));
   BUFCHD FE_PHC6959_n2934 (.O(FE_PHN6959_n2934), 
	.I(FE_PHN4389_n2934));
   BUFCHD FE_PHC6958_n892 (.O(FE_PHN6958_n892), 
	.I(FE_PHN3997_n892));
   BUFCKEHD FE_PHC6957_n4355 (.O(FE_PHN6957_n4355), 
	.I(FE_PHN3354_n4355));
   BUFCHD FE_PHC6956_n4003 (.O(FE_PHN6956_n4003), 
	.I(FE_PHN3294_n4003));
   BUFCKEHD FE_PHC6955_n2978 (.O(FE_PHN6955_n2978), 
	.I(FE_PHN3577_n2978));
   BUFCHD FE_PHC6954_n2946 (.O(FE_PHN6954_n2946), 
	.I(FE_PHN3951_n2946));
   BUFCHD FE_PHC6953_n4362 (.O(FE_PHN6953_n4362), 
	.I(FE_PHN3797_n4362));
   BUFCHD FE_PHC6952_n3103 (.O(FE_PHN6952_n3103), 
	.I(FE_PHN3434_n3103));
   BUFCHD FE_PHC6951_n3931 (.O(FE_PHN6951_n3931), 
	.I(FE_PHN3234_n3931));
   BUFCKEHD FE_PHC6950_n4410 (.O(FE_PHN6950_n4410), 
	.I(FE_PHN3914_n4410));
   BUFCKEHD FE_PHC6949_n4361 (.O(FE_PHN6949_n4361), 
	.I(FE_PHN3970_n4361));
   BUFCKEHD FE_PHC6948_n2987 (.O(FE_PHN6948_n2987), 
	.I(FE_PHN3556_n2987));
   BUFCHD FE_PHC6947_n4233 (.O(FE_PHN6947_n4233), 
	.I(FE_PHN3508_n4233));
   BUFCHD FE_PHC6946_n4387 (.O(FE_PHN6946_n4387), 
	.I(FE_PHN3943_n4387));
   BUFCHD FE_PHC6945_ram_153__11_ (.O(FE_PHN6945_ram_153__11_), 
	.I(FE_PHN3690_ram_153__11_));
   BUFCHD FE_PHC6944_n2399 (.O(FE_PHN6944_n2399), 
	.I(FE_PHN4345_n2399));
   BUFCKEHD FE_PHC6943_n3079 (.O(FE_PHN6943_n3079), 
	.I(FE_PHN4349_n3079));
   BUFCHD FE_PHC6942_n919 (.O(FE_PHN6942_n919), 
	.I(FE_PHN3757_n919));
   BUFCKEHD FE_PHC6941_n1020 (.O(FE_PHN6941_n1020), 
	.I(FE_PHN4595_n1020));
   BUFCHD FE_PHC6940_n2413 (.O(FE_PHN6940_n2413), 
	.I(n2413));
   BUFCHD FE_PHC6939_n957 (.O(FE_PHN6939_n957), 
	.I(FE_PHN4435_n957));
   BUFCHD FE_PHC6938_n2992 (.O(FE_PHN6938_n2992), 
	.I(FE_PHN4563_n2992));
   BUFCKEHD FE_PHC6937_n3952 (.O(FE_PHN6937_n3952), 
	.I(FE_PHN3517_n3952));
   BUFCHD FE_PHC6936_n3910 (.O(FE_PHN6936_n3910), 
	.I(FE_PHN3477_n3910));
   BUFCHD FE_PHC6935_n1093 (.O(FE_PHN6935_n1093), 
	.I(FE_PHN4053_n1093));
   BUFCKEHD FE_PHC6934_n4076 (.O(FE_PHN6934_n4076), 
	.I(FE_PHN3781_n4076));
   BUFCKEHD FE_PHC6933_ram_221__1_ (.O(FE_PHN6933_ram_221__1_), 
	.I(FE_PHN6248_ram_221__1_));
   BUFCKEHD FE_PHC6932_n4222 (.O(FE_PHN6932_n4222), 
	.I(FE_PHN3747_n4222));
   BUFCHD FE_PHC6931_n2916 (.O(FE_PHN6931_n2916), 
	.I(FE_PHN3852_n2916));
   BUFCKEHD FE_PHC6930_n3915 (.O(FE_PHN6930_n3915), 
	.I(FE_PHN4113_n3915));
   BUFCKEHD FE_PHC6929_n4295 (.O(FE_PHN6929_n4295), 
	.I(FE_PHN3539_n4295));
   BUFCKEHD FE_PHC6928_n1087 (.O(FE_PHN6928_n1087), 
	.I(FE_PHN4216_n1087));
   BUFCKEHD FE_PHC6927_n4169 (.O(FE_PHN6927_n4169), 
	.I(FE_PHN3543_n4169));
   BUFCHD FE_PHC6926_n4291 (.O(FE_PHN6926_n4291), 
	.I(FE_PHN3808_n4291));
   BUFCHD FE_PHC6925_n4202 (.O(FE_PHN6925_n4202), 
	.I(FE_PHN3988_n4202));
   BUFCKEHD FE_PHC6924_n3956 (.O(FE_PHN6924_n3956), 
	.I(FE_PHN3788_n3956));
   BUFCHD FE_PHC6923_n3060 (.O(FE_PHN6923_n3060), 
	.I(FE_PHN4303_n3060));
   BUFCHD FE_PHC6922_n3976 (.O(FE_PHN6922_n3976), 
	.I(FE_PHN3466_n3976));
   BUFCHD FE_PHC6921_n3996 (.O(FE_PHN6921_n3996), 
	.I(FE_PHN4413_n3996));
   BUFCKEHD FE_PHC6920_n3947 (.O(FE_PHN6920_n3947), 
	.I(FE_PHN4031_n3947));
   BUFCKEHD FE_PHC6919_n848 (.O(FE_PHN6919_n848), 
	.I(FE_PHN3376_n848));
   BUFCKEHD FE_PHC6918_n4183 (.O(FE_PHN6918_n4183), 
	.I(FE_PHN4558_n4183));
   BUFCKEHD FE_PHC6917_n2621 (.O(FE_PHN6917_n2621), 
	.I(FE_PHN3962_n2621));
   BUFCHD FE_PHC6916_n4111 (.O(FE_PHN6916_n4111), 
	.I(FE_PHN3818_n4111));
   BUFCHD FE_PHC6915_n4021 (.O(FE_PHN6915_n4021), 
	.I(FE_PHN3248_n4021));
   BUFCKEHD FE_PHC6914_n936 (.O(FE_PHN6914_n936), 
	.I(FE_PHN4468_n936));
   BUFCKEHD FE_PHC6913_ram_144__8_ (.O(FE_PHN6913_ram_144__8_), 
	.I(FE_PHN3641_ram_144__8_));
   BUFCHD FE_PHC6912_n3954 (.O(FE_PHN6912_n3954), 
	.I(FE_PHN4016_n3954));
   BUFCKEHD FE_PHC6911_n846 (.O(FE_PHN6911_n846), 
	.I(FE_PHN5173_n846));
   BUFCKEHD FE_PHC6910_n994 (.O(FE_PHN6910_n994), 
	.I(FE_PHN4315_n994));
   BUFCKEHD FE_PHC6909_n2936 (.O(FE_PHN6909_n2936), 
	.I(FE_PHN3257_n2936));
   BUFCHD FE_PHC6908_n4371 (.O(FE_PHN6908_n4371), 
	.I(FE_PHN3582_n4371));
   BUFCHD FE_PHC6907_n3936 (.O(FE_PHN6907_n3936), 
	.I(FE_PHN3429_n3936));
   BUFCHD FE_PHC6906_n2735 (.O(FE_PHN6906_n2735), 
	.I(FE_PHN3900_n2735));
   BUFCHD FE_PHC6905_n1899 (.O(FE_PHN6905_n1899), 
	.I(FE_PHN3864_n1899));
   BUFCKEHD FE_PHC6904_n4311 (.O(FE_PHN6904_n4311), 
	.I(FE_PHN3332_n4311));
   BUFCHD FE_PHC6903_n3984 (.O(FE_PHN6903_n3984), 
	.I(FE_PHN3693_n3984));
   BUFCHD FE_PHC6902_n876 (.O(FE_PHN6902_n876), 
	.I(FE_PHN4103_n876));
   BUFCHD FE_PHC6901_n2437 (.O(FE_PHN6901_n2437), 
	.I(FE_PHN3809_n2437));
   BUFCKEHD FE_PHC6900_n4239 (.O(FE_PHN6900_n4239), 
	.I(FE_PHN4153_n4239));
   BUFCKEHD FE_PHC6899_n872 (.O(FE_PHN6899_n872), 
	.I(FE_PHN3732_n872));
   BUFCHD FE_PHC6898_n3951 (.O(FE_PHN6898_n3951), 
	.I(FE_PHN3871_n3951));
   BUFCHD FE_PHC6897_n3959 (.O(FE_PHN6897_n3959), 
	.I(FE_PHN4180_n3959));
   BUFCHD FE_PHC6896_n3998 (.O(FE_PHN6896_n3998), 
	.I(FE_PHN4013_n3998));
   BUFCHD FE_PHC6895_n840 (.O(FE_PHN6895_n840), 
	.I(FE_PHN3857_n840));
   BUFCHD FE_PHC6894_n4252 (.O(FE_PHN6894_n4252), 
	.I(FE_PHN3239_n4252));
   BUFCHD FE_PHC6893_n988 (.O(FE_PHN6893_n988), 
	.I(FE_PHN5208_n988));
   BUFCHD FE_PHC6892_n961 (.O(FE_PHN6892_n961), 
	.I(FE_PHN4006_n961));
   BUFCHD FE_PHC6891_n4172 (.O(FE_PHN6891_n4172), 
	.I(FE_PHN3755_n4172));
   BUFCHD FE_PHC6890_n1106 (.O(FE_PHN6890_n1106), 
	.I(FE_PHN4636_n1106));
   BUFCHD FE_PHC6889_n3948 (.O(FE_PHN6889_n3948), 
	.I(FE_PHN3500_n3948));
   BUFCHD FE_PHC6888_n2158 (.O(FE_PHN6888_n2158), 
	.I(n2158));
   BUFCHD FE_PHC6887_n3027 (.O(FE_PHN6887_n3027), 
	.I(FE_PHN3583_n3027));
   BUFCKEHD FE_PHC6886_n4033 (.O(FE_PHN6886_n4033), 
	.I(FE_PHN3263_n4033));
   BUFCHD FE_PHC6885_n958 (.O(FE_PHN6885_n958), 
	.I(FE_PHN3436_n958));
   BUFCHD FE_PHC6884_n2967 (.O(FE_PHN6884_n2967), 
	.I(FE_PHN3859_n2967));
   BUFCKEHD FE_PHC6883_n4324 (.O(FE_PHN6883_n4324), 
	.I(FE_PHN3233_n4324));
   BUFCHD FE_PHC6882_n4017 (.O(FE_PHN6882_n4017), 
	.I(FE_PHN3397_n4017));
   BUFCHD FE_PHC6881_n2374 (.O(FE_PHN6881_n2374), 
	.I(FE_PHN5016_n2374));
   BUFCKEHD FE_PHC6880_n4028 (.O(FE_PHN6880_n4028), 
	.I(FE_PHN3361_n4028));
   BUFCKEHD FE_PHC6879_n3972 (.O(FE_PHN6879_n3972), 
	.I(FE_PHN4197_n3972));
   BUFCKEHD FE_PHC6878_n3914 (.O(FE_PHN6878_n3914), 
	.I(FE_PHN6187_n3914));
   BUFCHD FE_PHC6877_n1056 (.O(FE_PHN6877_n1056), 
	.I(FE_PHN3525_n1056));
   BUFCHD FE_PHC6876_n3063 (.O(FE_PHN6876_n3063), 
	.I(FE_PHN3290_n3063));
   BUFCHD FE_PHC6875_n3025 (.O(FE_PHN6875_n3025), 
	.I(FE_PHN4381_n3025));
   BUFCHD FE_PHC6874_n4005 (.O(FE_PHN6874_n4005), 
	.I(FE_PHN3412_n4005));
   BUFCHD FE_PHC6873_n1066 (.O(FE_PHN6873_n1066), 
	.I(FE_PHN3563_n1066));
   BUFCKEHD FE_PHC6872_n3257 (.O(FE_PHN6872_n3257), 
	.I(FE_PHN3985_n3257));
   BUFCKEHD FE_PHC6871_n4185 (.O(FE_PHN6871_n4185), 
	.I(FE_PHN3934_n4185));
   BUFCKEHD FE_PHC6870_n4166 (.O(FE_PHN6870_n4166), 
	.I(FE_PHN3378_n4166));
   BUFCHD FE_PHC6869_n4188 (.O(FE_PHN6869_n4188), 
	.I(FE_PHN3589_n4188));
   BUFCKEHD FE_PHC6868_n839 (.O(FE_PHN6868_n839), 
	.I(FE_PHN3660_n839));
   BUFCHD FE_PHC6867_n4327 (.O(FE_PHN6867_n4327), 
	.I(FE_PHN3458_n4327));
   BUFCHD FE_PHC6866_n851 (.O(FE_PHN6866_n851), 
	.I(FE_PHN3903_n851));
   BUFCHD FE_PHC6865_n3937 (.O(FE_PHN6865_n3937), 
	.I(FE_PHN3313_n3937));
   BUFCHD FE_PHC6864_n989 (.O(FE_PHN6864_n989), 
	.I(FE_PHN4225_n989));
   BUFCKEHD FE_PHC6863_n1078 (.O(FE_PHN6863_n1078), 
	.I(FE_PHN4148_n1078));
   BUFCHD FE_PHC6862_ram_133__9_ (.O(FE_PHN6862_ram_133__9_), 
	.I(FE_PHN4511_ram_133__9_));
   BUFCHD FE_PHC6861_n3987 (.O(FE_PHN6861_n3987), 
	.I(FE_PHN4219_n3987));
   BUFCHD FE_PHC6860_n2943 (.O(FE_PHN6860_n2943), 
	.I(FE_PHN3826_n2943));
   BUFCHD FE_PHC6859_n2998 (.O(FE_PHN6859_n2998), 
	.I(FE_PHN3666_n2998));
   BUFCKEHD FE_PHC6858_n902 (.O(FE_PHN6858_n902), 
	.I(FE_PHN6140_n902));
   BUFCHD FE_PHC6857_n4211 (.O(FE_PHN6857_n4211), 
	.I(FE_PHN3538_n4211));
   BUFCHD FE_PHC6856_n4377 (.O(FE_PHN6856_n4377), 
	.I(FE_PHN3304_n4377));
   BUFCHD FE_PHC6855_n3943 (.O(FE_PHN6855_n3943), 
	.I(FE_PHN4143_n3943));
   BUFCHD FE_PHC6854_n4226 (.O(FE_PHN6854_n4226), 
	.I(FE_PHN3550_n4226));
   BUFCHD FE_PHC6853_n855 (.O(FE_PHN6853_n855), 
	.I(FE_PHN3276_n855));
   BUFCHD FE_PHC6852_n1051 (.O(FE_PHN6852_n1051), 
	.I(FE_PHN5068_n1051));
   BUFCHD FE_PHC6851_n3029 (.O(FE_PHN6851_n3029), 
	.I(FE_PHN4521_n3029));
   BUFCHD FE_PHC6850_n3930 (.O(FE_PHN6850_n3930), 
	.I(FE_PHN3462_n3930));
   BUFCHD FE_PHC6849_n2971 (.O(FE_PHN6849_n2971), 
	.I(FE_PHN3651_n2971));
   BUFCHD FE_PHC6848_n852 (.O(FE_PHN6848_n852), 
	.I(FE_PHN3668_n852));
   BUFCHD FE_PHC6847_n3116 (.O(FE_PHN6847_n3116), 
	.I(FE_PHN4052_n3116));
   BUFCKEHD FE_PHC6846_n857 (.O(FE_PHN6846_n857), 
	.I(FE_PHN3529_n857));
   BUFCKEHD FE_PHC6845_n3963 (.O(FE_PHN6845_n3963), 
	.I(FE_PHN3815_n3963));
   BUFCHD FE_PHC6844_n1069 (.O(FE_PHN6844_n1069), 
	.I(FE_PHN3673_n1069));
   BUFCKEHD FE_PHC6843_n2258 (.O(FE_PHN6843_n2258), 
	.I(n2258));
   BUFCHD FE_PHC6842_n4217 (.O(FE_PHN6842_n4217), 
	.I(FE_PHN3902_n4217));
   BUFCHD FE_PHC6841_n3043 (.O(FE_PHN6841_n3043), 
	.I(FE_PHN4204_n3043));
   BUFCHD FE_PHC6840_n4323 (.O(FE_PHN6840_n4323), 
	.I(FE_PHN3503_n4323));
   BUFCKEHD FE_PHC6839_n2396 (.O(FE_PHN6839_n2396), 
	.I(n2396));
   BUFCHD FE_PHC6838_n2930 (.O(FE_PHN6838_n2930), 
	.I(FE_PHN3348_n2930));
   BUFCHD FE_PHC6837_n3207 (.O(FE_PHN6837_n3207), 
	.I(FE_PHN3908_n3207));
   BUFCKEHD FE_PHC6836_n2433 (.O(FE_PHN6836_n2433), 
	.I(FE_PHN3400_n2433));
   BUFCHD FE_PHC6835_n3052 (.O(FE_PHN6835_n3052), 
	.I(n3052));
   BUFCHD FE_PHC6834_n887 (.O(FE_PHN6834_n887), 
	.I(FE_PHN6045_n887));
   BUFCHD FE_PHC6833_n945 (.O(FE_PHN6833_n945), 
	.I(FE_PHN3892_n945));
   BUFCHD FE_PHC6832_n1896 (.O(FE_PHN6832_n1896), 
	.I(FE_PHN3814_n1896));
   BUFCHD FE_PHC6831_n965 (.O(FE_PHN6831_n965), 
	.I(FE_PHN3789_n965));
   BUFCKEHD FE_PHC6830_n2722 (.O(FE_PHN6830_n2722), 
	.I(FE_PHN3983_n2722));
   BUFCHD FE_PHC6829_n941 (.O(FE_PHN6829_n941), 
	.I(FE_PHN3708_n941));
   BUFCHD FE_PHC6828_n2127 (.O(FE_PHN6828_n2127), 
	.I(n2127));
   BUFCHD FE_PHC6827_n1034 (.O(FE_PHN6827_n1034), 
	.I(FE_PHN4445_n1034));
   BUFCHD FE_PHC6826_n2623 (.O(FE_PHN6826_n2623), 
	.I(FE_PHN3969_n2623));
   BUFCHD FE_PHC6825_n858 (.O(FE_PHN6825_n858), 
	.I(FE_PHN3311_n858));
   BUFCHD FE_PHC6824_n4220 (.O(FE_PHN6824_n4220), 
	.I(FE_PHN3513_n4220));
   BUFCHD FE_PHC6823_n3927 (.O(FE_PHN6823_n3927), 
	.I(FE_PHN4375_n3927));
   BUFCKEHD FE_PHC6822_n866 (.O(FE_PHN6822_n866), 
	.I(FE_PHN4124_n866));
   BUFCHD FE_PHC6821_n889 (.O(FE_PHN6821_n889), 
	.I(FE_PHN4590_n889));
   BUFCHD FE_PHC6820_n4393 (.O(FE_PHN6820_n4393), 
	.I(FE_PHN3325_n4393));
   BUFCHD FE_PHC6819_n4278 (.O(FE_PHN6819_n4278), 
	.I(FE_PHN3459_n4278));
   BUFCHD FE_PHC6818_n4036 (.O(FE_PHN6818_n4036), 
	.I(FE_PHN3952_n4036));
   BUFCKEHD FE_PHC6817_n1037 (.O(FE_PHN6817_n1037), 
	.I(FE_PHN3816_n1037));
   BUFCHD FE_PHC6816_n2932 (.O(FE_PHN6816_n2932), 
	.I(FE_PHN4247_n2932));
   BUFCHD FE_PHC6815_n920 (.O(FE_PHN6815_n920), 
	.I(FE_PHN4232_n920));
   BUFCHD FE_PHC6814_n4307 (.O(FE_PHN6814_n4307), 
	.I(FE_PHN3349_n4307));
   BUFCHD FE_PHC6813_n4029 (.O(FE_PHN6813_n4029), 
	.I(FE_PHN3402_n4029));
   BUFCHD FE_PHC6812_n864 (.O(FE_PHN6812_n864), 
	.I(FE_PHN4248_n864));
   BUFCHD FE_PHC6811_n2754 (.O(FE_PHN6811_n2754), 
	.I(FE_PHN4307_n2754));
   BUFCHD FE_PHC6810_n3988 (.O(FE_PHN6810_n3988), 
	.I(FE_PHN3314_n3988));
   BUFCHD FE_PHC6809_n3023 (.O(FE_PHN6809_n3023), 
	.I(FE_PHN4167_n3023));
   BUFCHD FE_PHC6808_n4195 (.O(FE_PHN6808_n4195), 
	.I(FE_PHN3277_n4195));
   BUFCHD FE_PHC6807_n972 (.O(FE_PHN6807_n972), 
	.I(FE_PHN3723_n972));
   BUFCHD FE_PHC6806_n878 (.O(FE_PHN6806_n878), 
	.I(FE_PHN3528_n878));
   BUFCKEHD FE_PHC6805_n856 (.O(FE_PHN6805_n856), 
	.I(FE_PHN4038_n856));
   BUFCHD FE_PHC6804_n2430 (.O(FE_PHN6804_n2430), 
	.I(FE_PHN3692_n2430));
   BUFCHD FE_PHC6803_n4299 (.O(FE_PHN6803_n4299), 
	.I(FE_PHN3598_n4299));
   BUFCHD FE_PHC6802_n3073 (.O(FE_PHN6802_n3073), 
	.I(FE_PHN3618_n3073));
   BUFCHD FE_PHC6801_n894 (.O(FE_PHN6801_n894), 
	.I(FE_PHN4450_n894));
   BUFCHD FE_PHC6800_n2141 (.O(FE_PHN6800_n2141), 
	.I(n2141));
   BUFCHD FE_PHC6799_n3916 (.O(FE_PHN6799_n3916), 
	.I(FE_PHN3801_n3916));
   BUFCKEHD FE_PHC6798_n4014 (.O(FE_PHN6798_n4014), 
	.I(FE_PHN4140_n4014));
   BUFCHD FE_PHC6797_n913 (.O(FE_PHN6797_n913), 
	.I(FE_PHN3846_n913));
   BUFCHD FE_PHC6796_n3055 (.O(FE_PHN6796_n3055), 
	.I(FE_PHN3631_n3055));
   BUFCHD FE_PHC6795_n861 (.O(FE_PHN6795_n861), 
	.I(FE_PHN3441_n861));
   BUFCHD FE_PHC6794_n943 (.O(FE_PHN6794_n943), 
	.I(FE_PHN5962_n943));
   BUFCHD FE_PHC6793_n4340 (.O(FE_PHN6793_n4340), 
	.I(FE_PHN4114_n4340));
   BUFCHD FE_PHC6792_n3071 (.O(FE_PHN6792_n3071), 
	.I(FE_PHN3407_n3071));
   BUFCHD FE_PHC6791_n929 (.O(FE_PHN6791_n929), 
	.I(FE_PHN3509_n929));
   BUFCHD FE_PHC6790_n2900 (.O(FE_PHN6790_n2900), 
	.I(FE_PHN3878_n2900));
   BUFCHD FE_PHC6789_n1079 (.O(FE_PHN6789_n1079), 
	.I(FE_PHN4342_n1079));
   BUFCHD FE_PHC6788_n4232 (.O(FE_PHN6788_n4232), 
	.I(FE_PHN3705_n4232));
   BUFCHD FE_PHC6787_n4209 (.O(FE_PHN6787_n4209), 
	.I(FE_PHN3834_n4209));
   BUFDHD FE_PHC6786_n1022 (.O(FE_PHN6786_n1022), 
	.I(FE_PHN4373_n1022));
   BUFCHD FE_PHC6785_n2178 (.O(FE_PHN6785_n2178), 
	.I(FE_PHN4058_n2178));
   BUFCHD FE_PHC6784_n4225 (.O(FE_PHN6784_n4225), 
	.I(FE_PHN4163_n4225));
   BUFCHD FE_PHC6783_n935 (.O(FE_PHN6783_n935), 
	.I(FE_PHN3573_n935));
   BUFCKEHD FE_PHC6782_n4001 (.O(FE_PHN6782_n4001), 
	.I(FE_PHN3327_n4001));
   BUFCKEHD FE_PHC6781_n4277 (.O(FE_PHN6781_n4277), 
	.I(FE_PHN3794_n4277));
   BUFCHD FE_PHC6780_n842 (.O(FE_PHN6780_n842), 
	.I(FE_PHN3664_n842));
   BUFCHD FE_PHC6779_n2927 (.O(FE_PHN6779_n2927), 
	.I(FE_PHN3554_n2927));
   BUFCHD FE_PHC6778_n925 (.O(FE_PHN6778_n925), 
	.I(FE_PHN3709_n925));
   BUFCHD FE_PHC6777_n2400 (.O(FE_PHN6777_n2400), 
	.I(FE_PHN4112_n2400));
   BUFCHD FE_PHC6776_n910 (.O(FE_PHN6776_n910), 
	.I(FE_PHN3790_n910));
   BUFCHD FE_PHC6775_n4240 (.O(FE_PHN6775_n4240), 
	.I(FE_PHN3657_n4240));
   BUFCKEHD FE_PHC6774_n2383 (.O(FE_PHN6774_n2383), 
	.I(FE_PHN4304_n2383));
   BUFCHD FE_PHC6773_n3992 (.O(FE_PHN6773_n3992), 
	.I(FE_PHN3578_n3992));
   BUFCKEHD FE_PHC6772_n4203 (.O(FE_PHN6772_n4203), 
	.I(n4203));
   BUFCHD FE_PHC6771_n1038 (.O(FE_PHN6771_n1038), 
	.I(FE_PHN4305_n1038));
   BUFCHD FE_PHC6770_n4000 (.O(FE_PHN6770_n4000), 
	.I(FE_PHN4207_n4000));
   BUFCKEHD FE_PHC6769_n4350 (.O(FE_PHN6769_n4350), 
	.I(FE_PHN3491_n4350));
   BUFCHD FE_PHC6768_n4194 (.O(FE_PHN6768_n4194), 
	.I(FE_PHN3317_n4194));
   BUFCHD FE_PHC6767_n4164 (.O(FE_PHN6767_n4164), 
	.I(FE_PHN3382_n4164));
   BUFCHD FE_PHC6766_n911 (.O(FE_PHN6766_n911), 
	.I(FE_PHN3595_n911));
   BUFCHD FE_PHC6765_n2405 (.O(FE_PHN6765_n2405), 
	.I(FE_PHN3701_n2405));
   BUFCHD FE_PHC6764_n3258 (.O(FE_PHN6764_n3258), 
	.I(FE_PHN3515_n3258));
   BUFCHD FE_PHC6763_n2945 (.O(FE_PHN6763_n2945), 
	.I(FE_PHN3929_n2945));
   BUFCHD FE_PHC6762_n4174 (.O(FE_PHN6762_n4174), 
	.I(FE_PHN7298_n4174));
   BUFCHD FE_PHC6761_n3129 (.O(FE_PHN6761_n3129), 
	.I(FE_PHN7455_n3129));
   BUFCHD FE_PHC6760_n3219 (.O(FE_PHN6760_n3219), 
	.I(FE_PHN4559_n3219));
   BUFCHD FE_PHC6759_n1920 (.O(FE_PHN6759_n1920), 
	.I(FE_PHN3717_n1920));
   BUFCHD FE_PHC6758_n2389 (.O(FE_PHN6758_n2389), 
	.I(FE_PHN3552_n2389));
   BUFCHD FE_PHC6757_n959 (.O(FE_PHN6757_n959), 
	.I(FE_PHN4235_n959));
   BUFCHD FE_PHC6756_n2564 (.O(FE_PHN6756_n2564), 
	.I(FE_PHN7306_n2564));
   BUFCHD FE_PHC6755_n3028 (.O(FE_PHN6755_n3028), 
	.I(FE_PHN7291_n3028));
   BUFCHD FE_PHC6754_n2420 (.O(FE_PHN6754_n2420), 
	.I(FE_PHN3639_n2420));
   BUFCKEHD FE_PHC6753_n928 (.O(FE_PHN6753_n928), 
	.I(FE_PHN7304_n928));
   BUFCHD FE_PHC6752_n905 (.O(FE_PHN6752_n905), 
	.I(FE_PHN7303_n905));
   BUFCHD FE_PHC6751_n3077 (.O(FE_PHN6751_n3077), 
	.I(FE_PHN3768_n3077));
   BUFCHD FE_PHC6750_n2385 (.O(FE_PHN6750_n2385), 
	.I(FE_PHN5234_n2385));
   BUFCHD FE_PHC6749_n4178 (.O(FE_PHN6749_n4178), 
	.I(FE_PHN5367_n4178));
   BUFCHD FE_PHC6748_n1014 (.O(FE_PHN6748_n1014), 
	.I(FE_PHN7288_n1014));
   BUFCHD FE_PHC6747_n4049 (.O(FE_PHN6747_n4049), 
	.I(FE_PHN3721_n4049));
   BUFCHD FE_PHC6746_n1870 (.O(FE_PHN6746_n1870), 
	.I(FE_PHN3551_n1870));
   BUFCHD FE_PHC6745_n1017 (.O(FE_PHN6745_n1017), 
	.I(FE_PHN7290_n1017));
   BUFCHD FE_PHC6744_n3072 (.O(FE_PHN6744_n3072), 
	.I(FE_PHN7308_n3072));
   BUFCHD FE_PHC6743_n4248 (.O(FE_PHN6743_n4248), 
	.I(FE_PHN3965_n4248));
   BUFCHD FE_PHC6742_n4214 (.O(FE_PHN6742_n4214), 
	.I(FE_PHN4145_n4214));
   BUFCHD FE_PHC6741_n2574 (.O(FE_PHN6741_n2574), 
	.I(FE_PHN7299_n2574));
   BUFCHD FE_PHC6740_n4334 (.O(FE_PHN6740_n4334), 
	.I(FE_PHN3610_n4334));
   BUFCHD FE_PHC6739_n2431 (.O(FE_PHN6739_n2431), 
	.I(FE_PHN3567_n2431));
   BUFCHD FE_PHC6738_n1902 (.O(FE_PHN6738_n1902), 
	.I(FE_PHN3764_n1902));
   BUFCHD FE_PHC6737_n3919 (.O(FE_PHN6737_n3919), 
	.I(FE_PHN7302_n3919));
   BUFCHD FE_PHC6736_n2415 (.O(FE_PHN6736_n2415), 
	.I(FE_PHN3782_n2415));
   BUFCHD FE_PHC6735_n4046 (.O(FE_PHN6735_n4046), 
	.I(FE_PHN7309_n4046));
   BUFCHD FE_PHC6734_n4255 (.O(FE_PHN6734_n4255), 
	.I(FE_PHN4540_n4255));
   BUFCHD FE_PHC6733_n3263 (.O(FE_PHN6733_n3263), 
	.I(FE_PHN3586_n3263));
   BUFCHD FE_PHC6732_n4343 (.O(FE_PHN6732_n4343), 
	.I(FE_PHN4023_n4343));
   BUFCHD FE_PHC6731_n3964 (.O(FE_PHN6731_n3964), 
	.I(FE_PHN7287_n3964));
   BUFCKEHD FE_PHC6730_n975 (.O(FE_PHN6730_n975), 
	.I(FE_PHN7297_n975));
   BUFCHD FE_PHC6729_n1905 (.O(FE_PHN6729_n1905), 
	.I(FE_PHN3752_n1905));
   BUFCKEHD FE_PHC6728_n4215 (.O(FE_PHN6728_n4215), 
	.I(FE_PHN7301_n4215));
   BUFCHD FE_PHC6727_n4180 (.O(FE_PHN6727_n4180), 
	.I(FE_PHN7305_n4180));
   BUFCHD FE_PHC6726_n946 (.O(FE_PHN6726_n946), 
	.I(FE_PHN4164_n946));
   BUFCHD FE_PHC6725_n2408 (.O(FE_PHN6725_n2408), 
	.I(FE_PHN3874_n2408));
   BUFCHD FE_PHC6724_n2580 (.O(FE_PHN6724_n2580), 
	.I(FE_PHN7292_n2580));
   BUFCHD FE_PHC6723_n3040 (.O(FE_PHN6723_n3040), 
	.I(n3040));
   BUFCKGHD FE_PHC6722_n2599 (.O(FE_PHN6722_n2599), 
	.I(FE_PHN7296_n2599));
   BUFCHD FE_PHC6721_n948 (.O(FE_PHN6721_n948), 
	.I(FE_PHN7294_n948));
   BUFCHD FE_PHC6720_n954 (.O(FE_PHN6720_n954), 
	.I(FE_PHN3899_n954));
   BUFCHD FE_PHC6719_n1013 (.O(FE_PHN6719_n1013), 
	.I(FE_PHN7285_n1013));
   BUFCHD FE_PHC6718_n4219 (.O(FE_PHN6718_n4219), 
	.I(FE_PHN7300_n4219));
   BUFCKEHD FE_PHC6717_n2964 (.O(FE_PHN6717_n2964), 
	.I(n2964));
   BUFCHD FE_PHC6716_n4229 (.O(FE_PHN6716_n4229), 
	.I(FE_PHN7289_n4229));
   BUFCHD FE_PHC6715_n1873 (.O(FE_PHN6715_n1873), 
	.I(FE_PHN3763_n1873));
   BUFCKEHD FE_PHC6714_n1082 (.O(FE_PHN6714_n1082), 
	.I(FE_PHN7295_n1082));
   BUFCHD FE_PHC6713_n974 (.O(FE_PHN6713_n974), 
	.I(FE_PHN7286_n974));
   BUFCHD FE_PHC6712_n3068 (.O(FE_PHN6712_n3068), 
	.I(FE_PHN7281_n3068));
   BUFCHD FE_PHC6711_n2133 (.O(FE_PHN6711_n2133), 
	.I(FE_PHN7277_n2133));
   BUFCKLHD FE_PHC6710_n2610 (.O(FE_PHN6710_n2610), 
	.I(n2610));
   BUFCHD FE_PHC6709_n2180 (.O(FE_PHN6709_n2180), 
	.I(FE_PHN7388_n2180));
   BUFEHD FE_PHC6708_n2166 (.O(FE_PHN6708_n2166), 
	.I(FE_PHN7221_n2166));
   BUFCHD FE_PHC6707_n2167 (.O(FE_PHN6707_n2167), 
	.I(FE_PHN7234_n2167));
   BUFCHD FE_PHC6706_n2890 (.O(FE_PHN6706_n2890), 
	.I(FE_PHN7390_n2890));
   BUFCHD FE_PHC6705_n4409 (.O(FE_PHN6705_n4409), 
	.I(FE_PHN7282_n4409));
   BUFCHD FE_PHC6704_n2887 (.O(FE_PHN6704_n2887), 
	.I(FE_PHN7430_n2887));
   BUFMHD FE_PHC6703_n2126 (.O(FE_PHN6703_n2126), 
	.I(FE_PHN7268_n2126));
   BUFCHD FE_PHC6702_n4013 (.O(FE_PHN6702_n4013), 
	.I(FE_PHN7278_n4013));
   BUFCHD FE_PHC6701_n4137 (.O(FE_PHN6701_n4137), 
	.I(FE_PHN7242_n4137));
   BUFCHD FE_PHC6700_n3953 (.O(FE_PHN6700_n3953), 
	.I(FE_PHN7262_n3953));
   BUFCHD FE_PHC6699_n2120 (.O(FE_PHN6699_n2120), 
	.I(FE_PHN7248_n2120));
   BUFCHD FE_PHC6698_n3230 (.O(FE_PHN6698_n3230), 
	.I(FE_PHN7238_n3230));
   BUFCHD FE_PHC6697_n2614 (.O(FE_PHN6697_n2614), 
	.I(FE_PHN7217_n2614));
   BUFMHD FE_PHC6696_n2570 (.O(FE_PHN6696_n2570), 
	.I(FE_PHN7261_n2570));
   BUFCHD FE_PHC6695_n2179 (.O(FE_PHN6695_n2179), 
	.I(FE_PHN7259_n2179));
   BUFCHD FE_PHC6694_n2175 (.O(FE_PHN6694_n2175), 
	.I(FE_PHN7255_n2175));
   BUFCKIHD FE_PHC6693_n2154 (.O(FE_PHN6693_n2154), 
	.I(FE_PHN7231_n2154));
   BUFCHD FE_PHC6692_n2972 (.O(FE_PHN6692_n2972), 
	.I(FE_PHN7283_n2972));
   BUFLHD FE_PHC6691_n2155 (.O(FE_PHN6691_n2155), 
	.I(FE_PHN4956_n2155));
   BUFMHD FE_PHC6690_n2135 (.O(FE_PHN6690_n2135), 
	.I(FE_PHN7260_n2135));
   BUFCHD FE_PHC6689_n2164 (.O(FE_PHN6689_n2164), 
	.I(FE_PHN7250_n2164));
   BUFHHD FE_PHC6688_n2592 (.O(FE_PHN6688_n2592), 
	.I(n2592));
   BUFCHD FE_PHC6687_n2394 (.O(FE_PHN6687_n2394), 
	.I(FE_PHN7229_n2394));
   BUFCHD FE_PHC6686_n4155 (.O(FE_PHN6686_n4155), 
	.I(FE_PHN7235_n4155));
   BUFMHD FE_PHC6685_n2379 (.O(FE_PHN6685_n2379), 
	.I(FE_PHN7274_n2379));
   BUFCHD FE_PHC6684_n4002 (.O(FE_PHN6684_n4002), 
	.I(FE_PHN7266_n4002));
   BUFCHD FE_PHC6683_n2604 (.O(FE_PHN6683_n2604), 
	.I(FE_PHN4862_n2604));
   BUFCHD FE_PHC6682_n2165 (.O(FE_PHN6682_n2165), 
	.I(FE_PHN7257_n2165));
   BUFCHD FE_PHC6681_n2625 (.O(FE_PHN6681_n2625), 
	.I(FE_PHN7227_n2625));
   BUFCHD FE_PHC6680_n2159 (.O(FE_PHN6680_n2159), 
	.I(FE_PHN7226_n2159));
   BUFCHD FE_PHC6679_n2132 (.O(FE_PHN6679_n2132), 
	.I(FE_PHN7239_n2132));
   BUFCKEHD FE_PHC6678_n4102 (.O(FE_PHN6678_n4102), 
	.I(FE_PHN7216_n4102));
   BUFCKLHD FE_PHC6677_n2603 (.O(FE_PHN6677_n2603), 
	.I(FE_PHN4890_n2603));
   BUFCHD FE_PHC6676_n3934 (.O(FE_PHN6676_n3934), 
	.I(FE_PHN7247_n3934));
   BUFCHD FE_PHC6675_n3960 (.O(FE_PHN6675_n3960), 
	.I(FE_PHN7243_n3960));
   BUFCKEHD FE_PHC6674_n1863 (.O(FE_PHN6674_n1863), 
	.I(FE_PHN7218_n1863));
   BUFCKLHD FE_PHC6673_n2582 (.O(FE_PHN6673_n2582), 
	.I(FE_PHN7224_n2582));
   BUFCHD FE_PHC6672_n2151 (.O(FE_PHN6672_n2151), 
	.I(FE_PHN7270_n2151));
   BUFCHD FE_PHC6671_n2119 (.O(FE_PHN6671_n2119), 
	.I(FE_PHN7271_n2119));
   BUFCKLHD FE_PHC6670_n2427 (.O(FE_PHN6670_n2427), 
	.I(FE_PHN7269_n2427));
   BUFCHD FE_PHC6669_n4147 (.O(FE_PHN6669_n4147), 
	.I(FE_PHN7222_n4147));
   BUFEHD FE_PHC6668_n4163 (.O(FE_PHN6668_n4163), 
	.I(FE_PHN7215_n4163));
   BUFCKEHD FE_PHC6667_n2628 (.O(FE_PHN6667_n2628), 
	.I(FE_PHN7219_n2628));
   BUFCHD FE_PHC6666_n4365 (.O(FE_PHN6666_n4365), 
	.I(FE_PHN7284_n4365));
   BUFCKLHD FE_PHC6665_n2417 (.O(FE_PHN6665_n2417), 
	.I(FE_PHN7236_n2417));
   BUFCHD FE_PHC6664_n2892 (.O(FE_PHN6664_n2892), 
	.I(FE_PHN7276_n2892));
   BUFMHD FE_PHC6663_n2393 (.O(FE_PHN6663_n2393), 
	.I(FE_PHN7253_n2393));
   BUFCHD FE_PHC6662_n2169 (.O(FE_PHN6662_n2169), 
	.I(FE_PHN7252_n2169));
   BUFCHD FE_PHC6661_n4153 (.O(FE_PHN6661_n4153), 
	.I(FE_PHN7245_n4153));
   BUFCKIHD FE_PHC6660_n2170 (.O(FE_PHN6660_n2170), 
	.I(FE_PHN7225_n2170));
   BUFCHD FE_PHC6659_n4139 (.O(FE_PHN6659_n4139), 
	.I(FE_PHN7399_n4139));
   BUFCKIHD FE_PHC6658_n2130 (.O(FE_PHN6658_n2130), 
	.I(n2130));
   BUFMHD FE_PHC6657_n2434 (.O(FE_PHN6657_n2434), 
	.I(FE_PHN7264_n2434));
   BUFMHD FE_PHC6656_n2118 (.O(FE_PHN6656_n2118), 
	.I(FE_PHN4866_n2118));
   BUFCKLHD FE_PHC6655_n2426 (.O(FE_PHN6655_n2426), 
	.I(FE_PHN7279_n2426));
   BUFCHD FE_PHC6654_n3968 (.O(FE_PHN6654_n3968), 
	.I(FE_PHN7237_n3968));
   BUFCKLHD FE_PHC6653_n2378 (.O(FE_PHN6653_n2378), 
	.I(FE_PHN7258_n2378));
   BUFCKLHD FE_PHC6652_n2578 (.O(FE_PHN6652_n2578), 
	.I(FE_PHN7241_n2578));
   BUFCHD FE_PHC6651_n3923 (.O(FE_PHN6651_n3923), 
	.I(FE_PHN7240_n3923));
   BUFCKLHD FE_PHC6650_n2571 (.O(FE_PHN6650_n2571), 
	.I(FE_PHN7246_n2571));
   BUFCHD FE_PHC6649_n2402 (.O(FE_PHN6649_n2402), 
	.I(FE_PHN7228_n2402));
   BUFCHD FE_PHC6648_n4121 (.O(FE_PHN6648_n4121), 
	.I(FE_PHN7233_n4121));
   BUFCKLHD FE_PHC6647_n2425 (.O(FE_PHN6647_n2425), 
	.I(FE_PHN7275_n2425));
   BUFCKLHD FE_PHC6646_n2395 (.O(FE_PHN6646_n2395), 
	.I(FE_PHN7267_n2395));
   BUFCKLHD FE_PHC6645_n2410 (.O(FE_PHN6645_n2410), 
	.I(FE_PHN4803_n2410));
   BUFCHD FE_PHC6644_n2168 (.O(FE_PHN6644_n2168), 
	.I(FE_PHN7256_n2168));
   BUFCKLHD FE_PHC6643_n2377 (.O(FE_PHN6643_n2377), 
	.I(FE_PHN7273_n2377));
   BUFCHD FE_PHC6642_n4011 (.O(FE_PHN6642_n4011), 
	.I(FE_PHN7272_n4011));
   BUFCHD FE_PHC6641_n2152 (.O(FE_PHN6641_n2152), 
	.I(FE_PHN7251_n2152));
   BUFCHD FE_PHC6640_n2414 (.O(FE_PHN6640_n2414), 
	.I(FE_PHN4936_n2414));
   BUFCHD FE_PHC6639_n2397 (.O(FE_PHN6639_n2397), 
	.I(FE_PHN4917_n2397));
   BUFCHD FE_PHC6638_n2921 (.O(FE_PHN6638_n2921), 
	.I(FE_PHN4899_n2921));
   BUFCKEHD FE_PHC6637_n2743 (.O(FE_PHN6637_n2743), 
	.I(FE_PHN7195_n2743));
   BUFCKEHD FE_PHC6636_n2749 (.O(FE_PHN6636_n2749), 
	.I(FE_PHN7191_n2749));
   BUFCKEHD FE_PHC6635_n2122 (.O(FE_PHN6635_n2122), 
	.I(FE_PHN7184_n2122));
   BUFCKEHD FE_PHC6634_n2176 (.O(FE_PHN6634_n2176), 
	.I(FE_PHN7172_n2176));
   BUFCKEHD FE_PHC6633_n2589 (.O(FE_PHN6633_n2589), 
	.I(FE_PHN7196_n2589));
   BUFCKEHD FE_PHC6632_n4158 (.O(FE_PHN6632_n4158), 
	.I(FE_PHN7173_n4158));
   BUFCKEHD FE_PHC6631_n4062 (.O(FE_PHN6631_n4062), 
	.I(FE_PHN7157_n4062));
   BUFCKEHD FE_PHC6630_n3965 (.O(FE_PHN6630_n3965), 
	.I(FE_PHN7162_n3965));
   BUFCHD FE_PHC6629_n1913 (.O(FE_PHN6629_n1913), 
	.I(FE_PHN7209_n1913));
   BUFCHD FE_PHC6628_n4135 (.O(FE_PHN6628_n4135), 
	.I(FE_PHN7211_n4135));
   BUFCHD FE_PHC6627_n2697 (.O(FE_PHN6627_n2697), 
	.I(FE_PHN7203_n2697));
   BUFCHD FE_PHC6626_n3033 (.O(FE_PHN6626_n3033), 
	.I(FE_PHN7165_n3033));
   BUFCKEHD FE_PHC6625_n2609 (.O(FE_PHN6625_n2609), 
	.I(FE_PHN7199_n2609));
   BUFCKEHD FE_PHC6624_n4107 (.O(FE_PHN6624_n4107), 
	.I(FE_PHN7207_n4107));
   BUFCKEHD FE_PHC6623_n3944 (.O(FE_PHN6623_n3944), 
	.I(FE_PHN7202_n3944));
   BUFCKEHD FE_PHC6622_n2123 (.O(FE_PHN6622_n2123), 
	.I(FE_PHN7198_n2123));
   BUFEHD FE_PHC6621_n3034 (.O(FE_PHN6621_n3034), 
	.I(FE_PHN4004_n3034));
   BUFCHD FE_PHC6620_n921 (.O(FE_PHN6620_n921), 
	.I(FE_PHN7200_n921));
   BUFCHD FE_PHC6619_n1908 (.O(FE_PHN6619_n1908), 
	.I(FE_PHN7187_n1908));
   BUFEHD FE_PHC6618_n1375 (.O(FE_PHN6618_n1375), 
	.I(FE_PHN4872_n1375));
   BUFEHD FE_PHC6617_n2908 (.O(FE_PHN6617_n2908), 
	.I(FE_PHN4808_n2908));
   BUFCKEHD FE_PHC6616_n2257 (.O(FE_PHN6616_n2257), 
	.I(FE_PHN7116_n2257));
   BUFCHD FE_PHC6615_n4151 (.O(FE_PHN6615_n4151), 
	.I(FE_PHN7182_n4151));
   BUFCHD FE_PHC6614_n2624 (.O(FE_PHN6614_n2624), 
	.I(FE_PHN7176_n2624));
   BUFEHD FE_PHC6613_n1865 (.O(FE_PHN6613_n1865), 
	.I(FE_PHN4949_n1865));
   BUFEHD FE_PHC6612_n2386 (.O(FE_PHN6612_n2386), 
	.I(FE_PHN4848_n2386));
   BUFCHD FE_PHC6611_n3004 (.O(FE_PHN6611_n3004), 
	.I(FE_PHN4001_n3004));
   BUFCHD FE_PHC6610_n4150 (.O(FE_PHN6610_n4150), 
	.I(FE_PHN7158_n4150));
   BUFEHD FE_PHC6609_n2390 (.O(FE_PHN6609_n2390), 
	.I(FE_PHN4814_n2390));
   BUFCHD FE_PHC6608_n3017 (.O(FE_PHN6608_n3017), 
	.I(FE_PHN7206_n3017));
   BUFCHD FE_PHC6607_n2626 (.O(FE_PHN6607_n2626), 
	.I(FE_PHN7146_n2626));
   BUFIHD FE_PHC6606_n2422 (.O(FE_PHN6606_n2422), 
	.I(FE_PHN7208_n2422));
   BUFCKEHD FE_PHC6605_n2876 (.O(FE_PHN6605_n2876), 
	.I(FE_PHN7111_n2876));
   BUFCHD FE_PHC6604_n2577 (.O(FE_PHN6604_n2577), 
	.I(FE_PHN7106_n2577));
   BUFCKEHD FE_PHC6603_n3150 (.O(FE_PHN6603_n3150), 
	.I(FE_PHN7212_n3150));
   BUFCHD FE_PHC6602_n3047 (.O(FE_PHN6602_n3047), 
	.I(FE_PHN7190_n3047));
   BUFCKEHD FE_PHC6601_n2177 (.O(FE_PHN6601_n2177), 
	.I(FE_PHN7197_n2177));
   BUFCHD FE_PHC6600_n2406 (.O(FE_PHN6600_n2406), 
	.I(FE_PHN7084_n2406));
   BUFCHD FE_PHC6599_n2587 (.O(FE_PHN6599_n2587), 
	.I(FE_PHN7119_n2587));
   BUFCHD FE_PHC6598_n1012 (.O(FE_PHN6598_n1012), 
	.I(FE_PHN7179_n1012));
   BUFEHD FE_PHC6597_n985 (.O(FE_PHN6597_n985), 
	.I(FE_PHN7129_n985));
   BUFCHD FE_PHC6596_n973 (.O(FE_PHN6596_n973), 
	.I(FE_PHN7192_n973));
   BUFCKEHD FE_PHC6595_n2701 (.O(FE_PHN6595_n2701), 
	.I(FE_PHN7170_n2701));
   BUFCHD FE_PHC6594_n1007 (.O(FE_PHN6594_n1007), 
	.I(FE_PHN7151_n1007));
   BUFCKEHD FE_PHC6593_n2873 (.O(FE_PHN6593_n2873), 
	.I(FE_PHN7194_n2873));
   BUFCHD FE_PHC6592_n2919 (.O(FE_PHN6592_n2919), 
	.I(FE_PHN7175_n2919));
   BUFCHD FE_PHC6591_n2398 (.O(FE_PHN6591_n2398), 
	.I(FE_PHN7112_n2398));
   BUFCKEHD FE_PHC6590_n2171 (.O(FE_PHN6590_n2171), 
	.I(FE_PHN7188_n2171));
   BUFCHD FE_PHC6589_n2938 (.O(FE_PHN6589_n2938), 
	.I(FE_PHN7134_n2938));
   BUFCHD FE_PHC6588_n1003 (.O(FE_PHN6588_n1003), 
	.I(FE_PHN7145_n1003));
   BUFCKEHD FE_PHC6587_n1286 (.O(FE_PHN6587_n1286), 
	.I(FE_PHN7149_n1286));
   BUFCHD FE_PHC6586_n2889 (.O(FE_PHN6586_n2889), 
	.I(FE_PHN7164_n2889));
   BUFCKEHD FE_PHC6585_n2161 (.O(FE_PHN6585_n2161), 
	.I(FE_PHN7142_n2161));
   BUFCHD FE_PHC6584_n3021 (.O(FE_PHN6584_n3021), 
	.I(FE_PHN7189_n3021));
   BUFCHD FE_PHC6583_n1028 (.O(FE_PHN6583_n1028), 
	.I(FE_PHN7193_n1028));
   BUFCHD FE_PHC6582_n2619 (.O(FE_PHN6582_n2619), 
	.I(FE_PHN7076_n2619));
   BUFCHD FE_PHC6581_n981 (.O(FE_PHN6581_n981), 
	.I(FE_PHN7177_n981));
   BUFCKEHD FE_PHC6580_n2590 (.O(FE_PHN6580_n2590), 
	.I(FE_PHN7186_n2590));
   BUFCHD FE_PHC6579_n977 (.O(FE_PHN6579_n977), 
	.I(FE_PHN4920_n977));
   BUFCHD FE_PHC6578_n2893 (.O(FE_PHN6578_n2893), 
	.I(FE_PHN7150_n2893));
   BUFCKEHD FE_PHC6577_n2616 (.O(FE_PHN6577_n2616), 
	.I(FE_PHN7180_n2616));
   BUFCKEHD FE_PHC6576_n2857 (.O(FE_PHN6576_n2857), 
	.I(FE_PHN7121_n2857));
   BUFCHD FE_PHC6575_n983 (.O(FE_PHN6575_n983), 
	.I(FE_PHN7127_n983));
   BUFCKEHD FE_PHC6574_n2428 (.O(FE_PHN6574_n2428), 
	.I(FE_PHN7066_n2428));
   BUFCHD FE_PHC6573_n2907 (.O(FE_PHN6573_n2907), 
	.I(FE_PHN7148_n2907));
   BUFCHD FE_PHC6572_n1086 (.O(FE_PHN6572_n1086), 
	.I(FE_PHN7205_n1086));
   BUFCHD FE_PHC6571_n2381 (.O(FE_PHN6571_n2381), 
	.I(FE_PHN7185_n2381));
   BUFCHD FE_PHC6570_n2925 (.O(FE_PHN6570_n2925), 
	.I(FE_PHN7140_n2925));
   BUFCHD FE_PHC6569_n2941 (.O(FE_PHN6569_n2941), 
	.I(FE_PHN7131_n2941));
   BUFCHD FE_PHC6568_n896 (.O(FE_PHN6568_n896), 
	.I(FE_PHN3998_n896));
   BUFCKEHD FE_PHC6567_n2750 (.O(FE_PHN6567_n2750), 
	.I(FE_PHN7086_n2750));
   BUFCKEHD FE_PHC6566_n2375 (.O(FE_PHN6566_n2375), 
	.I(FE_PHN7128_n2375));
   BUFCHD FE_PHC6565_n2696 (.O(FE_PHN6565_n2696), 
	.I(FE_PHN7123_n2696));
   BUFNHD FE_PHC6564_n1158 (.O(FE_PHN6564_n1158), 
	.I(n1158));
   BUFEHD FE_PHC6563_n4012 (.O(FE_PHN6563_n4012), 
	.I(FE_PHN7133_n4012));
   BUFCHD FE_PHC6562_n1019 (.O(FE_PHN6562_n1019), 
	.I(FE_PHN7147_n1019));
   BUFCKEHD FE_PHC6561_n2407 (.O(FE_PHN6561_n2407), 
	.I(FE_PHN7103_n2407));
   BUFCHD FE_PHC6560_n2181 (.O(FE_PHN6560_n2181), 
	.I(FE_PHN7095_n2181));
   BUFCHD FE_PHC6559_n996 (.O(FE_PHN6559_n996), 
	.I(FE_PHN7126_n996));
   BUFCHD FE_PHC6558_n1031 (.O(FE_PHN6558_n1031), 
	.I(FE_PHN7097_n1031));
   BUFEHD FE_PHC6557_n1094 (.O(FE_PHN6557_n1094), 
	.I(FE_PHN7064_n1094));
   BUFCHD FE_PHC6556_n2429 (.O(FE_PHN6556_n2429), 
	.I(FE_PHN7083_n2429));
   BUFCHD FE_PHC6555_n2566 (.O(FE_PHN6555_n2566), 
	.I(FE_PHN7099_n2566));
   BUFCHD FE_PHC6554_n2695 (.O(FE_PHN6554_n2695), 
	.I(FE_PHN7101_n2695));
   BUFCHD FE_PHC6553_n980 (.O(FE_PHN6553_n980), 
	.I(FE_PHN7094_n980));
   BUFCKEHD FE_PHC6552_n2144 (.O(FE_PHN6552_n2144), 
	.I(FE_PHN7139_n2144));
   BUFCHD FE_PHC6551_n2172 (.O(FE_PHN6551_n2172), 
	.I(FE_PHN7081_n2172));
   BUFCHD FE_PHC6550_n2125 (.O(FE_PHN6550_n2125), 
	.I(FE_PHN7125_n2125));
   BUFCKEHD FE_PHC6549_n2411 (.O(FE_PHN6549_n2411), 
	.I(FE_PHN7058_n2411));
   BUFCKIHD FE_PHC6548_n1015 (.O(FE_PHN6548_n1015), 
	.I(FE_PHN7071_n1015));
   BUFCHD FE_PHC6547_n967 (.O(FE_PHN6547_n967), 
	.I(FE_PHN7178_n967));
   BUFHHD FE_PHC6546_n979 (.O(FE_PHN6546_n979), 
	.I(FE_PHN7074_n979));
   BUFCHD FE_PHC6545_n880 (.O(FE_PHN6545_n880), 
	.I(FE_PHN7210_n880));
   BUFCHD FE_PHC6544_n2611 (.O(FE_PHN6544_n2611), 
	.I(FE_PHN7062_n2611));
   BUFCHD FE_PHC6543_n3945 (.O(FE_PHN6543_n3945), 
	.I(FE_PHN7155_n3945));
   BUFCHD FE_PHC6542_n4210 (.O(FE_PHN6542_n4210), 
	.I(FE_PHN7136_n4210));
   BUFCHD FE_PHC6541_n2148 (.O(FE_PHN6541_n2148), 
	.I(FE_PHN7102_n2148));
   BUFCHD FE_PHC6540_n1001 (.O(FE_PHN6540_n1001), 
	.I(FE_PHN7031_n1001));
   BUFCHD FE_PHC6539_n2747 (.O(FE_PHN6539_n2747), 
	.I(FE_PHN7091_n2747));
   BUFCHD FE_PHC6538_n2594 (.O(FE_PHN6538_n2594), 
	.I(FE_PHN7051_n2594));
   BUFCHD FE_PHC6537_n4018 (.O(FE_PHN6537_n4018), 
	.I(FE_PHN7075_n4018));
   BUFCHD FE_PHC6536_n2618 (.O(FE_PHN6536_n2618), 
	.I(FE_PHN7046_n2618));
   BUFCHD FE_PHC6535_n2424 (.O(FE_PHN6535_n2424), 
	.I(FE_PHN7105_n2424));
   BUFCHD FE_PHC6534_n1054 (.O(FE_PHN6534_n1054), 
	.I(FE_PHN7100_n1054));
   BUFCHD FE_PHC6533_n898 (.O(FE_PHN6533_n898), 
	.I(FE_PHN4005_n898));
   BUFCHD FE_PHC6532_n4403 (.O(FE_PHN6532_n4403), 
	.I(FE_PHN3981_n4403));
   BUFCHD FE_PHC6531_n3980 (.O(FE_PHN6531_n3980), 
	.I(FE_PHN7115_n3980));
   BUFCHD FE_PHC6530_n1154 (.O(FE_PHN6530_n1154), 
	.I(FE_PHN7042_n1154));
   BUFCHD FE_PHC6529_n3981 (.O(FE_PHN6529_n3981), 
	.I(FE_PHN7092_n3981));
   BUFCHD FE_PHC6528_n2602 (.O(FE_PHN6528_n2602), 
	.I(FE_PHN7037_n2602));
   BUFCHD FE_PHC6527_n1190 (.O(FE_PHN6527_n1190), 
	.I(FE_PHN7069_n1190));
   BUFCHD FE_PHC6526_n4016 (.O(FE_PHN6526_n4016), 
	.I(FE_PHN7204_n4016));
   BUFCHD FE_PHC6525_n962 (.O(FE_PHN6525_n962), 
	.I(FE_PHN7110_n962));
   BUFCHD FE_PHC6524_n2376 (.O(FE_PHN6524_n2376), 
	.I(FE_PHN7070_n2376));
   BUFCHD FE_PHC6523_n2576 (.O(FE_PHN6523_n2576), 
	.I(FE_PHN7035_n2576));
   BUFCHD FE_PHC6522_n2423 (.O(FE_PHN6522_n2423), 
	.I(FE_PHN7054_n2423));
   BUFCHD FE_PHC6521_n3932 (.O(FE_PHN6521_n3932), 
	.I(FE_PHN7053_n3932));
   BUFCHD FE_PHC6520_n4358 (.O(FE_PHN6520_n4358), 
	.I(FE_PHN7161_n4358));
   BUFCHD FE_PHC6519_n4259 (.O(FE_PHN6519_n4259), 
	.I(FE_PHN7163_n4259));
   BUFCHD FE_PHC6518_n1178 (.O(FE_PHN6518_n1178), 
	.I(FE_PHN7061_n1178));
   BUFCHD FE_PHC6517_n953 (.O(FE_PHN6517_n953), 
	.I(FE_PHN7040_n953));
   BUFCHD FE_PHC6516_n917 (.O(FE_PHN6516_n917), 
	.I(FE_PHN7118_n917));
   BUFCHD FE_PHC6515_n3962 (.O(FE_PHN6515_n3962), 
	.I(FE_PHN7201_n3962));
   BUFCHD FE_PHC6514_n2622 (.O(FE_PHN6514_n2622), 
	.I(FE_PHN7041_n2622));
   BUFCHD FE_PHC6513_n3971 (.O(FE_PHN6513_n3971), 
	.I(FE_PHN7089_n3971));
   BUFCHD FE_PHC6512_n2380 (.O(FE_PHN6512_n2380), 
	.I(FE_PHN7068_n2380));
   BUFCHD FE_PHC6511_n4274 (.O(FE_PHN6511_n4274), 
	.I(FE_PHN7122_n4274));
   BUFCHD FE_PHC6510_n2572 (.O(FE_PHN6510_n2572), 
	.I(FE_PHN7028_n2572));
   BUFCHD FE_PHC6509_n2156 (.O(FE_PHN6509_n2156), 
	.I(FE_PHN7072_n2156));
   BUFCHD FE_PHC6508_n888 (.O(FE_PHN6508_n888), 
	.I(FE_PHN7144_n888));
   BUFCHD FE_PHC6507_n4294 (.O(FE_PHN6507_n4294), 
	.I(FE_PHN7085_n4294));
   BUFHHD FE_PHC6506_n4114 (.O(FE_PHN6506_n4114), 
	.I(FE_PHN4857_n4114));
   BUFCHD FE_PHC6505_n949 (.O(FE_PHN6505_n949), 
	.I(FE_PHN7104_n949));
   BUFCHD FE_PHC6504_n4391 (.O(FE_PHN6504_n4391), 
	.I(FE_PHN3258_n4391));
   BUFCHD FE_PHC6503_n2251 (.O(FE_PHN6503_n2251), 
	.I(FE_PHN7027_n2251));
   BUFCHD FE_PHC6502_n3212 (.O(FE_PHN6502_n3212), 
	.I(FE_PHN7153_n3212));
   BUFCHD FE_PHC6501_n2412 (.O(FE_PHN6501_n2412), 
	.I(FE_PHN7030_n2412));
   BUFCHD FE_PHC6500_n4035 (.O(FE_PHN6500_n4035), 
	.I(FE_PHN7159_n4035));
   BUFCKMHD FE_PHC6499_n2615 (.O(FE_PHN6499_n2615), 
	.I(FE_PHN7093_n2615));
   BUFCHD FE_PHC6498_n2131 (.O(FE_PHN6498_n2131), 
	.I(FE_PHN7078_n2131));
   BUFCHD FE_PHC6497_n1872 (.O(FE_PHN6497_n1872), 
	.I(FE_PHN7060_n1872));
   BUFCHD FE_PHC6496_n4308 (.O(FE_PHN6496_n4308), 
	.I(FE_PHN7143_n4308));
   BUFHHD FE_PHC6495_n1874 (.O(FE_PHN6495_n1874), 
	.I(FE_PHN3853_n1874));
   BUFCHD FE_PHC6494_n2388 (.O(FE_PHN6494_n2388), 
	.I(FE_PHN7032_n2388));
   BUFCHD FE_PHC6493_n3970 (.O(FE_PHN6493_n3970), 
	.I(FE_PHN7080_n3970));
   BUFCHD FE_PHC6492_n4034 (.O(FE_PHN6492_n4034), 
	.I(FE_PHN7141_n4034));
   BUFCHD FE_PHC6491_n1922 (.O(FE_PHN6491_n1922), 
	.I(FE_PHN7038_n1922));
   BUFCHD FE_PHC6490_n3955 (.O(FE_PHN6490_n3955), 
	.I(FE_PHN7077_n3955));
   BUFCHD FE_PHC6489_n4404 (.O(FE_PHN6489_n4404), 
	.I(FE_PHN7169_n4404));
   BUFCHD FE_PHC6488_n4273 (.O(FE_PHN6488_n4273), 
	.I(FE_PHN7098_n4273));
   BUFCHD FE_PHC6487_n2935 (.O(FE_PHN6487_n2935), 
	.I(FE_PHN7183_n2935));
   BUFCHD FE_PHC6486_n2968 (.O(FE_PHN6486_n2968), 
	.I(FE_PHN3697_n2968));
   BUFCHD FE_PHC6485_n4374 (.O(FE_PHN6485_n4374), 
	.I(FE_PHN3287_n4374));
   BUFCHD FE_PHC6484_n3260 (.O(FE_PHN6484_n3260), 
	.I(FE_PHN7117_n3260));
   BUFCHD FE_PHC6483_n2138 (.O(FE_PHN6483_n2138), 
	.I(FE_PHN7048_n2138));
   BUFCHD FE_PHC6482_n4242 (.O(FE_PHN6482_n4242), 
	.I(FE_PHN7124_n4242));
   BUFCKLHD FE_PHC6481_n1906 (.O(FE_PHN6481_n1906), 
	.I(FE_PHN7114_n1906));
   BUFCHD FE_PHC6480_n1918 (.O(FE_PHN6480_n1918), 
	.I(FE_PHN7056_n1918));
   BUFCHD FE_PHC6479_n938 (.O(FE_PHN6479_n938), 
	.I(FE_PHN7034_n938));
   BUFCHD FE_PHC6478_n4370 (.O(FE_PHN6478_n4370), 
	.I(FE_PHN4000_n4370));
   BUFCHD FE_PHC6477_n964 (.O(FE_PHN6477_n964), 
	.I(FE_PHN7055_n964));
   BUFCHD FE_PHC6476_n906 (.O(FE_PHN6476_n906), 
	.I(FE_PHN7050_n906));
   BUFCHD FE_PHC6475_n2163 (.O(FE_PHN6475_n2163), 
	.I(FE_PHN7088_n2163));
   BUFCHD FE_PHC6474_n2598 (.O(FE_PHN6474_n2598), 
	.I(FE_PHN3769_n2598));
   BUFCHD FE_PHC6473_n950 (.O(FE_PHN6473_n950), 
	.I(FE_PHN7052_n950));
   BUFCHD FE_PHC6472_n901 (.O(FE_PHN6472_n901), 
	.I(FE_PHN7130_n901));
   BUFCHD FE_PHC6471_n2612 (.O(FE_PHN6471_n2612), 
	.I(FE_PHN7026_n2612));
   BUFCHD FE_PHC6470_n944 (.O(FE_PHN6470_n944), 
	.I(FE_PHN7065_n944));
   BUFCKLHD FE_PHC6469_n2121 (.O(FE_PHN6469_n2121), 
	.I(FE_PHN7079_n2121));
   BUFCHD FE_PHC6468_n933 (.O(FE_PHN6468_n933), 
	.I(FE_PHN7108_n933));
   BUFCKLHD FE_PHC6467_n2419 (.O(FE_PHN6467_n2419), 
	.I(FE_PHN7096_n2419));
   BUFCHD FE_PHC6466_n3983 (.O(FE_PHN6466_n3983), 
	.I(FE_PHN7120_n3983));
   BUFCHD FE_PHC6465_n2124 (.O(FE_PHN6465_n2124), 
	.I(FE_PHN7045_n2124));
   BUFCHD FE_PHC6464_n4116 (.O(FE_PHN6464_n4116), 
	.I(FE_PHN7059_n4116));
   BUFCKEHD FE_PHC6463_n1880 (.O(FE_PHN6463_n1880), 
	.I(FE_PHN7043_n1880));
   BUFCHD FE_PHC6462_n4032 (.O(FE_PHN6462_n4032), 
	.I(FE_PHN7135_n4032));
   BUFCHD FE_PHC6461_n3966 (.O(FE_PHN6461_n3966), 
	.I(FE_PHN7087_n3966));
   BUFCHD FE_PHC6460_n2137 (.O(FE_PHN6460_n2137), 
	.I(FE_PHN7049_n2137));
   BUFCHD FE_PHC6459_n3979 (.O(FE_PHN6459_n3979), 
	.I(FE_PHN7137_n3979));
   BUFCHD FE_PHC6458_n4148 (.O(FE_PHN6458_n4148), 
	.I(FE_PHN7057_n4148));
   BUFCKLHD FE_PHC6457_n2403 (.O(FE_PHN6457_n2403), 
	.I(FE_PHN7132_n2403));
   BUFCHD FE_PHC6456_n1919 (.O(FE_PHN6456_n1919), 
	.I(FE_PHN7036_n1919));
   BUFCHD FE_PHC6455_n927 (.O(FE_PHN6455_n927), 
	.I(FE_PHN7067_n927));
   BUFCHD FE_PHC6454_n4008 (.O(FE_PHN6454_n4008), 
	.I(FE_PHN7174_n4008));
   BUFCHD FE_PHC6453_n2904 (.O(FE_PHN6453_n2904), 
	.I(FE_PHN7171_n2904));
   BUFCHD FE_PHC6452_n2922 (.O(FE_PHN6452_n2922), 
	.I(FE_PHN7154_n2922));
   BUFCHD FE_PHC6451_n3000 (.O(FE_PHN6451_n3000), 
	.I(FE_PHN3738_n3000));
   BUFCHD FE_PHC6450_n4027 (.O(FE_PHN6450_n4027), 
	.I(FE_PHN7090_n4027));
   BUFCHD FE_PHC6449_n2985 (.O(FE_PHN6449_n2985), 
	.I(FE_PHN3646_n2985));
   BUFCKLHD FE_PHC6448_n2382 (.O(FE_PHN6448_n2382), 
	.I(FE_PHN7082_n2382));
   BUFCHD FE_PHC6447_n2149 (.O(FE_PHN6447_n2149), 
	.I(FE_PHN7047_n2149));
   BUFCHD FE_PHC6446_n4331 (.O(FE_PHN6446_n4331), 
	.I(FE_PHN7168_n4331));
   BUFCKLHD FE_PHC6445_n2401 (.O(FE_PHN6445_n2401), 
	.I(FE_PHN7073_n2401));
   BUFCKLHD FE_PHC6444_n2432 (.O(FE_PHN6444_n2432), 
	.I(FE_PHN7138_n2432));
   BUFCHD FE_PHC6443_n4142 (.O(FE_PHN6443_n4142), 
	.I(FE_PHN7044_n4142));
   BUFCHD FE_PHC6442_n4110 (.O(FE_PHN6442_n4110), 
	.I(FE_PHN7033_n4110));
   BUFCHD FE_PHC6441_n930 (.O(FE_PHN6441_n930), 
	.I(FE_PHN7109_n930));
   BUFCHD FE_PHC6440_n914 (.O(FE_PHN6440_n914), 
	.I(FE_PHN7107_n914));
   BUFCHD FE_PHC6439_n4031 (.O(FE_PHN6439_n4031), 
	.I(FE_PHN7113_n4031));
   BUFCKEHD FE_PHC6438_n2605 (.O(FE_PHN6438_n2605), 
	.I(FE_PHN3955_n2605));
   BUFCKEHD FE_PHC6437_n1904 (.O(FE_PHN6437_n1904), 
	.I(FE_PHN4236_n1904));
   BUFCKEHD FE_PHC6436_n904 (.O(FE_PHN6436_n904), 
	.I(FE_PHN4338_n904));
   BUFCKEHD FE_PHC6435_n3109 (.O(FE_PHN6435_n3109), 
	.I(FE_PHN3850_n3109));
   BUFCHD FE_PHC6434_n4123 (.O(FE_PHN6434_n4123), 
	.I(n4123));
   BUFCKEHD FE_PHC6433_n4244 (.O(FE_PHN6433_n4244), 
	.I(FE_PHN3474_n4244));
   BUFCHD FE_PHC6432_n3066 (.O(FE_PHN6432_n3066), 
	.I(FE_PHN3967_n3066));
   BUFCHD FE_PHC6431_n3911 (.O(FE_PHN6431_n3911), 
	.I(FE_PHN3561_n3911));
   BUFCKEHD FE_PHC6430_n3005 (.O(FE_PHN6430_n3005), 
	.I(FE_PHN4306_n3005));
   BUFCKEHD FE_PHC6429_n4285 (.O(FE_PHN6429_n4285), 
	.I(FE_PHN4496_n4285));
   BUFCHD FE_PHC6428_n3119 (.O(FE_PHN6428_n3119), 
	.I(FE_PHN3851_n3119));
   BUFCKEHD FE_PHC6427_ram_98__3_ (.O(FE_PHN6427_ram_98__3_), 
	.I(FE_PHN4087_ram_98__3_));
   BUFCKEHD FE_PHC6426_n3030 (.O(FE_PHN6426_n3030), 
	.I(FE_PHN3245_n3030));
   BUFCKEHD FE_PHC6425_n2262 (.O(FE_PHN6425_n2262), 
	.I(FE_PHN5637_n2262));
   BUFCKEHD FE_PHC6424_n4367 (.O(FE_PHN6424_n4367), 
	.I(FE_PHN3621_n4367));
   BUFCHD FE_PHC6423_n3140 (.O(FE_PHN6423_n3140), 
	.I(FE_PHN3547_n3140));
   BUFCKEHD FE_PHC6422_n2891 (.O(FE_PHN6422_n2891), 
	.I(FE_PHN3617_n2891));
   BUFCKEHD FE_PHC6421_n4146 (.O(FE_PHN6421_n4146), 
	.I(FE_PHN4115_n4146));
   BUFCKEHD FE_PHC6420_n2554 (.O(FE_PHN6420_n2554), 
	.I(FE_PHN3917_n2554));
   BUFCHD FE_PHC6419_n4363 (.O(FE_PHN6419_n4363), 
	.I(FE_PHN3417_n4363));
   BUFCHD FE_PHC6418_n3036 (.O(FE_PHN6418_n3036), 
	.I(FE_PHN3897_n3036));
   BUFCHD FE_PHC6417_n3241 (.O(FE_PHN6417_n3241), 
	.I(FE_PHN5612_n3241));
   BUFCHD FE_PHC6416_n2957 (.O(FE_PHN6416_n2957), 
	.I(FE_PHN3778_n2957));
   BUFCHD FE_PHC6415_n3135 (.O(FE_PHN6415_n3135), 
	.I(FE_PHN3995_n3135));
   BUFCHD FE_PHC6414_n4265 (.O(FE_PHN6414_n4265), 
	.I(FE_PHN3824_n4265));
   BUFCKEHD FE_PHC6413_n2910 (.O(FE_PHN6413_n2910), 
	.I(FE_PHN3265_n2910));
   BUFCHD FE_PHC6412_n2600 (.O(FE_PHN6412_n2600), 
	.I(FE_PHN3484_n2600));
   BUFCKEHD FE_PHC6411_n2974 (.O(FE_PHN6411_n2974), 
	.I(FE_PHN3448_n2974));
   BUFCHD FE_PHC6410_n4175 (.O(FE_PHN6410_n4175), 
	.I(FE_PHN3714_n4175));
   BUFCHD FE_PHC6409_n3123 (.O(FE_PHN6409_n3123), 
	.I(FE_PHN3468_n3123));
   BUFCKEHD FE_PHC6408_n2906 (.O(FE_PHN6408_n2906), 
	.I(FE_PHN6998_n2906));
   BUFCKEHD FE_PHC6407_n3999 (.O(FE_PHN6407_n3999), 
	.I(FE_PHN3240_n3999));
   BUFCKEHD FE_PHC6406_n3011 (.O(FE_PHN6406_n3011), 
	.I(FE_PHN3901_n3011));
   BUFCKEHD FE_PHC6405_n1023 (.O(FE_PHN6405_n1023), 
	.I(FE_PHN3882_n1023));
   BUFCHD FE_PHC6404_n4366 (.O(FE_PHN6404_n4366), 
	.I(FE_PHN3822_n4366));
   BUFCKEHD FE_PHC6403_n2960 (.O(FE_PHN6403_n2960), 
	.I(FE_PHN3677_n2960));
   BUFCHD FE_PHC6402_n3046 (.O(FE_PHN6402_n3046), 
	.I(FE_PHN3793_n3046));
   BUFCKEHD FE_PHC6401_n841 (.O(FE_PHN6401_n841), 
	.I(FE_PHN3811_n841));
   BUFCKEHD FE_PHC6400_n3265 (.O(FE_PHN6400_n3265), 
	.I(FE_PHN6984_n3265));
   BUFCKEHD FE_PHC6399_n1206 (.O(FE_PHN6399_n1206), 
	.I(FE_PHN5632_n1206));
   BUFCKEHD FE_PHC6398_n3139 (.O(FE_PHN6398_n3139), 
	.I(FE_PHN3942_n3139));
   BUFCHD FE_PHC6397_n3090 (.O(FE_PHN6397_n3090), 
	.I(FE_PHN3838_n3090));
   BUFCHD FE_PHC6396_n4261 (.O(FE_PHN6396_n4261), 
	.I(FE_PHN4472_n4261));
   BUFCKEHD FE_PHC6395_ram_17__14_ (.O(FE_PHN6395_ram_17__14_), 
	.I(FE_PHN3451_ram_17__14_));
   BUFCKEHD FE_PHC6394_n951 (.O(FE_PHN6394_n951), 
	.I(FE_PHN6980_n951));
   BUFCKEHD FE_PHC6393_n4170 (.O(FE_PHN6393_n4170), 
	.I(FE_PHN5628_n4170));
   BUFCHD FE_PHC6392_n4187 (.O(FE_PHN6392_n4187), 
	.I(FE_PHN4637_n4187));
   BUFCHD FE_PHC6391_n3091 (.O(FE_PHN6391_n3091), 
	.I(FE_PHN4531_n3091));
   BUFCKEHD FE_PHC6390_n3115 (.O(FE_PHN6390_n3115), 
	.I(FE_PHN3336_n3115));
   BUFCHD FE_PHC6389_n3085 (.O(FE_PHN6389_n3085), 
	.I(FE_PHN3911_n3085));
   BUFCHD FE_PHC6388_n2963 (.O(FE_PHN6388_n2963), 
	.I(FE_PHN3987_n2963));
   BUFCHD FE_PHC6387_n4267 (.O(FE_PHN6387_n4267), 
	.I(FE_PHN3632_n4267));
   BUFCHD FE_PHC6386_n4168 (.O(FE_PHN6386_n4168), 
	.I(FE_PHN4543_n4168));
   BUFCHD FE_PHC6385_n871 (.O(FE_PHN6385_n871), 
	.I(FE_PHN4234_n871));
   BUFCKEHD FE_PHC6384_n4138 (.O(FE_PHN6384_n4138), 
	.I(FE_PHN3493_n4138));
   BUFCKEHD FE_PHC6383_n4241 (.O(FE_PHN6383_n4241), 
	.I(FE_PHN3933_n4241));
   BUFCKEHD FE_PHC6382_n4266 (.O(FE_PHN6382_n4266), 
	.I(FE_PHN6975_n4266));
   BUFCKEHD FE_PHC6381_n863 (.O(FE_PHN6381_n863), 
	.I(FE_PHN3654_n863));
   BUFCHD FE_PHC6380_n2391 (.O(FE_PHN6380_n2391), 
	.I(FE_PHN3246_n2391));
   BUFCKEHD FE_PHC6379_n4201 (.O(FE_PHN6379_n4201), 
	.I(FE_PHN6981_n4201));
   BUFCHD FE_PHC6378_n3031 (.O(FE_PHN6378_n3031), 
	.I(FE_PHN3362_n3031));
   BUFCHD FE_PHC6377_n4254 (.O(FE_PHN6377_n4254), 
	.I(FE_PHN3360_n4254));
   BUFCHD FE_PHC6376_n976 (.O(FE_PHN6376_n976), 
	.I(FE_PHN3989_n976));
   BUFCKEHD FE_PHC6375_n991 (.O(FE_PHN6375_n991), 
	.I(FE_PHN3711_n991));
   BUFCKEHD FE_PHC6374_n3931 (.O(FE_PHN6374_n3931), 
	.I(FE_PHN6951_n3931));
   BUFCKEHD FE_PHC6373_n4316 (.O(FE_PHN6373_n4316), 
	.I(FE_PHN3615_n4316));
   BUFCKEHD FE_PHC6372_n3132 (.O(FE_PHN6372_n3132), 
	.I(FE_PHN3558_n3132));
   BUFCKEHD FE_PHC6371_n3083 (.O(FE_PHN6371_n3083), 
	.I(FE_PHN3719_n3083));
   BUFCHD FE_PHC6370_n4395 (.O(FE_PHN6370_n4395), 
	.I(FE_PHN3728_n4395));
   BUFCKEHD FE_PHC6369_n3137 (.O(FE_PHN6369_n3137), 
	.I(n3137));
   BUFCKEHD FE_PHC6368_n3117 (.O(FE_PHN6368_n3117), 
	.I(FE_PHN3609_n3117));
   BUFCHD FE_PHC6367_n4227 (.O(FE_PHN6367_n4227), 
	.I(FE_PHN4643_n4227));
   BUFCHD FE_PHC6366_n4276 (.O(FE_PHN6366_n4276), 
	.I(FE_PHN3961_n4276));
   BUFCKEHD FE_PHC6365_n952 (.O(FE_PHN6365_n952), 
	.I(FE_PHN3845_n952));
   BUFCKEHD FE_PHC6364_n3920 (.O(FE_PHN6364_n3920), 
	.I(FE_PHN5620_n3920));
   BUFCKEHD FE_PHC6363_n4231 (.O(FE_PHN6363_n4231), 
	.I(FE_PHN3800_n4231));
   BUFCHD FE_PHC6362_n4382 (.O(FE_PHN6362_n4382), 
	.I(FE_PHN4554_n4382));
   BUFCKEHD FE_PHC6361_n3064 (.O(FE_PHN6361_n3064), 
	.I(FE_PHN4460_n3064));
   BUFCKEHD FE_PHC6360_n1911 (.O(FE_PHN6360_n1911), 
	.I(FE_PHN3974_n1911));
   BUFCHD FE_PHC6359_n2990 (.O(FE_PHN6359_n2990), 
	.I(FE_PHN3805_n2990));
   BUFCHD FE_PHC6358_n3038 (.O(FE_PHN6358_n3038), 
	.I(FE_PHN3381_n3038));
   BUFCHD FE_PHC6357_n4213 (.O(FE_PHN6357_n4213), 
	.I(FE_PHN4451_n4213));
   BUFCHD FE_PHC6356_n968 (.O(FE_PHN6356_n968), 
	.I(FE_PHN3940_n968));
   BUFCHD FE_PHC6355_n4236 (.O(FE_PHN6355_n4236), 
	.I(FE_PHN3731_n4236));
   BUFCHD FE_PHC6354_n4375 (.O(FE_PHN6354_n4375), 
	.I(FE_PHN3425_n4375));
   BUFCKEHD FE_PHC6353_n3947 (.O(FE_PHN6353_n3947), 
	.I(FE_PHN6920_n3947));
   BUFCHD FE_PHC6352_n3118 (.O(FE_PHN6352_n3118), 
	.I(FE_PHN3472_n3118));
   BUFCKEHD FE_PHC6351_n3111 (.O(FE_PHN6351_n3111), 
	.I(FE_PHN3422_n3111));
   BUFCHD FE_PHC6350_n877 (.O(FE_PHN6350_n877), 
	.I(FE_PHN3464_n877));
   BUFCHD FE_PHC6349_n3065 (.O(FE_PHN6349_n3065), 
	.I(FE_PHN3489_n3065));
   BUFCKEHD FE_PHC6348_n4270 (.O(FE_PHN6348_n4270), 
	.I(FE_PHN3364_n4270));
   BUFCKEHD FE_PHC6347_n2703 (.O(FE_PHN6347_n2703), 
	.I(FE_PHN4274_n2703));
   BUFCKEHD FE_PHC6346_n966 (.O(FE_PHN6346_n966), 
	.I(FE_PHN4676_n966));
   BUFCHD FE_PHC6345_n4290 (.O(FE_PHN6345_n4290), 
	.I(FE_PHN3674_n4290));
   BUFCKEHD FE_PHC6344_n922 (.O(FE_PHN6344_n922), 
	.I(FE_PHN3633_n922));
   BUFCHD FE_PHC6343_n1016 (.O(FE_PHN6343_n1016), 
	.I(FE_PHN3420_n1016));
   BUFCKEHD FE_PHC6342_n2926 (.O(FE_PHN6342_n2926), 
	.I(FE_PHN6973_n2926));
   BUFCHD FE_PHC6341_n3126 (.O(FE_PHN6341_n3126), 
	.I(FE_PHN3761_n3126));
   BUFCHD FE_PHC6340_n3939 (.O(FE_PHN6340_n3939), 
	.I(FE_PHN3303_n3939));
   BUFCHD FE_PHC6339_n3089 (.O(FE_PHN6339_n3089), 
	.I(FE_PHN3485_n3089));
   BUFCKEHD FE_PHC6338_n4356 (.O(FE_PHN6338_n4356), 
	.I(FE_PHN3523_n4356));
   BUFCKEHD FE_PHC6337_n3105 (.O(FE_PHN6337_n3105), 
	.I(FE_PHN3300_n3105));
   BUFCHD FE_PHC6336_n4420 (.O(FE_PHN6336_n4420), 
	.I(FE_PHN3945_n4420));
   BUFCKEHD FE_PHC6335_n1864 (.O(FE_PHN6335_n1864), 
	.I(FE_PHN3760_n1864));
   BUFCKEHD FE_PHC6334_ram_237__7_ (.O(FE_PHN6334_ram_237__7_), 
	.I(FE_PHN3389_ram_237__7_));
   BUFCHD FE_PHC6333_n4286 (.O(FE_PHN6333_n4286), 
	.I(FE_PHN3306_n4286));
   BUFCHD FE_PHC6332_n909 (.O(FE_PHN6332_n909), 
	.I(FE_PHN4440_n909));
   BUFCKEHD FE_PHC6331_n4412 (.O(FE_PHN6331_n4412), 
	.I(FE_PHN3505_n4412));
   BUFEHD FE_PHC6330_n3008 (.O(FE_PHN6330_n3008), 
	.I(FE_PHN3433_n3008));
   BUFCHD FE_PHC6329_n3917 (.O(FE_PHN6329_n3917), 
	.I(FE_PHN3564_n3917));
   BUFCKEHD FE_PHC6328_n4384 (.O(FE_PHN6328_n4384), 
	.I(FE_PHN3254_n4384));
   BUFCHD FE_PHC6327_n2966 (.O(FE_PHN6327_n2966), 
	.I(FE_PHN3272_n2966));
   BUFCHD FE_PHC6326_n4406 (.O(FE_PHN6326_n4406), 
	.I(FE_PHN3326_n4406));
   BUFCKEHD FE_PHC6325_n4414 (.O(FE_PHN6325_n4414), 
	.I(FE_PHN3536_n4414));
   BUFCHD FE_PHC6324_n4181 (.O(FE_PHN6324_n4181), 
	.I(FE_PHN3678_n4181));
   BUFCHD FE_PHC6323_n3058 (.O(FE_PHN6323_n3058), 
	.I(FE_PHN4599_n3058));
   BUFCKEHD FE_PHC6322_n3223 (.O(FE_PHN6322_n3223), 
	.I(FE_PHN3410_n3223));
   BUFEHD FE_PHC6321_n3127 (.O(FE_PHN6321_n3127), 
	.I(FE_PHN4088_n3127));
   BUFCKEHD FE_PHC6320_n3141 (.O(FE_PHN6320_n3141), 
	.I(FE_PHN3946_n3141));
   BUFEHD FE_PHC6319_ram_158__11_ (.O(FE_PHN6319_ram_158__11_), 
	.I(FE_PHN3374_ram_158__11_));
   BUFCKEHD FE_PHC6318_n4025 (.O(FE_PHN6318_n4025), 
	.I(FE_PHN3655_n4025));
   BUFCHD FE_PHC6317_n3950 (.O(FE_PHN6317_n3950), 
	.I(FE_PHN3591_n3950));
   BUFEHD FE_PHC6316_n843 (.O(FE_PHN6316_n843), 
	.I(FE_PHN3776_n843));
   BUFCHD FE_PHC6315_n4368 (.O(FE_PHN6315_n4368), 
	.I(FE_PHN3923_n4368));
   BUFCKEHD FE_PHC6314_n958 (.O(FE_PHN6314_n958), 
	.I(FE_PHN6885_n958));
   BUFEHD FE_PHC6313_n2898 (.O(FE_PHN6313_n2898), 
	.I(FE_PHN3785_n2898));
   BUFCHD FE_PHC6312_n4218 (.O(FE_PHN6312_n4218), 
	.I(FE_PHN5121_n4218));
   BUFCHD FE_PHC6311_n4171 (.O(FE_PHN6311_n4171), 
	.I(FE_PHN3604_n4171));
   BUFCHD FE_PHC6310_n850 (.O(FE_PHN6310_n850), 
	.I(FE_PHN3890_n850));
   BUFCKEHD FE_PHC6309_n4383 (.O(FE_PHN6309_n4383), 
	.I(FE_PHN3252_n4383));
   BUFCHD FE_PHC6308_n3099 (.O(FE_PHN6308_n3099), 
	.I(FE_PHN6990_n3099));
   BUFCKEHD FE_PHC6307_n1024 (.O(FE_PHN6307_n1024), 
	.I(FE_PHN3885_n1024));
   BUFCKEHD FE_PHC6306_n1002 (.O(FE_PHN6306_n1002), 
	.I(FE_PHN3791_n1002));
   BUFCKEHD FE_PHC6305_n3138 (.O(FE_PHN6305_n3138), 
	.I(FE_PHN3344_n3138));
   BUFCKEHD FE_PHC6304_n4094 (.O(FE_PHN6304_n4094), 
	.I(FE_PHN7003_n4094));
   BUFCHD FE_PHC6303_n4212 (.O(FE_PHN6303_n4212), 
	.I(FE_PHN3540_n4212));
   BUFCKEHD FE_PHC6302_n4283 (.O(FE_PHN6302_n4283), 
	.I(FE_PHN3825_n4283));
   BUFCKEHD FE_PHC6301_n3015 (.O(FE_PHN6301_n3015), 
	.I(FE_PHN3830_n3015));
   BUFCHD FE_PHC6300_n3918 (.O(FE_PHN6300_n3918), 
	.I(FE_PHN6987_n3918));
   BUFCKEHD FE_PHC6299_n1000 (.O(FE_PHN6299_n1000), 
	.I(FE_PHN3984_n1000));
   BUFCHD FE_PHC6298_n3114 (.O(FE_PHN6298_n3114), 
	.I(FE_PHN3973_n3114));
   BUFCHD FE_PHC6297_n4364 (.O(FE_PHN6297_n4364), 
	.I(FE_PHN3548_n4364));
   BUFEHD FE_PHC6296_n934 (.O(FE_PHN6296_n934), 
	.I(FE_PHN4283_n934));
   BUFCHD FE_PHC6295_n4103 (.O(FE_PHN6295_n4103), 
	.I(FE_PHN4295_n4103));
   BUFCKEHD FE_PHC6294_n4023 (.O(FE_PHN6294_n4023), 
	.I(FE_PHN3446_n4023));
   BUFCKEHD FE_PHC6293_n1029 (.O(FE_PHN6293_n1029), 
	.I(FE_PHN3727_n1029));
   BUFCKEHD FE_PHC6292_n4166 (.O(FE_PHN6292_n4166), 
	.I(FE_PHN6870_n4166));
   BUFCKEHD FE_PHC6291_n3026 (.O(FE_PHN6291_n3026), 
	.I(FE_PHN3779_n3026));
   BUFCHD FE_PHC6290_n3120 (.O(FE_PHN6290_n3120), 
	.I(FE_PHN3416_n3120));
   BUFCKEHD FE_PHC6289_n4185 (.O(FE_PHN6289_n4185), 
	.I(FE_PHN6871_n4185));
   BUFGHD FE_PHC6288_n895 (.O(FE_PHN6288_n895), 
	.I(FE_PHN3884_n895));
   BUFCHD FE_PHC6287_n847 (.O(FE_PHN6287_n847), 
	.I(FE_PHN3636_n847));
   BUFCKEHD FE_PHC6286_n4398 (.O(FE_PHN6286_n4398), 
	.I(n4398));
   BUFCHD FE_PHC6285_n1062 (.O(FE_PHN6285_n1062), 
	.I(n1062));
   BUFCHD FE_PHC6284_n4396 (.O(FE_PHN6284_n4396), 
	.I(FE_PHN3457_n4396));
   BUFCHD FE_PHC6283_n4373 (.O(FE_PHN6283_n4373), 
	.I(FE_PHN3912_n4373));
   BUFCHD FE_PHC6282_n2413 (.O(FE_PHN6282_n2413), 
	.I(FE_PHN6940_n2413));
   BUFCKEHD FE_PHC6281_n997 (.O(FE_PHN6281_n997), 
	.I(FE_PHN3568_n997));
   BUFCHD FE_PHC6280_n3946 (.O(FE_PHN6280_n3946), 
	.I(FE_PHN3860_n3946));
   BUFCHD FE_PHC6279_n986 (.O(FE_PHN6279_n986), 
	.I(FE_PHN3907_n986));
   BUFCHD FE_PHC6278_n886 (.O(FE_PHN6278_n886), 
	.I(FE_PHN3926_n886));
   BUFCHD FE_PHC6277_n4372 (.O(FE_PHN6277_n4372), 
	.I(FE_PHN3384_n4372));
   BUFCHD FE_PHC6276_n869 (.O(FE_PHN6276_n869), 
	.I(FE_PHN4553_n869));
   BUFCHD FE_PHC6275_n4245 (.O(FE_PHN6275_n4245), 
	.I(FE_PHN7008_n4245));
   BUFCKEHD FE_PHC6274_n960 (.O(FE_PHN6274_n960), 
	.I(FE_PHN3365_n960));
   BUFCKEHD FE_PHC6273_n3095 (.O(FE_PHN6273_n3095), 
	.I(FE_PHN3562_n3095));
   BUFCHD FE_PHC6272_n4269 (.O(FE_PHN6272_n4269), 
	.I(FE_PHN6972_n4269));
   BUFCHD FE_PHC6271_n978 (.O(FE_PHN6271_n978), 
	.I(FE_PHN3734_n978));
   BUFCHD FE_PHC6270_n4134 (.O(FE_PHN6270_n4134), 
	.I(FE_PHN6991_n4134));
   BUFCHD FE_PHC6269_ram_31__2_ (.O(FE_PHN6269_ram_31__2_), 
	.I(FE_PHN4414_ram_31__2_));
   BUFCHD FE_PHC6268_ram_145__1_ (.O(FE_PHN6268_ram_145__1_), 
	.I(FE_PHN4134_ram_145__1_));
   BUFCKEHD FE_PHC6267_n1916 (.O(FE_PHN6267_n1916), 
	.I(FE_PHN3817_n1916));
   BUFCHD FE_PHC6266_n3012 (.O(FE_PHN6266_n3012), 
	.I(FE_PHN3740_n3012));
   BUFCKEHD FE_PHC6265_n1921 (.O(FE_PHN6265_n1921), 
	.I(FE_PHN3869_n1921));
   BUFCHD FE_PHC6264_n3042 (.O(FE_PHN6264_n3042), 
	.I(FE_PHN3758_n3042));
   BUFCHD FE_PHC6263_n3032 (.O(FE_PHN6263_n3032), 
	.I(FE_PHN4029_n3032));
   BUFCHD FE_PHC6262_n854 (.O(FE_PHN6262_n854), 
	.I(FE_PHN3295_n854));
   BUFCHD FE_PHC6261_n3133 (.O(FE_PHN6261_n3133), 
	.I(FE_PHN3637_n3133));
   BUFCHD FE_PHC6260_n4097 (.O(FE_PHN6260_n4097), 
	.I(FE_PHN3950_n4097));
   BUFCHD FE_PHC6259_n3062 (.O(FE_PHN6259_n3062), 
	.I(FE_PHN3807_n3062));
   BUFCHD FE_PHC6258_n2986 (.O(FE_PHN6258_n2986), 
	.I(FE_PHN3843_n2986));
   BUFCKEHD FE_PHC6257_n3262 (.O(FE_PHN6257_n3262), 
	.I(FE_PHN3835_n3262));
   BUFCKEHD FE_PHC6256_n849 (.O(FE_PHN6256_n849), 
	.I(FE_PHN3555_n849));
   BUFCHD FE_PHC6255_n3035 (.O(FE_PHN6255_n3035), 
	.I(FE_PHN4042_n3035));
   BUFCHD FE_PHC6254_n1008 (.O(FE_PHN6254_n1008), 
	.I(FE_PHN3393_n1008));
   BUFCHD FE_PHC6253_n2982 (.O(FE_PHN6253_n2982), 
	.I(FE_PHN3733_n2982));
   BUFCHD FE_PHC6252_n2297 (.O(FE_PHN6252_n2297), 
	.I(FE_PHN5296_n2297));
   BUFEHD FE_PHC6251_n3922 (.O(FE_PHN6251_n3922), 
	.I(FE_PHN4028_n3922));
   BUFEHD FE_PHC6250_n3100 (.O(FE_PHN6250_n3100), 
	.I(FE_PHN4041_n3100));
   BUFCHD FE_PHC6249_n4003 (.O(FE_PHN6249_n4003), 
	.I(FE_PHN6956_n4003));
   BUFEHD FE_PHC6248_ram_221__1_ (.O(FE_PHN6248_ram_221__1_), 
	.I(FE_PHN4105_ram_221__1_));
   BUFEHD FE_PHC6247_n4339 (.O(FE_PHN6247_n4339), 
	.I(FE_PHN6962_n4339));
   BUFCHD FE_PHC6246_n993 (.O(FE_PHN6246_n993), 
	.I(FE_PHN3409_n993));
   BUFCKEHD FE_PHC6245_n947 (.O(FE_PHN6245_n947), 
	.I(FE_PHN3767_n947));
   BUFCHD FE_PHC6244_n3084 (.O(FE_PHN6244_n3084), 
	.I(FE_PHN6965_n3084));
   BUFCKIHD FE_PHC6243_n4233 (.O(FE_PHN6243_n4233), 
	.I(FE_PHN6947_n4233));
   BUFCHD FE_PHC6242_n2952 (.O(FE_PHN6242_n2952), 
	.I(FE_PHN3980_n2952));
   BUFCKEHD FE_PHC6241_n919 (.O(FE_PHN6241_n919), 
	.I(FE_PHN6942_n919));
   BUFCHD FE_PHC6240_n3080 (.O(FE_PHN6240_n3080), 
	.I(FE_PHN3954_n3080));
   BUFCHD FE_PHC6239_n3054 (.O(FE_PHN6239_n3054), 
	.I(FE_PHN3849_n3054));
   BUFCHD FE_PHC6238_n3094 (.O(FE_PHN6238_n3094), 
	.I(FE_PHN3324_n3094));
   BUFCKEHD FE_PHC6237_n897 (.O(FE_PHN6237_n897), 
	.I(FE_PHN3533_n897));
   BUFCHD FE_PHC6236_n3014 (.O(FE_PHN6236_n3014), 
	.I(FE_PHN3301_n3014));
   BUFEHD FE_PHC6235_n845 (.O(FE_PHN6235_n845), 
	.I(FE_PHN4330_n845));
   BUFCHD FE_PHC6234_n1005 (.O(FE_PHN6234_n1005), 
	.I(FE_PHN4073_n1005));
   BUFCHD FE_PHC6233_n3130 (.O(FE_PHN6233_n3130), 
	.I(FE_PHN3991_n3130));
   BUFCHD FE_PHC6232_n3125 (.O(FE_PHN6232_n3125), 
	.I(FE_PHN3247_n3125));
   BUFCHD FE_PHC6231_n1042 (.O(FE_PHN6231_n1042), 
	.I(FE_PHN4625_n1042));
   BUFEHD FE_PHC6230_n4167 (.O(FE_PHN6230_n4167), 
	.I(FE_PHN3288_n4167));
   BUFCHD FE_PHC6229_n3110 (.O(FE_PHN6229_n3110), 
	.I(FE_PHN4231_n3110));
   BUFCHD FE_PHC6228_n3092 (.O(FE_PHN6228_n3092), 
	.I(FE_PHN3312_n3092));
   BUFCKEHD FE_PHC6227_n3063 (.O(FE_PHN6227_n3063), 
	.I(FE_PHN6876_n3063));
   BUFEHD FE_PHC6226_n3078 (.O(FE_PHN6226_n3078), 
	.I(FE_PHN7014_n3078));
   BUFCHD FE_PHC6225_n3108 (.O(FE_PHN6225_n3108), 
	.I(FE_PHN6977_n3108));
   BUFCKEHD FE_PHC6224_n4289 (.O(FE_PHN6224_n4289), 
	.I(FE_PHN3975_n4289));
   BUFCHD FE_PHC6223_n4235 (.O(FE_PHN6223_n4235), 
	.I(FE_PHN3369_n4235));
   BUFCKEHD FE_PHC6222_n4199 (.O(FE_PHN6222_n4199), 
	.I(FE_PHN3414_n4199));
   BUFCHD FE_PHC6221_n2258 (.O(FE_PHN6221_n2258), 
	.I(FE_PHN6843_n2258));
   BUFCKEHD FE_PHC6220_n3104 (.O(FE_PHN6220_n3104), 
	.I(n3104));
   BUFCKGHD FE_PHC6219_ram_20__10_ (.O(FE_PHN6219_ram_20__10_), 
	.I(FE_PHN3924_ram_20__10_));
   BUFCHD FE_PHC6218_n3102 (.O(FE_PHN6218_n3102), 
	.I(FE_PHN4101_n3102));
   BUFCKEHD FE_PHC6217_n3124 (.O(FE_PHN6217_n3124), 
	.I(FE_PHN3339_n3124));
   BUFCHD FE_PHC6216_n4238 (.O(FE_PHN6216_n4238), 
	.I(FE_PHN7007_n4238));
   BUFCKEHD FE_PHC6215_n4397 (.O(FE_PHN6215_n4397), 
	.I(FE_PHN3848_n4397));
   BUFCKEHD FE_PHC6214_n1018 (.O(FE_PHN6214_n1018), 
	.I(FE_PHN4566_n1018));
   BUFCHD FE_PHC6213_n2896 (.O(FE_PHN6213_n2896), 
	.I(FE_PHN7009_n2896));
   BUFCHD FE_PHC6212_ram_238__0_ (.O(FE_PHN6212_ram_238__0_), 
	.I(FE_PHN3854_ram_238__0_));
   BUFCHD FE_PHC6211_n3001 (.O(FE_PHN6211_n3001), 
	.I(FE_PHN4059_n3001));
   BUFCKEHD FE_PHC6210_n903 (.O(FE_PHN6210_n903), 
	.I(FE_PHN3726_n903));
   BUFCHD FE_PHC6209_n2886 (.O(FE_PHN6209_n2886), 
	.I(FE_PHN3426_n2886));
   BUFCHD FE_PHC6208_n4327 (.O(FE_PHN6208_n4327), 
	.I(FE_PHN6867_n4327));
   BUFCHD FE_PHC6207_n4388 (.O(FE_PHN6207_n4388), 
	.I(FE_PHN4056_n4388));
   BUFCHD FE_PHC6206_n4076 (.O(FE_PHN6206_n4076), 
	.I(FE_PHN6934_n4076));
   BUFCHD FE_PHC6205_n2158 (.O(FE_PHN6205_n2158), 
	.I(FE_PHN6888_n2158));
   BUFCHD FE_PHC6204_n838 (.O(FE_PHN6204_n838), 
	.I(FE_PHN3366_n838));
   BUFCHD FE_PHC6203_n1068 (.O(FE_PHN6203_n1068), 
	.I(FE_PHN6986_n1068));
   BUFCKEHD FE_PHC6202_n4179 (.O(FE_PHN6202_n4179), 
	.I(FE_PHN5382_n4179));
   BUFCHD FE_PHC6201_n2753 (.O(FE_PHN6201_n2753), 
	.I(FE_PHN5311_n2753));
   BUFCHD FE_PHC6200_n4026 (.O(FE_PHN6200_n4026), 
	.I(FE_PHN3443_n4026));
   BUFCHD FE_PHC6199_n4329 (.O(FE_PHN6199_n4329), 
	.I(FE_PHN3645_n4329));
   BUFGHD FE_PHC6198_n882 (.O(FE_PHN6198_n882), 
	.I(FE_PHN7017_n882));
   BUFCHD FE_PHC6197_n2959 (.O(FE_PHN6197_n2959), 
	.I(FE_PHN3978_n2959));
   BUFCHD FE_PHC6196_n3079 (.O(FE_PHN6196_n3079), 
	.I(FE_PHN6943_n3079));
   BUFCHD FE_PHC6195_n844 (.O(FE_PHN6195_n844), 
	.I(FE_PHN7025_n844));
   BUFCHD FE_PHC6194_n3940 (.O(FE_PHN6194_n3940), 
	.I(FE_PHN6983_n3940));
   BUFCHD FE_PHC6193_n2928 (.O(FE_PHN6193_n2928), 
	.I(FE_PHN7016_n2928));
   BUFGHD FE_PHC6192_n3952 (.O(FE_PHN6192_n3952), 
	.I(FE_PHN6937_n3952));
   BUFCHD FE_PHC6191_n4230 (.O(FE_PHN6191_n4230), 
	.I(FE_PHN4035_n4230));
   BUFCKEHD FE_PHC6190_n4333 (.O(FE_PHN6190_n4333), 
	.I(FE_PHN6978_n4333));
   BUFCKEHD FE_PHC6189_n3074 (.O(FE_PHN6189_n3074), 
	.I(FE_PHN3866_n3074));
   BUFCHD FE_PHC6188_n3936 (.O(FE_PHN6188_n3936), 
	.I(FE_PHN6907_n3936));
   BUFEHD FE_PHC6187_n3914 (.O(FE_PHN6187_n3914), 
	.I(FE_PHN4036_n3914));
   BUFCKEHD FE_PHC6186_n3985 (.O(FE_PHN6186_n3985), 
	.I(FE_PHN3243_n3985));
   BUFCHD FE_PHC6185_n918 (.O(FE_PHN6185_n918), 
	.I(FE_PHN4033_n918));
   BUFCKEHD FE_PHC6184_n2933 (.O(FE_PHN6184_n2933), 
	.I(FE_PHN6967_n2933));
   BUFCHD FE_PHC6183_n3122 (.O(FE_PHN6183_n3122), 
	.I(FE_PHN3958_n3122));
   BUFCHD FE_PHC6182_n3136 (.O(FE_PHN6182_n3136), 
	.I(FE_PHN3712_n3136));
   BUFCHD FE_PHC6181_n3974 (.O(FE_PHN6181_n3974), 
	.I(FE_PHN3271_n3974));
   BUFCHD FE_PHC6180_n3989 (.O(FE_PHN6180_n3989), 
	.I(FE_PHN3751_n3989));
   BUFCHD FE_PHC6179_n3003 (.O(FE_PHN6179_n3003), 
	.I(FE_PHN3614_n3003));
   BUFCHD FE_PHC6178_n982 (.O(FE_PHN6178_n982), 
	.I(FE_PHN3511_n982));
   BUFCHD FE_PHC6177_n2127 (.O(FE_PHN6177_n2127), 
	.I(FE_PHN6828_n2127));
   BUFCHD FE_PHC6176_n4416 (.O(FE_PHN6176_n4416), 
	.I(FE_PHN4007_n4416));
   BUFCKEHD FE_PHC6175_n1064 (.O(FE_PHN6175_n1064), 
	.I(FE_PHN3250_n1064));
   BUFCHD FE_PHC6174_n2993 (.O(FE_PHN6174_n2993), 
	.I(FE_PHN3895_n2993));
   BUFCHD FE_PHC6173_n3096 (.O(FE_PHN6173_n3096), 
	.I(FE_PHN4020_n3096));
   BUFCHD FE_PHC6172_n3951 (.O(FE_PHN6172_n3951), 
	.I(FE_PHN6898_n3951));
   BUFCKEHD FE_PHC6171_n2965 (.O(FE_PHN6171_n2965), 
	.I(FE_PHN3904_n2965));
   BUFCHD FE_PHC6170_n2396 (.O(FE_PHN6170_n2396), 
	.I(FE_PHN6839_n2396));
   BUFCHD FE_PHC6169_n4408 (.O(FE_PHN6169_n4408), 
	.I(FE_PHN3377_n4408));
   BUFCHD FE_PHC6168_n3954 (.O(FE_PHN6168_n3954), 
	.I(FE_PHN6912_n3954));
   BUFCKIHD FE_PHC6167_n4228 (.O(FE_PHN6167_n4228), 
	.I(FE_PHN3594_n4228));
   BUFCKEHD FE_PHC6166_n4417 (.O(FE_PHN6166_n4417), 
	.I(FE_PHN3394_n4417));
   BUFCHD FE_PHC6165_ram_214__13_ (.O(FE_PHN6165_ram_214__13_), 
	.I(FE_PHN6976_ram_214__13_));
   BUFCHD FE_PHC6164_n3006 (.O(FE_PHN6164_n3006), 
	.I(FE_PHN3671_n3006));
   BUFCKEHD FE_PHC6163_n4196 (.O(FE_PHN6163_n4196), 
	.I(FE_PHN7002_n4196));
   BUFCHD FE_PHC6162_n865 (.O(FE_PHN6162_n865), 
	.I(FE_PHN3308_n865));
   BUFCHD FE_PHC6161_n3013 (.O(FE_PHN6161_n3013), 
	.I(FE_PHN3669_n3013));
   BUFEHD FE_PHC6160_n4239 (.O(FE_PHN6160_n4239), 
	.I(FE_PHN6900_n4239));
   BUFCHD FE_PHC6159_n2973 (.O(FE_PHN6159_n2973), 
	.I(FE_PHN3320_n2973));
   BUFCHD FE_PHC6158_n1088 (.O(FE_PHN6158_n1088), 
	.I(FE_PHN3695_n1088));
   BUFCHD FE_PHC6157_n3942 (.O(FE_PHN6157_n3942), 
	.I(FE_PHN3799_n3942));
   BUFCHD FE_PHC6156_n1899 (.O(FE_PHN6156_n1899), 
	.I(FE_PHN6905_n1899));
   BUFCHD FE_PHC6155_n3019 (.O(FE_PHN6155_n3019), 
	.I(FE_PHN3787_n3019));
   BUFCHD FE_PHC6154_n3088 (.O(FE_PHN6154_n3088), 
	.I(FE_PHN3656_n3088));
   BUFCKEHD FE_PHC6153_n3961 (.O(FE_PHN6153_n3961), 
	.I(FE_PHN3307_n3961));
   BUFCKEHD FE_PHC6152_n3086 (.O(FE_PHN6152_n3086), 
	.I(FE_PHN3642_n3086));
   BUFCHD FE_PHC6151_n2991 (.O(FE_PHN6151_n2991), 
	.I(FE_PHN3737_n2991));
   BUFCHD FE_PHC6150_n2920 (.O(FE_PHN6150_n2920), 
	.I(FE_PHN3387_n2920));
   BUFCHD FE_PHC6149_n992 (.O(FE_PHN6149_n992), 
	.I(FE_PHN4285_n992));
   BUFCHD FE_PHC6148_n4281 (.O(FE_PHN6148_n4281), 
	.I(FE_PHN6996_n4281));
   BUFCHD FE_PHC6147_n2969 (.O(FE_PHN6147_n2969), 
	.I(FE_PHN3756_n2969));
   BUFCKEHD FE_PHC6146_n4271 (.O(FE_PHN6146_n4271), 
	.I(FE_PHN6963_n4271));
   BUFCHD FE_PHC6145_n969 (.O(FE_PHN6145_n969), 
	.I(FE_PHN6988_n969));
   BUFCHD FE_PHC6144_n874 (.O(FE_PHN6144_n874), 
	.I(FE_PHN3557_n874));
   BUFCHD FE_PHC6143_n2918 (.O(FE_PHN6143_n2918), 
	.I(FE_PHN3424_n2918));
   BUFCHD FE_PHC6142_n4415 (.O(FE_PHN6142_n4415), 
	.I(FE_PHN4536_n4415));
   BUFCHD FE_PHC6141_n3070 (.O(FE_PHN6141_n3070), 
	.I(FE_PHN3703_n3070));
   BUFEHD FE_PHC6140_n902 (.O(FE_PHN6140_n902), 
	.I(FE_PHN4329_n902));
   BUFCHD FE_PHC6139_n2141 (.O(FE_PHN6139_n2141), 
	.I(FE_PHN6800_n2141));
   BUFCHD FE_PHC6138_n3069 (.O(FE_PHN6138_n3069), 
	.I(FE_PHN5250_n3069));
   BUFCHD FE_PHC6137_n885 (.O(FE_PHN6137_n885), 
	.I(FE_PHN3960_n885));
   BUFCHD FE_PHC6136_n900 (.O(FE_PHN6136_n900), 
	.I(FE_PHN4490_n900));
   BUFCHD FE_PHC6135_n3210 (.O(FE_PHN6135_n3210), 
	.I(FE_PHN3812_n3210));
   BUFCHD FE_PHC6134_n4202 (.O(FE_PHN6134_n4202), 
	.I(FE_PHN6925_n4202));
   BUFCHD FE_PHC6133_n1026 (.O(FE_PHN6133_n1026), 
	.I(FE_PHN3242_n1026));
   BUFCHD FE_PHC6132_n3972 (.O(FE_PHN6132_n3972), 
	.I(FE_PHN6879_n3972));
   BUFCHD FE_PHC6131_n2984 (.O(FE_PHN6131_n2984), 
	.I(FE_PHN3423_n2984));
   BUFCHD FE_PHC6130_n2977 (.O(FE_PHN6130_n2977), 
	.I(FE_PHN3367_n2977));
   BUFCKEHD FE_PHC6129_n3107 (.O(FE_PHN6129_n3107), 
	.I(FE_PHN3275_n3107));
   BUFCHD FE_PHC6128_n3087 (.O(FE_PHN6128_n3087), 
	.I(FE_PHN7010_n3087));
   BUFCKEHD FE_PHC6127_n2979 (.O(FE_PHN6127_n2979), 
	.I(FE_PHN3343_n2979));
   BUFCHD FE_PHC6126_n2934 (.O(FE_PHN6126_n2934), 
	.I(FE_PHN6959_n2934));
   BUFCHD FE_PHC6125_n4394 (.O(FE_PHN6125_n4394), 
	.I(FE_PHN3455_n4394));
   BUFCHD FE_PHC6124_n3009 (.O(FE_PHN6124_n3009), 
	.I(FE_PHN3559_n3009));
   BUFCHD FE_PHC6123_n4380 (.O(FE_PHN6123_n4380), 
	.I(FE_PHN3296_n4380));
   BUFCHD FE_PHC6122_n2997 (.O(FE_PHN6122_n2997), 
	.I(FE_PHN6989_n2997));
   BUFCHD FE_PHC6121_n3050 (.O(FE_PHN6121_n3050), 
	.I(FE_PHN3932_n3050));
   BUFCHD FE_PHC6120_n2980 (.O(FE_PHN6120_n2980), 
	.I(FE_PHN7011_n2980));
   BUFCHD FE_PHC6119_n3921 (.O(FE_PHN6119_n3921), 
	.I(FE_PHN7000_n3921));
   BUFCKEHD FE_PHC6118_n4300 (.O(FE_PHN6118_n4300), 
	.I(FE_PHN4462_n4300));
   BUFCHD FE_PHC6117_n853 (.O(FE_PHN6117_n853), 
	.I(FE_PHN3784_n853));
   BUFCHD FE_PHC6116_n2946 (.O(FE_PHN6116_n2946), 
	.I(FE_PHN6954_n2946));
   BUFCHD FE_PHC6115_ram_229__12_ (.O(FE_PHN6115_ram_229__12_), 
	.I(FE_PHN7018_ram_229__12_));
   BUFCHD FE_PHC6114_n4169 (.O(FE_PHN6114_n4169), 
	.I(FE_PHN6927_n4169));
   BUFCHD FE_PHC6113_n3956 (.O(FE_PHN6113_n3956), 
	.I(FE_PHN6924_n3956));
   BUFCHD FE_PHC6112_n3024 (.O(FE_PHN6112_n3024), 
	.I(FE_PHN6968_n3024));
   BUFCHD FE_PHC6111_n3993 (.O(FE_PHN6111_n3993), 
	.I(FE_PHN4015_n3993));
   BUFCHD FE_PHC6110_n899 (.O(FE_PHN6110_n899), 
	.I(FE_PHN4963_n899));
   BUFCHD FE_PHC6109_n4262 (.O(FE_PHN6109_n4262), 
	.I(FE_PHN7001_n4262));
   BUFCHD FE_PHC6108_n3116 (.O(FE_PHN6108_n3116), 
	.I(FE_PHN6847_n3116));
   BUFCHD FE_PHC6107_n839 (.O(FE_PHN6107_n839), 
	.I(FE_PHN6868_n839));
   BUFCHD FE_PHC6106_n4284 (.O(FE_PHN6106_n4284), 
	.I(FE_PHN3495_n4284));
   BUFCHD FE_PHC6105_n4402 (.O(FE_PHN6105_n4402), 
	.I(FE_PHN3297_n4402));
   BUFCHD FE_PHC6104_n1074 (.O(FE_PHN6104_n1074), 
	.I(FE_PHN3281_n1074));
   BUFCHD FE_PHC6103_n2981 (.O(FE_PHN6103_n2981), 
	.I(FE_PHN3478_n2981));
   BUFCKEHD FE_PHC6102_ram_153__7_ (.O(FE_PHN6102_ram_153__7_), 
	.I(FE_PHN3373_ram_153__7_));
   BUFCKEHD FE_PHC6101_n2621 (.O(FE_PHN6101_n2621), 
	.I(FE_PHN6917_n2621));
   BUFCHD FE_PHC6100_n984 (.O(FE_PHN6100_n984), 
	.I(FE_PHN3546_n984));
   BUFCKEHD FE_PHC6099_n4111 (.O(FE_PHN6099_n4111), 
	.I(FE_PHN6916_n4111));
   BUFCHD FE_PHC6098_n1020 (.O(FE_PHN6098_n1020), 
	.I(FE_PHN6941_n1020));
   BUFCHD FE_PHC6097_n3959 (.O(FE_PHN6097_n3959), 
	.I(FE_PHN6897_n3959));
   BUFCHD FE_PHC6096_n2983 (.O(FE_PHN6096_n2983), 
	.I(FE_PHN3706_n2983));
   BUFCHD FE_PHC6095_n2996 (.O(FE_PHN6095_n2996), 
	.I(FE_PHN3608_n2996));
   BUFCKEHD FE_PHC6094_n3977 (.O(FE_PHN6094_n3977), 
	.I(FE_PHN3986_n3977));
   BUFCHD FE_PHC6093_n4007 (.O(FE_PHN6093_n4007), 
	.I(FE_PHN3661_n4007));
   BUFCKEHD FE_PHC6092_n3103 (.O(FE_PHN6092_n3103), 
	.I(FE_PHN6952_n3103));
   BUFCHD FE_PHC6091_n2944 (.O(FE_PHN6091_n2944), 
	.I(FE_PHN4634_n2944));
   BUFCHD FE_PHC6090_n4022 (.O(FE_PHN6090_n4022), 
	.I(FE_PHN3510_n4022));
   BUFCHD FE_PHC6089_n3975 (.O(FE_PHN6089_n3975), 
	.I(FE_PHN4341_n3975));
   BUFCHD FE_PHC6088_n2954 (.O(FE_PHN6088_n2954), 
	.I(FE_PHN3993_n2954));
   BUFCHD FE_PHC6087_n1009 (.O(FE_PHN6087_n1009), 
	.I(FE_PHN4368_n1009));
   BUFCHD FE_PHC6086_n2975 (.O(FE_PHN6086_n2975), 
	.I(FE_PHN3765_n2975));
   BUFCHD FE_PHC6085_n2888 (.O(FE_PHN6085_n2888), 
	.I(FE_PHN3333_n2888));
   BUFCHD FE_PHC6084_n4291 (.O(FE_PHN6084_n4291), 
	.I(FE_PHN6926_n4291));
   BUFCHD FE_PHC6083_n2916 (.O(FE_PHN6083_n2916), 
	.I(FE_PHN6931_n2916));
   BUFCHD FE_PHC6082_n1032 (.O(FE_PHN6082_n1032), 
	.I(FE_PHN3359_n1032));
   BUFCKEHD FE_PHC6081_n961 (.O(FE_PHN6081_n961), 
	.I(FE_PHN6892_n961));
   BUFCHD FE_PHC6080_n3044 (.O(FE_PHN6080_n3044), 
	.I(FE_PHN3575_n3044));
   BUFCHD FE_PHC6079_n4183 (.O(FE_PHN6079_n4183), 
	.I(FE_PHN6918_n4183));
   BUFCHD FE_PHC6078_n1077 (.O(FE_PHN6078_n1077), 
	.I(FE_PHN3796_n1077));
   BUFCHD FE_PHC6077_n3943 (.O(FE_PHN6077_n3943), 
	.I(FE_PHN6855_n3943));
   BUFCKEHD FE_PHC6076_n4386 (.O(FE_PHN6076_n4386), 
	.I(FE_PHN3292_n4386));
   BUFCHD FE_PHC6075_n3007 (.O(FE_PHN6075_n3007), 
	.I(FE_PHN3730_n3007));
   BUFCHD FE_PHC6074_n4251 (.O(FE_PHN6074_n4251), 
	.I(FE_PHN6994_n4251));
   BUFCHD FE_PHC6073_n3969 (.O(FE_PHN6073_n3969), 
	.I(FE_PHN6985_n3969));
   BUFCHD FE_PHC6072_n4222 (.O(FE_PHN6072_n4222), 
	.I(FE_PHN6932_n4222));
   BUFCHD FE_PHC6071_n4037 (.O(FE_PHN6071_n4037), 
	.I(FE_PHN3804_n4037));
   BUFCHD FE_PHC6070_n970 (.O(FE_PHN6070_n970), 
	.I(FE_PHN3323_n970));
   BUFCHD FE_PHC6069_n3998 (.O(FE_PHN6069_n3998), 
	.I(FE_PHN6896_n3998));
   BUFCHD FE_PHC6068_n3022 (.O(FE_PHN6068_n3022), 
	.I(FE_PHN3398_n3022));
   BUFCHD FE_PHC6067_n3255 (.O(FE_PHN6067_n3255), 
	.I(FE_PHN3968_n3255));
   BUFCHD FE_PHC6066_n3924 (.O(FE_PHN6066_n3924), 
	.I(FE_PHN7023_n3924));
   BUFCHD FE_PHC6065_n2953 (.O(FE_PHN6065_n2953), 
	.I(FE_PHN3663_n2953));
   BUFCHD FE_PHC6064_ram_145__7_ (.O(FE_PHN6064_ram_145__7_), 
	.I(FE_PHN7005_ram_145__7_));
   BUFCHD FE_PHC6063_n4204 (.O(FE_PHN6063_n4204), 
	.I(FE_PHN7022_n4204));
   BUFCKEHD FE_PHC6062_n3081 (.O(FE_PHN6062_n3081), 
	.I(FE_PHN3329_n3081));
   BUFCHD FE_PHC6061_n1072 (.O(FE_PHN6061_n1072), 
	.I(FE_PHN3725_n1072));
   BUFCHD FE_PHC6060_n1048 (.O(FE_PHN6060_n1048), 
	.I(FE_PHN3545_n1048));
   BUFCHD FE_PHC6059_n3112 (.O(FE_PHN6059_n3112), 
	.I(FE_PHN7019_n3112));
   BUFCHD FE_PHC6058_n2950 (.O(FE_PHN6058_n2950), 
	.I(FE_PHN3379_n2950));
   BUFCHD FE_PHC6057_n1896 (.O(FE_PHN6057_n1896), 
	.I(FE_PHN6832_n1896));
   BUFCHD FE_PHC6056_n4006 (.O(FE_PHN6056_n4006), 
	.I(FE_PHN3241_n4006));
   BUFCHD FE_PHC6055_n3996 (.O(FE_PHN6055_n3996), 
	.I(FE_PHN6921_n3996));
   BUFCHD FE_PHC6054_n3067 (.O(FE_PHN6054_n3067), 
	.I(FE_PHN4335_n3067));
   BUFCHD FE_PHC6053_n4260 (.O(FE_PHN6053_n4260), 
	.I(FE_PHN3428_n4260));
   BUFEHD FE_PHC6052_n941 (.O(FE_PHN6052_n941), 
	.I(FE_PHN6829_n941));
   BUFCHD FE_PHC6051_n3098 (.O(FE_PHN6051_n3098), 
	.I(FE_PHN6970_n3098));
   BUFCHD FE_PHC6050_n999 (.O(FE_PHN6050_n999), 
	.I(FE_PHN6999_n999));
   BUFCHD FE_PHC6049_n4279 (.O(FE_PHN6049_n4279), 
	.I(FE_PHN3638_n4279));
   BUFEHD FE_PHC6048_n856 (.O(FE_PHN6048_n856), 
	.I(FE_PHN6805_n856));
   BUFCHD FE_PHC6047_n3982 (.O(FE_PHN6047_n3982), 
	.I(FE_PHN3592_n3982));
   BUFCHD FE_PHC6046_n1025 (.O(FE_PHN6046_n1025), 
	.I(FE_PHN3625_n1025));
   BUFCKJHD FE_PHC6045_n887 (.O(FE_PHN6045_n887), 
	.I(FE_PHN3696_n887));
   BUFCKEHD FE_PHC6044_n1021 (.O(FE_PHN6044_n1021), 
	.I(FE_PHN7020_n1021));
   BUFCHD FE_PHC6043_n3910 (.O(FE_PHN6043_n3910), 
	.I(FE_PHN6936_n3910));
   BUFCKEHD FE_PHC6042_n4203 (.O(FE_PHN6042_n4203), 
	.I(FE_PHN6772_n4203));
   BUFCHD FE_PHC6041_n3134 (.O(FE_PHN6041_n3134), 
	.I(FE_PHN3588_n3134));
   BUFCHD FE_PHC6040_n2943 (.O(FE_PHN6040_n2943), 
	.I(FE_PHN6860_n2943));
   BUFCKEHD FE_PHC6039_n4332 (.O(FE_PHN6039_n4332), 
	.I(FE_PHN3260_n4332));
   BUFCHD FE_PHC6038_n4211 (.O(FE_PHN6038_n4211), 
	.I(FE_PHN6857_n4211));
   BUFCHD FE_PHC6037_n1066 (.O(FE_PHN6037_n1066), 
	.I(FE_PHN6873_n1066));
   BUFCHD FE_PHC6036_n3131 (.O(FE_PHN6036_n3131), 
	.I(FE_PHN7024_n3131));
   BUFCKEHD FE_PHC6035_n1014 (.O(FE_PHN6035_n1014), 
	.I(FE_PHN6748_n1014));
   BUFCHD FE_PHC6034_ram_145__10_ (.O(FE_PHN6034_ram_145__10_), 
	.I(FE_PHN3286_ram_145__10_));
   BUFCHD FE_PHC6033_n3060 (.O(FE_PHN6033_n3060), 
	.I(FE_PHN6923_n3060));
   BUFCHD FE_PHC6032_n998 (.O(FE_PHN6032_n998), 
	.I(FE_PHN4350_n998));
   BUFCHD FE_PHC6031_n890 (.O(FE_PHN6031_n890), 
	.I(FE_PHN6979_n890));
   BUFCHD FE_PHC6030_n989 (.O(FE_PHN6030_n989), 
	.I(FE_PHN6864_n989));
   BUFCHD FE_PHC6029_n1006 (.O(FE_PHN6029_n1006), 
	.I(FE_PHN6974_n1006));
   BUFCHD FE_PHC6028_n3053 (.O(FE_PHN6028_n3053), 
	.I(FE_PHN3350_n3053));
   BUFCHD FE_PHC6027_n889 (.O(FE_PHN6027_n889), 
	.I(FE_PHN6821_n889));
   BUFCHD FE_PHC6026_n4311 (.O(FE_PHN6026_n4311), 
	.I(FE_PHN6904_n4311));
   BUFCHD FE_PHC6025_n4418 (.O(FE_PHN6025_n4418), 
	.I(FE_PHN3479_n4418));
   BUFCHD FE_PHC6024_ram_145__0_ (.O(FE_PHN6024_ram_145__0_), 
	.I(FE_PHN3358_ram_145__0_));
   BUFCHD FE_PHC6023_n892 (.O(FE_PHN6023_n892), 
	.I(FE_PHN6958_n892));
   BUFCKEHD FE_PHC6022_n879 (.O(FE_PHN6022_n879), 
	.I(FE_PHN4480_n879));
   BUFCHD FE_PHC6021_ram_133__9_ (.O(FE_PHN6021_ram_133__9_), 
	.I(FE_PHN6862_ram_133__9_));
   BUFCHD FE_PHC6020_n3076 (.O(FE_PHN6020_n3076), 
	.I(FE_PHN6966_n3076));
   BUFCHD FE_PHC6019_n840 (.O(FE_PHN6019_n840), 
	.I(FE_PHN6895_n840));
   BUFCKEHD FE_PHC6018_n2976 (.O(FE_PHN6018_n2976), 
	.I(FE_PHN3475_n2976));
   BUFCHD FE_PHC6017_n3025 (.O(FE_PHN6017_n3025), 
	.I(FE_PHN6875_n3025));
   BUFCKLHD FE_PHC6016_n884 (.O(FE_PHN6016_n884), 
	.I(FE_PHN6982_n884));
   BUFCHD FE_PHC6015_n4405 (.O(FE_PHN6015_n4405), 
	.I(FE_PHN3355_n4405));
   BUFCHD FE_PHC6014_n3056 (.O(FE_PHN6014_n3056), 
	.I(FE_PHN6992_n3056));
   BUFCHD FE_PHC6013_n4419 (.O(FE_PHN6013_n4419), 
	.I(FE_PHN3473_n4419));
   BUFCHD FE_PHC6012_n2989 (.O(FE_PHN6012_n2989), 
	.I(FE_PHN3653_n2989));
   BUFCHD FE_PHC6011_n846 (.O(FE_PHN6011_n846), 
	.I(FE_PHN6911_n846));
   BUFCHD FE_PHC6010_n3929 (.O(FE_PHN6010_n3929), 
	.I(FE_PHN3244_n3929));
   BUFEHD FE_PHC6009_n4225 (.O(FE_PHN6009_n4225), 
	.I(FE_PHN6784_n4225));
   BUFCHD FE_PHC6008_n2994 (.O(FE_PHN6008_n2994), 
	.I(FE_PHN6971_n2994));
   BUFCHD FE_PHC6007_n4010 (.O(FE_PHN6007_n4010), 
	.I(FE_PHN3251_n4010));
   BUFCHD FE_PHC6006_n881 (.O(FE_PHN6006_n881), 
	.I(FE_PHN3309_n881));
   BUFGHD FE_PHC6005_n2930 (.O(FE_PHN6005_n2930), 
	.I(FE_PHN6838_n2930));
   BUFCHD FE_PHC6004_n4379 (.O(FE_PHN6004_n4379), 
	.I(FE_PHN3280_n4379));
   BUFCHD FE_PHC6003_n4360 (.O(FE_PHN6003_n4360), 
	.I(FE_PHN4479_n4360));
   BUFCHD FE_PHC6002_n1045 (.O(FE_PHN6002_n1045), 
	.I(FE_PHN3405_n1045));
   BUFCHD FE_PHC6001_n3093 (.O(FE_PHN6001_n3093), 
	.I(FE_PHN3421_n3093));
   BUFCHD FE_PHC6000_n893 (.O(FE_PHN6000_n893), 
	.I(FE_PHN3494_n893));
   BUFCHD FE_PHC5999_n848 (.O(FE_PHN5999_n848), 
	.I(FE_PHN6919_n848));
   BUFCHD FE_PHC5998_n3958 (.O(FE_PHN5998_n3958), 
	.I(FE_PHN6964_n3958));
   BUFCHD FE_PHC5997_n870 (.O(FE_PHN5997_n870), 
	.I(FE_PHN7006_n870));
   BUFGHD FE_PHC5996_n866 (.O(FE_PHN5996_n866), 
	.I(FE_PHN6822_n866));
   BUFCHD FE_PHC5995_n4009 (.O(FE_PHN5995_n4009), 
	.I(FE_PHN3634_n4009));
   BUFCHD FE_PHC5994_n1110 (.O(FE_PHN5994_n1110), 
	.I(FE_PHN6960_n1110));
   BUFCHD FE_PHC5993_n2992 (.O(FE_PHN5993_n2992), 
	.I(FE_PHN6938_n2992));
   BUFCKEHD FE_PHC5992_n2995 (.O(FE_PHN5992_n2995), 
	.I(FE_PHN7021_n2995));
   BUFCHD FE_PHC5991_n994 (.O(FE_PHN5991_n994), 
	.I(FE_PHN6910_n994));
   BUFCHD FE_PHC5990_n3976 (.O(FE_PHN5990_n3976), 
	.I(FE_PHN6922_n3976));
   BUFGHD FE_PHC5989_n3023 (.O(FE_PHN5989_n3023), 
	.I(FE_PHN6809_n3023));
   BUFCKGHD FE_PHC5988_n4188 (.O(FE_PHN5988_n4188), 
	.I(FE_PHN6869_n4188));
   BUFCHD FE_PHC5987_n3010 (.O(FE_PHN5987_n3010), 
	.I(FE_PHN3544_n3010));
   BUFCHD FE_PHC5986_ram_153__11_ (.O(FE_PHN5986_ram_153__11_), 
	.I(FE_PHN6945_ram_153__11_));
   BUFCHD FE_PHC5985_n2970 (.O(FE_PHN5985_n2970), 
	.I(FE_PHN7013_n2970));
   BUFCHD FE_PHC5984_n3987 (.O(FE_PHN5984_n3987), 
	.I(FE_PHN6861_n3987));
   BUFCHD FE_PHC5983_n913 (.O(FE_PHN5983_n913), 
	.I(FE_PHN6797_n913));
   BUFCHD FE_PHC5982_n1040 (.O(FE_PHN5982_n1040), 
	.I(FE_PHN3659_n1040));
   BUFCHD FE_PHC5981_n2961 (.O(FE_PHN5981_n2961), 
	.I(FE_PHN3729_n2961));
   BUFCHD FE_PHC5980_n3129 (.O(FE_PHN5980_n3129), 
	.I(FE_PHN6761_n3129));
   BUFCKGHD FE_PHC5979_n3984 (.O(FE_PHN5979_n3984), 
	.I(FE_PHN6903_n3984));
   BUFCHD FE_PHC5978_n3027 (.O(FE_PHN5978_n3027), 
	.I(FE_PHN6887_n3027));
   BUFCHD FE_PHC5977_n2978 (.O(FE_PHN5977_n2978), 
	.I(FE_PHN6955_n2978));
   BUFCKEHD FE_PHC5976_n3018 (.O(FE_PHN5976_n3018), 
	.I(FE_PHN3549_n3018));
   BUFCHD FE_PHC5975_n2374 (.O(FE_PHN5975_n2374), 
	.I(FE_PHN6881_n2374));
   BUFCKEHD FE_PHC5974_n4030 (.O(FE_PHN5974_n4030), 
	.I(FE_PHN3392_n4030));
   BUFCKEHD FE_PHC5973_n2430 (.O(FE_PHN5973_n2430), 
	.I(FE_PHN6804_n2430));
   BUFCHD FE_PHC5972_n876 (.O(FE_PHN5972_n876), 
	.I(FE_PHN6902_n876));
   BUFCKEHD FE_PHC5971_n4401 (.O(FE_PHN5971_n4401), 
	.I(FE_PHN3964_n4401));
   BUFCHD FE_PHC5970_n957 (.O(FE_PHN5970_n957), 
	.I(FE_PHN6939_n957));
   BUFCHD FE_PHC5969_n4172 (.O(FE_PHN5969_n4172), 
	.I(FE_PHN6891_n4172));
   BUFCHD FE_PHC5968_n2897 (.O(FE_PHN5968_n2897), 
	.I(FE_PHN6969_n2897));
   BUFCHD FE_PHC5967_n3916 (.O(FE_PHN5967_n3916), 
	.I(FE_PHN6799_n3916));
   BUFCHD FE_PHC5966_n3128 (.O(FE_PHN5966_n3128), 
	.I(FE_PHN3649_n3128));
   BUFCHD FE_PHC5965_n3978 (.O(FE_PHN5965_n3978), 
	.I(FE_PHN3662_n3978));
   BUFCHD FE_PHC5964_n4195 (.O(FE_PHN5964_n4195), 
	.I(FE_PHN6808_n4195));
   BUFCHD FE_PHC5963_n2998 (.O(FE_PHN5963_n2998), 
	.I(FE_PHN6859_n2998));
   BUFEHD FE_PHC5962_n943 (.O(FE_PHN5962_n943), 
	.I(FE_PHN3783_n943));
   BUFCHD FE_PHC5961_n4217 (.O(FE_PHN5961_n4217), 
	.I(FE_PHN6842_n4217));
   BUFCHD FE_PHC5960_n3075 (.O(FE_PHN5960_n3075), 
	.I(FE_PHN6995_n3075));
   BUFCHD FE_PHC5959_n4389 (.O(FE_PHN5959_n4389), 
	.I(FE_PHN3255_n4389));
   BUFCHD FE_PHC5958_n4355 (.O(FE_PHN5958_n4355), 
	.I(FE_PHN6957_n4355));
   BUFCHD FE_PHC5957_n929 (.O(FE_PHN5957_n929), 
	.I(FE_PHN6791_n929));
   BUFCHD FE_PHC5956_n4340 (.O(FE_PHN5956_n4340), 
	.I(FE_PHN6793_n4340));
   BUFCKIHD FE_PHC5955_n4219 (.O(FE_PHN5955_n4219), 
	.I(n4219));
   BUFGHD FE_PHC5954_n1079 (.O(FE_PHN5954_n1079), 
	.I(FE_PHN6789_n1079));
   BUFCHD FE_PHC5953_n861 (.O(FE_PHN5953_n861), 
	.I(FE_PHN6795_n861));
   BUFCHD FE_PHC5952_n3020 (.O(FE_PHN5952_n3020), 
	.I(FE_PHN3879_n3020));
   BUFCHD FE_PHC5951_n3082 (.O(FE_PHN5951_n3082), 
	.I(FE_PHN3888_n3082));
   BUFCHD FE_PHC5950_n4295 (.O(FE_PHN5950_n4295), 
	.I(FE_PHN6929_n4295));
   BUFCHD FE_PHC5949_n4399 (.O(FE_PHN5949_n4399), 
	.I(FE_PHN3447_n4399));
   BUFCHD FE_PHC5948_n3963 (.O(FE_PHN5948_n3963), 
	.I(FE_PHN6845_n3963));
   BUFCKEHD FE_PHC5947_n1013 (.O(FE_PHN5947_n1013), 
	.I(FE_PHN6719_n1013));
   BUFCHD FE_PHC5946_n3029 (.O(FE_PHN5946_n3029), 
	.I(FE_PHN6851_n3029));
   BUFCHD FE_PHC5945_n4021 (.O(FE_PHN5945_n4021), 
	.I(FE_PHN6915_n4021));
   BUFCHD FE_PHC5944_n4263 (.O(FE_PHN5944_n4263), 
	.I(FE_PHN3302_n4263));
   BUFCHD FE_PHC5943_n3002 (.O(FE_PHN5943_n3002), 
	.I(FE_PHN4419_n3002));
   BUFCHD FE_PHC5942_n2987 (.O(FE_PHN5942_n2987), 
	.I(FE_PHN6948_n2987));
   BUFCHD FE_PHC5941_n3028 (.O(FE_PHN5941_n3028), 
	.I(FE_PHN6755_n3028));
   BUFCHD FE_PHC5940_n4029 (.O(FE_PHN5940_n4029), 
	.I(FE_PHN6813_n4029));
   BUFCHD FE_PHC5939_n3048 (.O(FE_PHN5939_n3048), 
	.I(FE_PHN4085_n3048));
   BUFCHD FE_PHC5938_n4243 (.O(FE_PHN5938_n4243), 
	.I(FE_PHN7012_n4243));
   BUFCHD FE_PHC5937_n4369 (.O(FE_PHN5937_n4369), 
	.I(FE_PHN4334_n4369));
   BUFCHD FE_PHC5936_n2735 (.O(FE_PHN5936_n2735), 
	.I(FE_PHN6906_n2735));
   BUFCHD FE_PHC5935_n4378 (.O(FE_PHN5935_n4378), 
	.I(FE_PHN3456_n4378));
   BUFCHD FE_PHC5934_n4033 (.O(FE_PHN5934_n4033), 
	.I(FE_PHN6886_n4033));
   BUFCHD FE_PHC5933_n911 (.O(FE_PHN5933_n911), 
	.I(FE_PHN6766_n911));
   BUFCHD FE_PHC5932_n4400 (.O(FE_PHN5932_n4400), 
	.I(FE_PHN3828_n4400));
   BUFCHD FE_PHC5931_n2962 (.O(FE_PHN5931_n2962), 
	.I(FE_PHN4075_n2962));
   BUFGHD FE_PHC5930_n3055 (.O(FE_PHN5930_n3055), 
	.I(FE_PHN6796_n3055));
   BUFCHD FE_PHC5929_n4240 (.O(FE_PHN5929_n4240), 
	.I(FE_PHN6775_n4240));
   BUFCHD FE_PHC5928_n4220 (.O(FE_PHN5928_n4220), 
	.I(FE_PHN6824_n4220));
   BUFCHD FE_PHC5927_n4421 (.O(FE_PHN5927_n4421), 
	.I(FE_PHN4125_n4421));
   BUFCHD FE_PHC5926_n975 (.O(FE_PHN5926_n975), 
	.I(FE_PHN6730_n975));
   BUFCHD FE_PHC5925_n1037 (.O(FE_PHN5925_n1037), 
	.I(FE_PHN6817_n1037));
   BUFCHD FE_PHC5924_n2722 (.O(FE_PHN5924_n2722), 
	.I(FE_PHN6830_n2722));
   BUFCHD FE_PHC5923_n3257 (.O(FE_PHN5923_n3257), 
	.I(FE_PHN6872_n3257));
   BUFCHD FE_PHC5922_n3258 (.O(FE_PHN5922_n3258), 
	.I(FE_PHN6764_n3258));
   BUFCHD FE_PHC5921_n3043 (.O(FE_PHN5921_n3043), 
	.I(FE_PHN6841_n3043));
   BUFCHD FE_PHC5920_n864 (.O(FE_PHN5920_n864), 
	.I(FE_PHN6812_n864));
   BUFCKIHD FE_PHC5919_n965 (.O(FE_PHN5919_n965), 
	.I(FE_PHN6831_n965));
   BUFCHD FE_PHC5918_n1090 (.O(FE_PHN5918_n1090), 
	.I(FE_PHN4037_n1090));
   BUFCHD FE_PHC5917_n4028 (.O(FE_PHN5917_n4028), 
	.I(FE_PHN6880_n4028));
   BUFCHD FE_PHC5916_n1030 (.O(FE_PHN5916_n1030), 
	.I(FE_PHN7015_n1030));
   BUFCHD FE_PHC5915_n3964 (.O(FE_PHN5915_n3964), 
	.I(FE_PHN6731_n3964));
   BUFCHD FE_PHC5914_n4324 (.O(FE_PHN5914_n4324), 
	.I(FE_PHN6883_n4324));
   BUFCHD FE_PHC5913_n4361 (.O(FE_PHN5913_n4361), 
	.I(FE_PHN6949_n4361));
   BUFCHD FE_PHC5912_n857 (.O(FE_PHN5912_n857), 
	.I(FE_PHN6846_n857));
   BUFCKIHD FE_PHC5911_n4215 (.O(FE_PHN5911_n4215), 
	.I(FE_PHN6728_n4215));
   BUFCHD FE_PHC5910_n3915 (.O(FE_PHN5910_n3915), 
	.I(FE_PHN6930_n3915));
   BUFCHD FE_PHC5909_n4164 (.O(FE_PHN5909_n4164), 
	.I(FE_PHN6767_n4164));
   BUFCKIHD FE_PHC5908_n4180 (.O(FE_PHN5908_n4180), 
	.I(n4180));
   BUFCHD FE_PHC5907_n4299 (.O(FE_PHN5907_n4299), 
	.I(FE_PHN6803_n4299));
   BUFCHD FE_PHC5906_n910 (.O(FE_PHN5906_n910), 
	.I(FE_PHN6776_n910));
   BUFCHD FE_PHC5905_n3937 (.O(FE_PHN5905_n3937), 
	.I(FE_PHN6865_n3937));
   BUFCHD FE_PHC5904_n2964 (.O(FE_PHN5904_n2964), 
	.I(FE_PHN6717_n2964));
   BUFCHD FE_PHC5903_n2936 (.O(FE_PHN5903_n2936), 
	.I(FE_PHN6909_n2936));
   BUFCHD FE_PHC5902_n855 (.O(FE_PHN5902_n855), 
	.I(FE_PHN6853_n855));
   BUFCHD FE_PHC5901_n3207 (.O(FE_PHN5901_n3207), 
	.I(FE_PHN6837_n3207));
   BUFCHD FE_PHC5900_n1056 (.O(FE_PHN5900_n1056), 
	.I(FE_PHN6877_n1056));
   BUFCHD FE_PHC5899_n3926 (.O(FE_PHN5899_n3926), 
	.I(FE_PHN6993_n3926));
   BUFCHD FE_PHC5898_n4252 (.O(FE_PHN5898_n4252), 
	.I(FE_PHN6894_n4252));
   BUFCHD FE_PHC5897_n2754 (.O(FE_PHN5897_n2754), 
	.I(FE_PHN6811_n2754));
   BUFCHD FE_PHC5896_n4377 (.O(FE_PHN5896_n4377), 
	.I(FE_PHN6856_n4377));
   BUFCHD FE_PHC5895_n1051 (.O(FE_PHN5895_n1051), 
	.I(FE_PHN6852_n1051));
   BUFCHD FE_PHC5894_n2420 (.O(FE_PHN5894_n2420), 
	.I(FE_PHN6754_n2420));
   BUFCHD FE_PHC5893_n4226 (.O(FE_PHN5893_n4226), 
	.I(FE_PHN6854_n4226));
   BUFCHD FE_PHC5892_n4017 (.O(FE_PHN5892_n4017), 
	.I(FE_PHN6882_n4017));
   BUFCHD FE_PHC5891_n925 (.O(FE_PHN5891_n925), 
	.I(FE_PHN6778_n925));
   BUFCHD FE_PHC5890_n3948 (.O(FE_PHN5890_n3948), 
	.I(FE_PHN6889_n3948));
   BUFCHD FE_PHC5889_n3994 (.O(FE_PHN5889_n3994), 
	.I(FE_PHN6961_n3994));
   BUFCHD FE_PHC5888_n3049 (.O(FE_PHN5888_n3049), 
	.I(FE_PHN4357_n3049));
   BUFCHD FE_PHC5887_n4209 (.O(FE_PHN5887_n4209), 
	.I(FE_PHN6787_n4209));
   BUFCHD FE_PHC5886_n2958 (.O(FE_PHN5886_n2958), 
	.I(FE_PHN3762_n2958));
   BUFCHD FE_PHC5885_n4014 (.O(FE_PHN5885_n4014), 
	.I(FE_PHN6798_n4014));
   BUFCHD FE_PHC5884_n935 (.O(FE_PHN5884_n935), 
	.I(FE_PHN6783_n935));
   BUFCHD FE_PHC5883_n858 (.O(FE_PHN5883_n858), 
	.I(FE_PHN6825_n858));
   BUFCHD FE_PHC5882_n905 (.O(FE_PHN5882_n905), 
	.I(FE_PHN6752_n905));
   BUFCHD FE_PHC5881_n2564 (.O(FE_PHN5881_n2564), 
	.I(FE_PHN6756_n2564));
   BUFCHD FE_PHC5880_n2927 (.O(FE_PHN5880_n2927), 
	.I(FE_PHN6779_n2927));
   BUFCKEHD FE_PHC5879_n3052 (.O(FE_PHN5879_n3052), 
	.I(FE_PHN6835_n3052));
   BUFCHD FE_PHC5878_ram_144__8_ (.O(FE_PHN5878_ram_144__8_), 
	.I(FE_PHN6913_ram_144__8_));
   BUFCHD FE_PHC5877_n3992 (.O(FE_PHN5877_n3992), 
	.I(FE_PHN6773_n3992));
   BUFCHD FE_PHC5876_n4307 (.O(FE_PHN5876_n4307), 
	.I(FE_PHN6814_n4307));
   BUFCHD FE_PHC5875_n4385 (.O(FE_PHN5875_n4385), 
	.I(FE_PHN3236_n4385));
   BUFCKKHD FE_PHC5874_n2384 (.O(FE_PHN5874_n2384), 
	.I(FE_PHN3839_n2384));
   BUFCHD FE_PHC5873_n1920 (.O(FE_PHN5873_n1920), 
	.I(FE_PHN6759_n1920));
   BUFCHD FE_PHC5872_n1034 (.O(FE_PHN5872_n1034), 
	.I(FE_PHN6827_n1034));
   BUFCHD FE_PHC5871_n988 (.O(FE_PHN5871_n988), 
	.I(FE_PHN6893_n988));
   BUFCHD FE_PHC5870_n3927 (.O(FE_PHN5870_n3927), 
	.I(FE_PHN6823_n3927));
   BUFCHD FE_PHC5869_n851 (.O(FE_PHN5869_n851), 
	.I(FE_PHN6866_n851));
   BUFCHD FE_PHC5868_n4178 (.O(FE_PHN5868_n4178), 
	.I(FE_PHN6749_n4178));
   BUFCHD FE_PHC5867_n1106 (.O(FE_PHN5867_n1106), 
	.I(FE_PHN6890_n1106));
   BUFCHD FE_PHC5866_n945 (.O(FE_PHN5866_n945), 
	.I(FE_PHN6833_n945));
   BUFCHD FE_PHC5865_n894 (.O(FE_PHN5865_n894), 
	.I(FE_PHN6801_n894));
   BUFCHD FE_PHC5864_n852 (.O(FE_PHN5864_n852), 
	.I(FE_PHN6848_n852));
   BUFCHD FE_PHC5863_n1093 (.O(FE_PHN5863_n1093), 
	.I(FE_PHN6935_n1093));
   BUFCHD FE_PHC5862_n842 (.O(FE_PHN5862_n842), 
	.I(FE_PHN6780_n842));
   BUFCHD FE_PHC5861_n2385 (.O(FE_PHN5861_n2385), 
	.I(FE_PHN6750_n2385));
   BUFCHD FE_PHC5860_n4393 (.O(FE_PHN5860_n4393), 
	.I(FE_PHN6820_n4393));
   BUFCHD FE_PHC5859_n959 (.O(FE_PHN5859_n959), 
	.I(FE_PHN6757_n959));
   BUFCHD FE_PHC5858_n4277 (.O(FE_PHN5858_n4277), 
	.I(FE_PHN6781_n4277));
   BUFCHD FE_PHC5857_n4194 (.O(FE_PHN5857_n4194), 
	.I(FE_PHN6768_n4194));
   BUFCHD FE_PHC5856_n4046 (.O(FE_PHN5856_n4046), 
	.I(FE_PHN6735_n4046));
   BUFCHD FE_PHC5855_n4387 (.O(FE_PHN5855_n4387), 
	.I(FE_PHN6946_n4387));
   BUFCHD FE_PHC5854_n2955 (.O(FE_PHN5854_n2955), 
	.I(FE_PHN3707_n2955));
   BUFCHD FE_PHC5853_n1022 (.O(FE_PHN5853_n1022), 
	.I(FE_PHN6786_n1022));
   BUFCHD FE_PHC5852_n4350 (.O(FE_PHN5852_n4350), 
	.I(FE_PHN6769_n4350));
   BUFCHD FE_PHC5851_n1017 (.O(FE_PHN5851_n1017), 
	.I(FE_PHN6745_n1017));
   BUFCHD FE_PHC5850_n2178 (.O(FE_PHN5850_n2178), 
	.I(FE_PHN6785_n2178));
   BUFCHD FE_PHC5849_n2932 (.O(FE_PHN5849_n2932), 
	.I(FE_PHN6816_n2932));
   BUFCHD FE_PHC5848_n2956 (.O(FE_PHN5848_n2956), 
	.I(FE_PHN3430_n2956));
   BUFCHD FE_PHC5847_n3930 (.O(FE_PHN5847_n3930), 
	.I(FE_PHN6850_n3930));
   BUFCHD FE_PHC5846_n3071 (.O(FE_PHN5846_n3071), 
	.I(FE_PHN6792_n3071));
   BUFCHD FE_PHC5845_n2951 (.O(FE_PHN5845_n2951), 
	.I(FE_PHN3580_n2951));
   BUFCHD FE_PHC5844_n3988 (.O(FE_PHN5844_n3988), 
	.I(FE_PHN6810_n3988));
   BUFCHD FE_PHC5843_n2574 (.O(FE_PHN5843_n2574), 
	.I(FE_PHN6741_n2574));
   BUFCHD FE_PHC5842_n972 (.O(FE_PHN5842_n972), 
	.I(FE_PHN6807_n972));
   BUFCHD FE_PHC5841_n3072 (.O(FE_PHN5841_n3072), 
	.I(FE_PHN6744_n3072));
   BUFCHD FE_PHC5840_n2971 (.O(FE_PHN5840_n2971), 
	.I(FE_PHN6849_n2971));
   BUFCHD FE_PHC5839_n2405 (.O(FE_PHN5839_n2405), 
	.I(FE_PHN6765_n2405));
   BUFCHD FE_PHC5838_n2945 (.O(FE_PHN5838_n2945), 
	.I(FE_PHN6763_n2945));
   BUFCHD FE_PHC5837_n1087 (.O(FE_PHN5837_n1087), 
	.I(FE_PHN6928_n1087));
   BUFCHD FE_PHC5836_n1069 (.O(FE_PHN5836_n1069), 
	.I(FE_PHN6844_n1069));
   BUFCHD FE_PHC5835_n3073 (.O(FE_PHN5835_n3073), 
	.I(FE_PHN6802_n3073));
   BUFCHD FE_PHC5834_n2580 (.O(FE_PHN5834_n2580), 
	.I(FE_PHN6724_n2580));
   BUFCHD FE_PHC5833_n3040 (.O(FE_PHN5833_n3040), 
	.I(FE_PHN6723_n3040));
   BUFCHD FE_PHC5832_n4174 (.O(FE_PHN5832_n4174), 
	.I(FE_PHN6762_n4174));
   BUFCHD FE_PHC5831_n4334 (.O(FE_PHN5831_n4334), 
	.I(FE_PHN6740_n4334));
   BUFCHD FE_PHC5830_n4005 (.O(FE_PHN5830_n4005), 
	.I(FE_PHN6874_n4005));
   BUFCHD FE_PHC5829_n4323 (.O(FE_PHN5829_n4323), 
	.I(FE_PHN6840_n4323));
   BUFCHD FE_PHC5828_n2900 (.O(FE_PHN5828_n2900), 
	.I(FE_PHN6790_n2900));
   BUFCHD FE_PHC5827_n878 (.O(FE_PHN5827_n878), 
	.I(FE_PHN6806_n878));
   BUFCHD FE_PHC5826_n4001 (.O(FE_PHN5826_n4001), 
	.I(FE_PHN6782_n4001));
   BUFCHD FE_PHC5825_n4049 (.O(FE_PHN5825_n4049), 
	.I(FE_PHN6747_n4049));
   BUFCHD FE_PHC5824_n4278 (.O(FE_PHN5824_n4278), 
	.I(FE_PHN6819_n4278));
   BUFCHD FE_PHC5823_n4214 (.O(FE_PHN5823_n4214), 
	.I(FE_PHN6742_n4214));
   BUFCHD FE_PHC5822_n1870 (.O(FE_PHN5822_n1870), 
	.I(FE_PHN6746_n1870));
   BUFCHD FE_PHC5821_n4410 (.O(FE_PHN5821_n4410), 
	.I(FE_PHN6950_n4410));
   BUFCHD FE_PHC5820_n4232 (.O(FE_PHN5820_n4232), 
	.I(FE_PHN6788_n4232));
   BUFCKLHD FE_PHC5819_n2421 (.O(FE_PHN5819_n2421), 
	.I(FE_PHN3298_n2421));
   BUFCHD FE_PHC5818_n4359 (.O(FE_PHN5818_n4359), 
	.I(FE_PHN7004_n4359));
   BUFCHD FE_PHC5817_n4036 (.O(FE_PHN5817_n4036), 
	.I(FE_PHN6818_n4036));
   BUFCHD FE_PHC5816_n2383 (.O(FE_PHN5816_n2383), 
	.I(FE_PHN6774_n2383));
   BUFCHD FE_PHC5815_n4362 (.O(FE_PHN5815_n4362), 
	.I(FE_PHN6953_n4362));
   BUFCKLHD FE_PHC5814_n2437 (.O(FE_PHN5814_n2437), 
	.I(FE_PHN6901_n2437));
   BUFCHD FE_PHC5813_n4407 (.O(FE_PHN5813_n4407), 
	.I(FE_PHN3994_n4407));
   BUFCHD FE_PHC5812_n3919 (.O(FE_PHN5812_n3919), 
	.I(FE_PHN6737_n3919));
   BUFCHD FE_PHC5811_n1082 (.O(FE_PHN5811_n1082), 
	.I(FE_PHN6714_n1082));
   BUFCKKHD FE_PHC5810_n872 (.O(FE_PHN5810_n872), 
	.I(FE_PHN6899_n872));
   BUFCHD FE_PHC5809_n4371 (.O(FE_PHN5809_n4371), 
	.I(FE_PHN6908_n4371));
   BUFCHD FE_PHC5808_n4255 (.O(FE_PHN5808_n4255), 
	.I(FE_PHN6734_n4255));
   BUFCHD FE_PHC5807_n3219 (.O(FE_PHN5807_n3219), 
	.I(FE_PHN6760_n3219));
   BUFCHD FE_PHC5806_n948 (.O(FE_PHN5806_n948), 
	.I(FE_PHN6721_n948));
   BUFCHD FE_PHC5805_n4248 (.O(FE_PHN5805_n4248), 
	.I(FE_PHN6743_n4248));
   BUFCKKHD FE_PHC5804_n2400 (.O(FE_PHN5804_n2400), 
	.I(FE_PHN6777_n2400));
   BUFCHD FE_PHC5803_n1038 (.O(FE_PHN5803_n1038), 
	.I(FE_PHN6771_n1038));
   BUFCHD FE_PHC5802_n3263 (.O(FE_PHN5802_n3263), 
	.I(FE_PHN6733_n3263));
   BUFCKLHD FE_PHC5801_n2399 (.O(FE_PHN5801_n2399), 
	.I(FE_PHN6944_n2399));
   BUFCKLHD FE_PHC5800_n936 (.O(FE_PHN5800_n936), 
	.I(FE_PHN6914_n936));
   BUFCHD FE_PHC5799_n2389 (.O(FE_PHN5799_n2389), 
	.I(FE_PHN6758_n2389));
   BUFCKLHD FE_PHC5798_n2433 (.O(FE_PHN5798_n2433), 
	.I(FE_PHN6836_n2433));
   BUFCKMHD FE_PHC5797_n891 (.O(FE_PHN5797_n891), 
	.I(FE_PHN6997_n891));
   BUFCHD FE_PHC5796_n1078 (.O(FE_PHN5796_n1078), 
	.I(FE_PHN6863_n1078));
   BUFCHD FE_PHC5795_n1905 (.O(FE_PHN5795_n1905), 
	.I(FE_PHN6729_n1905));
   BUFCHD FE_PHC5794_n2599 (.O(FE_PHN5794_n2599), 
	.I(FE_PHN6722_n2599));
   BUFCHD FE_PHC5793_n4343 (.O(FE_PHN5793_n4343), 
	.I(FE_PHN6732_n4343));
   BUFCHD FE_PHC5792_n974 (.O(FE_PHN5792_n974), 
	.I(FE_PHN6713_n974));
   BUFCHD FE_PHC5791_n1902 (.O(FE_PHN5791_n1902), 
	.I(FE_PHN6738_n1902));
   BUFCHD FE_PHC5790_n2408 (.O(FE_PHN5790_n2408), 
	.I(FE_PHN6725_n2408));
   BUFCHD FE_PHC5789_n4000 (.O(FE_PHN5789_n4000), 
	.I(FE_PHN6770_n4000));
   BUFCKMHD FE_PHC5788_n2623 (.O(FE_PHN5788_n2623), 
	.I(FE_PHN6826_n2623));
   BUFCHD FE_PHC5787_n4229 (.O(FE_PHN5787_n4229), 
	.I(FE_PHN6716_n4229));
   BUFCHD FE_PHC5786_n946 (.O(FE_PHN5786_n946), 
	.I(FE_PHN6726_n946));
   BUFCHD FE_PHC5785_n2431 (.O(FE_PHN5785_n2431), 
	.I(FE_PHN6739_n2431));
   BUFCHD FE_PHC5784_n1873 (.O(FE_PHN5784_n1873), 
	.I(FE_PHN6715_n1873));
   BUFCHD FE_PHC5783_n2967 (.O(FE_PHN5783_n2967), 
	.I(FE_PHN6884_n2967));
   BUFCHD FE_PHC5782_n954 (.O(FE_PHN5782_n954), 
	.I(FE_PHN6720_n954));
   BUFCHD FE_PHC5781_n2415 (.O(FE_PHN5781_n2415), 
	.I(FE_PHN6736_n2415));
   BUFCHD FE_PHC5780_n3077 (.O(FE_PHN5780_n3077), 
	.I(FE_PHN6751_n3077));
   BUFCKLHD FE_PHC5779_n920 (.O(FE_PHN5779_n920), 
	.I(FE_PHN6815_n920));
   BUFCKLHD FE_PHC5778_n928 (.O(FE_PHN5778_n928), 
	.I(FE_PHN6753_n928));
   BUFCHD FE_PHC5777_n3068 (.O(FE_PHN5777_n3068), 
	.I(FE_PHN6712_n3068));
   BUFCKEHD FE_PHC5776_n3017 (.O(FE_PHN5776_n3017), 
	.I(FE_PHN6608_n3017));
   BUFCKEHD FE_PHC5775_n2577 (.O(FE_PHN5775_n2577), 
	.I(FE_PHN6604_n2577));
   BUFCKEHD FE_PHC5774_n3033 (.O(FE_PHN5774_n3033), 
	.I(FE_PHN6626_n3033));
   BUFCKEHD FE_PHC5773_n2406 (.O(FE_PHN5773_n2406), 
	.I(FE_PHN6600_n2406));
   BUFCKEHD FE_PHC5772_n3047 (.O(FE_PHN5772_n3047), 
	.I(FE_PHN6602_n3047));
   BUFCKEHD FE_PHC5771_n2414 (.O(FE_PHN5771_n2414), 
	.I(FE_PHN6640_n2414));
   BUFCKEHD FE_PHC5770_n2397 (.O(FE_PHN5770_n2397), 
	.I(FE_PHN6639_n2397));
   BUFCKEHD FE_PHC5769_n2422 (.O(FE_PHN5769_n2422), 
	.I(FE_PHN6606_n2422));
   BUFCKEHD FE_PHC5768_n2938 (.O(FE_PHN5768_n2938), 
	.I(FE_PHN6589_n2938));
   BUFCKEHD FE_PHC5767_n2619 (.O(FE_PHN5767_n2619), 
	.I(FE_PHN6582_n2619));
   BUFCKEHD FE_PHC5766_n2889 (.O(FE_PHN5766_n2889), 
	.I(FE_PHN6586_n2889));
   BUFCKEHD FE_PHC5765_n1913 (.O(FE_PHN5765_n1913), 
	.I(FE_PHN6629_n1913));
   BUFCKEHD FE_PHC5764_n2921 (.O(FE_PHN5764_n2921), 
	.I(FE_PHN6638_n2921));
   BUFCKEHD FE_PHC5763_n4135 (.O(FE_PHN5763_n4135), 
	.I(FE_PHN6628_n4135));
   BUFCHD FE_PHC5762_n1908 (.O(FE_PHN5762_n1908), 
	.I(FE_PHN6619_n1908));
   BUFCKEHD FE_PHC5761_n2697 (.O(FE_PHN5761_n2697), 
	.I(FE_PHN6627_n2697));
   BUFCHD FE_PHC5760_n1375 (.O(FE_PHN5760_n1375), 
	.I(FE_PHN7181_n1375));
   BUFCKEHD FE_PHC5759_n921 (.O(FE_PHN5759_n921), 
	.I(FE_PHN6620_n921));
   BUFCHD FE_PHC5758_n4151 (.O(FE_PHN5758_n4151), 
	.I(FE_PHN6615_n4151));
   BUFCHD FE_PHC5757_n1865 (.O(FE_PHN5757_n1865), 
	.I(FE_PHN7167_n1865));
   BUFCHD FE_PHC5756_n2908 (.O(FE_PHN5756_n2908), 
	.I(FE_PHN7166_n2908));
   BUFCHD FE_PHC5755_n2624 (.O(FE_PHN5755_n2624), 
	.I(FE_PHN6614_n2624));
   BUFCHD FE_PHC5754_n2386 (.O(FE_PHN5754_n2386), 
	.I(FE_PHN7156_n2386));
   BUFCHD FE_PHC5753_n4150 (.O(FE_PHN5753_n4150), 
	.I(FE_PHN6610_n4150));
   BUFCHD FE_PHC5752_n2390 (.O(FE_PHN5752_n2390), 
	.I(FE_PHN7152_n2390));
   BUFCHD FE_PHC5751_n2626 (.O(FE_PHN5751_n2626), 
	.I(FE_PHN6607_n2626));
   BUFCHD FE_PHC5750_n1012 (.O(FE_PHN5750_n1012), 
	.I(FE_PHN6598_n1012));
   BUFCHD FE_PHC5749_n2919 (.O(FE_PHN5749_n2919), 
	.I(FE_PHN6592_n2919));
   BUFCHD FE_PHC5748_n2587 (.O(FE_PHN5748_n2587), 
	.I(FE_PHN6599_n2587));
   BUFCHD FE_PHC5747_n2398 (.O(FE_PHN5747_n2398), 
	.I(FE_PHN6591_n2398));
   BUFCHD FE_PHC5746_n1003 (.O(FE_PHN5746_n1003), 
	.I(FE_PHN6588_n1003));
   BUFCHD FE_PHC5745_n973 (.O(FE_PHN5745_n973), 
	.I(FE_PHN6596_n973));
   BUFCHD FE_PHC5744_n2893 (.O(FE_PHN5744_n2893), 
	.I(FE_PHN6578_n2893));
   BUFJHD FE_PHC5743_n1007 (.O(FE_PHN5743_n1007), 
	.I(FE_PHN6594_n1007));
   BUFCHD FE_PHC5742_n2381 (.O(FE_PHN5742_n2381), 
	.I(FE_PHN6571_n2381));
   BUFCHD FE_PHC5741_n2907 (.O(FE_PHN5741_n2907), 
	.I(FE_PHN6573_n2907));
   BUFJHD FE_PHC5740_n981 (.O(FE_PHN5740_n981), 
	.I(n981));
   BUFCHD FE_PHC5739_n1028 (.O(FE_PHN5739_n1028), 
	.I(FE_PHN6583_n1028));
   BUFCHD FE_PHC5738_n2941 (.O(FE_PHN5738_n2941), 
	.I(FE_PHN6569_n2941));
   BUFCHD FE_PHC5737_n2181 (.O(FE_PHN5737_n2181), 
	.I(FE_PHN6560_n2181));
   BUFCHD FE_PHC5736_n2172 (.O(FE_PHN5736_n2172), 
	.I(FE_PHN6551_n2172));
   BUFLHD FE_PHC5735_n3021 (.O(FE_PHN5735_n3021), 
	.I(n3021));
   BUFCHD FE_PHC5734_n2925 (.O(FE_PHN5734_n2925), 
	.I(FE_PHN6570_n2925));
   BUFCHD FE_PHC5733_n983 (.O(FE_PHN5733_n983), 
	.I(FE_PHN6575_n983));
   BUFCHD FE_PHC5732_n4012 (.O(FE_PHN5732_n4012), 
	.I(FE_PHN6563_n4012));
   DELCKHD FE_PHC5731_n1142 (.O(FE_PHN5731_n1142), 
	.I(FE_PHN4871_n1142));
   BUFCHD FE_PHC5730_n2611 (.O(FE_PHN5730_n2611), 
	.I(FE_PHN6544_n2611));
   BUFCHD FE_PHC5729_n1094 (.O(FE_PHN5729_n1094), 
	.I(FE_PHN6557_n1094));
   BUFCHD FE_PHC5728_n2618 (.O(FE_PHN5728_n2618), 
	.I(FE_PHN6536_n2618));
   BUFCHD FE_PHC5727_n2747 (.O(FE_PHN5727_n2747), 
	.I(FE_PHN6539_n2747));
   BUFCHD FE_PHC5726_n985 (.O(FE_PHN5726_n985), 
	.I(FE_PHN6597_n985));
   BUFCHD FE_PHC5725_n977 (.O(FE_PHN5725_n977), 
	.I(FE_PHN6579_n977));
   BUFCHD FE_PHC5724_n2125 (.O(FE_PHN5724_n2125), 
	.I(FE_PHN6550_n2125));
   BUFCHD FE_PHC5723_n1019 (.O(FE_PHN5723_n1019), 
	.I(FE_PHN6562_n1019));
   BUFCHD FE_PHC5722_n2602 (.O(FE_PHN5722_n2602), 
	.I(FE_PHN6528_n2602));
   BUFCHD FE_PHC5721_n2594 (.O(FE_PHN5721_n2594), 
	.I(FE_PHN6538_n2594));
   BUFCHD FE_PHC5720_n2424 (.O(FE_PHN5720_n2424), 
	.I(FE_PHN6535_n2424));
   BUFCHD FE_PHC5719_n2376 (.O(FE_PHN5719_n2376), 
	.I(FE_PHN6524_n2376));
   BUFLHD FE_PHC5718_n2696 (.O(FE_PHN5718_n2696), 
	.I(FE_PHN4923_n2696));
   BUFCHD FE_PHC5717_n1031 (.O(FE_PHN5717_n1031), 
	.I(FE_PHN6558_n1031));
   BUFJHD FE_PHC5716_n996 (.O(FE_PHN5716_n996), 
	.I(n996));
   BUFCHD FE_PHC5715_n2576 (.O(FE_PHN5715_n2576), 
	.I(FE_PHN6523_n2576));
   BUFCHD FE_PHC5714_n2423 (.O(FE_PHN5714_n2423), 
	.I(FE_PHN6522_n2423));
   BUFCHD FE_PHC5713_n3034 (.O(FE_PHN5713_n3034), 
	.I(FE_PHN6621_n3034));
   BUFCKEHD FE_PHC5712_n1001 (.O(FE_PHN5712_n1001), 
	.I(FE_PHN6540_n1001));
   BUFCHD FE_PHC5711_n2251 (.O(FE_PHN5711_n2251), 
	.I(FE_PHN6503_n2251));
   BUFCHD FE_PHC5710_n2148 (.O(FE_PHN5710_n2148), 
	.I(FE_PHN6541_n2148));
   BUFCHD FE_PHC5709_n3981 (.O(FE_PHN5709_n3981), 
	.I(FE_PHN6529_n3981));
   BUFCHD FE_PHC5708_n2695 (.O(FE_PHN5708_n2695), 
	.I(FE_PHN6554_n2695));
   DELBKHD FE_PHC5707_n2740 (.O(FE_PHN5707_n2740), 
	.I(FE_PHN4952_n2740));
   BUFCHD FE_PHC5706_n2380 (.O(FE_PHN5706_n2380), 
	.I(FE_PHN6512_n2380));
   BUFCHD FE_PHC5705_n953 (.O(FE_PHN5705_n953), 
	.I(FE_PHN6517_n953));
   BUFCHD FE_PHC5704_n2412 (.O(FE_PHN5704_n2412), 
	.I(FE_PHN6501_n2412));
   BUFEHD FE_PHC5703_n2156 (.O(FE_PHN5703_n2156), 
	.I(FE_PHN6509_n2156));
   BUFCHD FE_PHC5702_n2572 (.O(FE_PHN5702_n2572), 
	.I(FE_PHN6510_n2572));
   BUFCHD FE_PHC5701_n2615 (.O(FE_PHN5701_n2615), 
	.I(FE_PHN6499_n2615));
   BUFCHD FE_PHC5700_n2622 (.O(FE_PHN5700_n2622), 
	.I(FE_PHN6514_n2622));
   BUFCHD FE_PHC5699_n2138 (.O(FE_PHN5699_n2138), 
	.I(FE_PHN6483_n2138));
   BUFCKMHD FE_PHC5698_n3965 (.O(FE_PHN5698_n3965), 
	.I(FE_PHN6630_n3965));
   BUFCHD FE_PHC5697_n1158 (.O(FE_PHN5697_n1158), 
	.I(FE_PHN7160_n1158));
   BUFCHD FE_PHC5696_n980 (.O(FE_PHN5696_n980), 
	.I(FE_PHN6553_n980));
   BUFCHD FE_PHC5695_n4018 (.O(FE_PHN5695_n4018), 
	.I(FE_PHN6537_n4018));
   BUFCKMHD FE_PHC5694_n2257 (.O(FE_PHN5694_n2257), 
	.I(FE_PHN6616_n2257));
   BUFCHD FE_PHC5693_n1086 (.O(FE_PHN5693_n1086), 
	.I(FE_PHN6572_n1086));
   BUFMHD FE_PHC5692_n2566 (.O(FE_PHN5692_n2566), 
	.I(FE_PHN4915_n2566));
   BUFCKEHD FE_PHC5691_n1178 (.O(FE_PHN5691_n1178), 
	.I(FE_PHN6518_n1178));
   BUFCHD FE_PHC5690_n2124 (.O(FE_PHN5690_n2124), 
	.I(FE_PHN6465_n2124));
   BUFCKMHD FE_PHC5689_n2743 (.O(FE_PHN5689_n2743), 
	.I(FE_PHN6637_n2743));
   BUFCKMHD FE_PHC5688_n3150 (.O(FE_PHN5688_n3150), 
	.I(FE_PHN6603_n3150));
   BUFCKMHD FE_PHC5687_n2589 (.O(FE_PHN5687_n2589), 
	.I(FE_PHN6633_n2589));
   BUFCKMHD FE_PHC5686_n2749 (.O(FE_PHN5686_n2749), 
	.I(FE_PHN6636_n2749));
   BUFCKMHD FE_PHC5685_n2873 (.O(FE_PHN5685_n2873), 
	.I(FE_PHN4913_n2873));
   BUFCHD FE_PHC5684_n2612 (.O(FE_PHN5684_n2612), 
	.I(FE_PHN6471_n2612));
   BUFEHD FE_PHC5683_n1054 (.O(FE_PHN5683_n1054), 
	.I(FE_PHN6534_n1054));
   BUFCKMHD FE_PHC5682_n4158 (.O(FE_PHN5682_n4158), 
	.I(FE_PHN6632_n4158));
   BUFCKMHD FE_PHC5681_n2876 (.O(FE_PHN5681_n2876), 
	.I(FE_PHN6605_n2876));
   BUFCHD FE_PHC5680_n3004 (.O(FE_PHN5680_n3004), 
	.I(FE_PHN6611_n3004));
   BUFCHD FE_PHC5679_n2149 (.O(FE_PHN5679_n2149), 
	.I(FE_PHN6447_n2149));
   BUFCKMHD FE_PHC5678_n2609 (.O(FE_PHN5678_n2609), 
	.I(FE_PHN6625_n2609));
   BUFCKGHD FE_PHC5677_n967 (.O(FE_PHN5677_n967), 
	.I(FE_PHN6547_n967));
   BUFCKEHD FE_PHC5676_n1190 (.O(FE_PHN5676_n1190), 
	.I(FE_PHN6527_n1190));
   BUFCKMHD FE_PHC5675_n4062 (.O(FE_PHN5675_n4062), 
	.I(FE_PHN6631_n4062));
   BUFCKGHD FE_PHC5674_n1154 (.O(FE_PHN5674_n1154), 
	.I(FE_PHN6530_n1154));
   BUFCKMHD FE_PHC5673_n2857 (.O(FE_PHN5673_n2857), 
	.I(FE_PHN6576_n2857));
   BUFCKMHD FE_PHC5672_n2590 (.O(FE_PHN5672_n2590), 
	.I(FE_PHN6580_n2590));
   BUFCKGHD FE_PHC5671_n1015 (.O(FE_PHN5671_n1015), 
	.I(FE_PHN6548_n1015));
   BUFCKMHD FE_PHC5670_n3944 (.O(FE_PHN5670_n3944), 
	.I(FE_PHN6623_n3944));
   BUFCHD FE_PHC5669_n979 (.O(FE_PHN5669_n979), 
	.I(FE_PHN6546_n979));
   BUFCHD FE_PHC5668_n4114 (.O(FE_PHN5668_n4114), 
	.I(FE_PHN7029_n4114));
   BUFCKMHD FE_PHC5667_n2616 (.O(FE_PHN5667_n2616), 
	.I(FE_PHN6577_n2616));
   BUFCKMHD FE_PHC5666_n2177 (.O(FE_PHN5666_n2177), 
	.I(FE_PHN6601_n2177));
   BUFCKMHD FE_PHC5665_n2161 (.O(FE_PHN5665_n2161), 
	.I(FE_PHN6585_n2161));
   BUFCKMHD FE_PHC5664_n2122 (.O(FE_PHN5664_n2122), 
	.I(FE_PHN6635_n2122));
   BUFCKMHD FE_PHC5663_n2750 (.O(FE_PHN5663_n2750), 
	.I(FE_PHN6567_n2750));
   BUFCKMHD FE_PHC5662_n2176 (.O(FE_PHN5662_n2176), 
	.I(FE_PHN6634_n2176));
   BUFCKMHD FE_PHC5661_n2701 (.O(FE_PHN5661_n2701), 
	.I(FE_PHN6595_n2701));
   BUFCKMHD FE_PHC5660_n1286 (.O(FE_PHN5660_n1286), 
	.I(FE_PHN6587_n1286));
   BUFCKEHD FE_PHC5659_n2382 (.O(FE_PHN5659_n2382), 
	.I(FE_PHN6448_n2382));
   BUFCKMHD FE_PHC5658_n2123 (.O(FE_PHN5658_n2123), 
	.I(FE_PHN6622_n2123));
   BUFCKEHD FE_PHC5657_n2121 (.O(FE_PHN5657_n2121), 
	.I(FE_PHN6469_n2121));
   BUFCKMHD FE_PHC5656_n4107 (.O(FE_PHN5656_n4107), 
	.I(FE_PHN6624_n4107));
   BUFCKMHD FE_PHC5655_n2144 (.O(FE_PHN5655_n2144), 
	.I(n2144));
   BUFCKLHD FE_PHC5654_n2375 (.O(FE_PHN5654_n2375), 
	.I(FE_PHN6566_n2375));
   BUFCKEHD FE_PHC5653_n2137 (.O(FE_PHN5653_n2137), 
	.I(FE_PHN6460_n2137));
   BUFCKMHD FE_PHC5652_n2171 (.O(FE_PHN5652_n2171), 
	.I(FE_PHN6590_n2171));
   BUFCKLHD FE_PHC5651_n2407 (.O(FE_PHN5651_n2407), 
	.I(FE_PHN6561_n2407));
   BUFCKLHD FE_PHC5650_n2428 (.O(FE_PHN5650_n2428), 
	.I(FE_PHN6574_n2428));
   BUFCKLHD FE_PHC5649_n2411 (.O(FE_PHN5649_n2411), 
	.I(FE_PHN6549_n2411));
   BUFCKLHD FE_PHC5648_n2429 (.O(FE_PHN5648_n2429), 
	.I(FE_PHN4812_n2429));
   BUFCKGHD FE_PHC5647_n2401 (.O(FE_PHN5647_n2401), 
	.I(FE_PHN6445_n2401));
   BUFCHD FE_PHC5646_n2923 (.O(FE_PHN5646_n2923), 
	.I(FE_PHN3530_n2923));
   BUFCHD FE_PHC5645_n2727 (.O(FE_PHN5645_n2727), 
	.I(FE_PHN3602_n2727));
   BUFCKEHD FE_PHC5644_n1027 (.O(FE_PHN5644_n1027), 
	.I(n1027));
   BUFCHD FE_PHC5643_n2733 (.O(FE_PHN5643_n2733), 
	.I(FE_PHN3702_n2733));
   BUFCHD FE_PHC5642_n2732 (.O(FE_PHN5642_n2732), 
	.I(FE_PHN3777_n2732));
   BUFCKEHD FE_PHC5641_n3132 (.O(FE_PHN5641_n3132), 
	.I(FE_PHN6372_n3132));
   BUFCHD FE_PHC5640_n2605 (.O(FE_PHN5640_n2605), 
	.I(FE_PHN6438_n2605));
   BUFCKEHD FE_PHC5639_n3117 (.O(FE_PHN5639_n3117), 
	.I(FE_PHN6368_n3117));
   BUFCKEHD FE_PHC5638_n4270 (.O(FE_PHN5638_n4270), 
	.I(FE_PHN6348_n4270));
   BUFCKEHD FE_PHC5637_n2262 (.O(FE_PHN5637_n2262), 
	.I(n2262));
   BUFCKEHD FE_PHC5636_n2554 (.O(FE_PHN5636_n2554), 
	.I(FE_PHN6420_n2554));
   BUFCKEHD FE_PHC5635_n4123 (.O(FE_PHN5635_n4123), 
	.I(FE_PHN6434_n4123));
   BUFCKEHD FE_PHC5634_n3913 (.O(FE_PHN5634_n3913), 
	.I(FE_PHN3534_n3913));
   BUFCKEHD FE_PHC5633_n4181 (.O(FE_PHN5633_n4181), 
	.I(FE_PHN6324_n4181));
   BUFEHD FE_PHC5632_n1206 (.O(FE_PHN5632_n1206), 
	.I(FE_PHN3626_n1206));
   BUFCHD FE_PHC5631_n2600 (.O(FE_PHN5631_n2600), 
	.I(FE_PHN6412_n2600));
   BUFCHD FE_PHC5630_n4175 (.O(FE_PHN5630_n4175), 
	.I(FE_PHN6410_n4175));
   BUFCHD FE_PHC5629_n1046 (.O(FE_PHN5629_n1046), 
	.I(FE_PHN3285_n1046));
   BUFEHD FE_PHC5628_n4170 (.O(FE_PHN5628_n4170), 
	.I(FE_PHN3698_n4170));
   BUFCHD FE_PHC5627_n4015 (.O(FE_PHN5627_n4015), 
	.I(FE_PHN3235_n4015));
   BUFCHD FE_PHC5626_n971 (.O(FE_PHN5626_n971), 
	.I(n971));
   BUFCKEHD FE_PHC5625_n3016 (.O(FE_PHN5625_n3016), 
	.I(FE_PHN3886_n3016));
   BUFCKEHD FE_PHC5624_n3095 (.O(FE_PHN5624_n3095), 
	.I(FE_PHN6273_n3095));
   BUFCHD FE_PHC5623_n2391 (.O(FE_PHN5623_n2391), 
	.I(FE_PHN6380_n2391));
   BUFCKEHD FE_PHC5622_n3111 (.O(FE_PHN5622_n3111), 
	.I(FE_PHN6351_n3111));
   BUFCHD FE_PHC5621_n2413 (.O(FE_PHN5621_n2413), 
	.I(FE_PHN6282_n2413));
   BUFEHD FE_PHC5620_n3920 (.O(FE_PHN5620_n3920), 
	.I(FE_PHN3982_n3920));
   BUFCHD FE_PHC5619_n1062 (.O(FE_PHN5619_n1062), 
	.I(FE_PHN6285_n1062));
   BUFCHD FE_PHC5618_n2926 (.O(FE_PHN5618_n2926), 
	.I(FE_PHN6342_n2926));
   BUFCKEHD FE_PHC5617_n4268 (.O(FE_PHN5617_n4268), 
	.I(FE_PHN3953_n4268));
   BUFCKEHD FE_PHC5616_n3066 (.O(FE_PHN5616_n3066), 
	.I(FE_PHN6432_n3066));
   BUFCKEHD FE_PHC5615_n4290 (.O(FE_PHN5615_n4290), 
	.I(FE_PHN6345_n4290));
   BUFCKEHD FE_PHC5614_n3036 (.O(FE_PHN5614_n3036), 
	.I(FE_PHN6418_n3036));
   BUFCHD FE_PHC5613_n2910 (.O(FE_PHN5613_n2910), 
	.I(FE_PHN6413_n2910));
   BUFJHD FE_PHC5612_n3241 (.O(FE_PHN5612_n3241), 
	.I(n3241));
   BUFEHD FE_PHC5611_n4094 (.O(FE_PHN5611_n4094), 
	.I(FE_PHN3913_n4094));
   BUFCKEHD FE_PHC5610_n3911 (.O(FE_PHN5610_n3911), 
	.I(FE_PHN6431_n3911));
   BUFCHD FE_PHC5609_n1068 (.O(FE_PHN5609_n1068), 
	.I(FE_PHN6203_n1068));
   BUFCHD FE_PHC5608_n2258 (.O(FE_PHN5608_n2258), 
	.I(FE_PHN6221_n2258));
   BUFCKEHD FE_PHC5607_n3031 (.O(FE_PHN5607_n3031), 
	.I(FE_PHN6378_n3031));
   BUFCKEHD FE_PHC5606_ram_154__5_ (.O(FE_PHN5606_ram_154__5_), 
	.I(FE_PHN3722_ram_154__5_));
   BUFCHD FE_PHC5605_n2127 (.O(FE_PHN5605_n2127), 
	.I(FE_PHN6177_n2127));
   BUFCHD FE_PHC5604_n2158 (.O(FE_PHN5604_n2158), 
	.I(FE_PHN6205_n2158));
   BUFCHD FE_PHC5603_n2396 (.O(FE_PHN5603_n2396), 
	.I(FE_PHN6170_n2396));
   BUFCKEHD FE_PHC5602_n3083 (.O(FE_PHN5602_n3083), 
	.I(FE_PHN6371_n3083));
   BUFCKEHD FE_PHC5601_n3085 (.O(FE_PHN5601_n3085), 
	.I(FE_PHN6389_n3085));
   BUFCHD FE_PHC5600_n3950 (.O(FE_PHN5600_n3950), 
	.I(FE_PHN6317_n3950));
   BUFCKEHD FE_PHC5599_n4231 (.O(FE_PHN5599_n4231), 
	.I(FE_PHN6363_n4231));
   BUFCHD FE_PHC5598_n4097 (.O(FE_PHN5598_n4097), 
	.I(FE_PHN6260_n4097));
   BUFCHD FE_PHC5597_n2141 (.O(FE_PHN5597_n2141), 
	.I(FE_PHN6139_n2141));
   BUFCKEHD FE_PHC5596_ram_20__10_ (.O(FE_PHN5596_ram_20__10_), 
	.I(FE_PHN6219_ram_20__10_));
   BUFCKEHD FE_PHC5595_n4138 (.O(FE_PHN5595_n4138), 
	.I(FE_PHN6384_n4138));
   BUFCHD FE_PHC5594_n3917 (.O(FE_PHN5594_n3917), 
	.I(FE_PHN6329_n3917));
   BUFCKEHD FE_PHC5593_n4398 (.O(FE_PHN5593_n4398), 
	.I(FE_PHN6286_n4398));
   BUFEHD FE_PHC5592_n2990 (.O(FE_PHN5592_n2990), 
	.I(FE_PHN6359_n2990));
   BUFEHD FE_PHC5591_n4076 (.O(FE_PHN5591_n4076), 
	.I(FE_PHN6206_n4076));
   BUFCKEHD FE_PHC5590_n4292 (.O(FE_PHN5590_n4292), 
	.I(FE_PHN3512_n4292));
   BUFCHD FE_PHC5589_n4267 (.O(FE_PHN5589_n4267), 
	.I(FE_PHN6387_n4267));
   BUFCKEHD FE_PHC5588_n3115 (.O(FE_PHN5588_n3115), 
	.I(FE_PHN6390_n3115));
   BUFCKEHD FE_PHC5587_n4417 (.O(FE_PHN5587_n4417), 
	.I(FE_PHN6166_n4417));
   BUFCHD FE_PHC5586_n4265 (.O(FE_PHN5586_n4265), 
	.I(FE_PHN6414_n4265));
   BUFCKEHD FE_PHC5585_n4261 (.O(FE_PHN5585_n4261), 
	.I(FE_PHN6396_n4261));
   BUFCHD FE_PHC5584_n4168 (.O(FE_PHN5584_n4168), 
	.I(FE_PHN6386_n4168));
   BUFCKEHD FE_PHC5583_n3005 (.O(FE_PHN5583_n3005), 
	.I(FE_PHN6430_n3005));
   BUFCKEHD FE_PHC5582_n3114 (.O(FE_PHN5582_n3114), 
	.I(FE_PHN6298_n3114));
   BUFCKEHD FE_PHC5581_n4397 (.O(FE_PHN5581_n4397), 
	.I(FE_PHN6215_n4397));
   BUFEHD FE_PHC5580_n4235 (.O(FE_PHN5580_n4235), 
	.I(FE_PHN6223_n4235));
   BUFCKEHD FE_PHC5579_n4413 (.O(FE_PHN5579_n4413), 
	.I(FE_PHN3596_n4413));
   BUFCKEHD FE_PHC5578_n3081 (.O(FE_PHN5578_n3081), 
	.I(FE_PHN6062_n3081));
   BUFCHD FE_PHC5577_n3952 (.O(FE_PHN5577_n3952), 
	.I(FE_PHN6192_n3952));
   BUFEHD FE_PHC5576_n3951 (.O(FE_PHN5576_n3951), 
	.I(FE_PHN6172_n3951));
   BUFCKEHD FE_PHC5575_n3120 (.O(FE_PHN5575_n3120), 
	.I(FE_PHN6290_n3120));
   BUFCKEHD FE_PHC5574_n4254 (.O(FE_PHN5574_n4254), 
	.I(FE_PHN6377_n4254));
   BUFCHD FE_PHC5573_n3091 (.O(FE_PHN5573_n3091), 
	.I(FE_PHN6391_n3091));
   BUFCHD FE_PHC5572_n3135 (.O(FE_PHN5572_n3135), 
	.I(FE_PHN6415_n3135));
   BUFCKEHD FE_PHC5571_n3946 (.O(FE_PHN5571_n3946), 
	.I(FE_PHN6280_n3946));
   BUFCHD FE_PHC5570_n871 (.O(FE_PHN5570_n871), 
	.I(FE_PHN6385_n871));
   BUFCKEHD FE_PHC5569_n2999 (.O(FE_PHN5569_n2999), 
	.I(FE_PHN3470_n2999));
   BUFCKEHD FE_PHC5568_n3133 (.O(FE_PHN5568_n3133), 
	.I(FE_PHN6261_n3133));
   BUFCHD FE_PHC5567_n3936 (.O(FE_PHN5567_n3936), 
	.I(FE_PHN6188_n3936));
   DELAKHD FE_PHC5566_n873 (.O(FE_PHN5566_n873), 
	.I(FE_PHN3872_n873));
   BUFCHD FE_PHC5565_n3038 (.O(FE_PHN5565_n3038), 
	.I(FE_PHN6358_n3038));
   BUFCHD FE_PHC5564_n4236 (.O(FE_PHN5564_n4236), 
	.I(FE_PHN6355_n4236));
   BUFCKEHD FE_PHC5563_n4187 (.O(FE_PHN5563_n4187), 
	.I(FE_PHN6392_n4187));
   BUFCKEHD FE_PHC5562_ram_237__7_ (.O(FE_PHN5562_ram_237__7_), 
	.I(FE_PHN6334_ram_237__7_));
   BUFCHD FE_PHC5561_n4382 (.O(FE_PHN5561_n4382), 
	.I(FE_PHN6362_n4382));
   BUFCKEHD FE_PHC5560_n3030 (.O(FE_PHN5560_n3030), 
	.I(FE_PHN6426_n3030));
   BUFCKEHD FE_PHC5559_n884 (.O(FE_PHN5559_n884), 
	.I(FE_PHN6016_n884));
   BUFCKEHD FE_PHC5558_n4227 (.O(FE_PHN5558_n4227), 
	.I(FE_PHN6367_n4227));
   BUFCKEHD FE_PHC5557_n3939 (.O(FE_PHN5557_n3939), 
	.I(FE_PHN6340_n3939));
   BUFCHD FE_PHC5556_n4366 (.O(FE_PHN5556_n4366), 
	.I(FE_PHN6404_n4366));
   BUFCHD FE_PHC5555_n909 (.O(FE_PHN5555_n909), 
	.I(FE_PHN6332_n909));
   BUFCHD FE_PHC5554_n4103 (.O(FE_PHN5554_n4103), 
	.I(FE_PHN6295_n4103));
   BUFCHD FE_PHC5553_n838 (.O(FE_PHN5553_n838), 
	.I(FE_PHN6204_n838));
   BUFCKEHD FE_PHC5552_ram_238__0_ (.O(FE_PHN5552_ram_238__0_), 
	.I(FE_PHN6212_ram_238__0_));
   BUFCKEHD FE_PHC5551_n2969 (.O(FE_PHN5551_n2969), 
	.I(FE_PHN6147_n2969));
   BUFEHD FE_PHC5550_n863 (.O(FE_PHN5550_n863), 
	.I(FE_PHN6381_n863));
   BUFCHD FE_PHC5549_n4213 (.O(FE_PHN5549_n4213), 
	.I(FE_PHN6357_n4213));
   BUFCHD FE_PHC5548_n3062 (.O(FE_PHN5548_n3062), 
	.I(FE_PHN6259_n3062));
   BUFCKEHD FE_PHC5547_n4384 (.O(FE_PHN5547_n4384), 
	.I(FE_PHN6328_n4384));
   BUFCKEHD FE_PHC5546_n4244 (.O(FE_PHN5546_n4244), 
	.I(FE_PHN6433_n4244));
   BUFCHD FE_PHC5545_n3127 (.O(FE_PHN5545_n3127), 
	.I(FE_PHN6321_n3127));
   BUFCHD FE_PHC5544_n3100 (.O(FE_PHN5544_n3100), 
	.I(FE_PHN6250_n3100));
   BUFCKEHD FE_PHC5543_n1899 (.O(FE_PHN5543_n1899), 
	.I(FE_PHN6156_n1899));
   BUFCHD FE_PHC5542_n2957 (.O(FE_PHN5542_n2957), 
	.I(FE_PHN6416_n2957));
   BUFCKEHD FE_PHC5541_n3129 (.O(FE_PHN5541_n3129), 
	.I(FE_PHN5980_n3129));
   BUFEHD FE_PHC5540_n895 (.O(FE_PHN5540_n895), 
	.I(FE_PHN6288_n895));
   BUFCHD FE_PHC5539_n3008 (.O(FE_PHN5539_n3008), 
	.I(FE_PHN6330_n3008));
   BUFCKEHD FE_PHC5538_n3019 (.O(FE_PHN5538_n3019), 
	.I(FE_PHN6155_n3019));
   BUFCHD FE_PHC5537_n934 (.O(FE_PHN5537_n934), 
	.I(FE_PHN6296_n934));
   BUFCHD FE_PHC5536_n4233 (.O(FE_PHN5536_n4233), 
	.I(FE_PHN6243_n4233));
   BUFCHD FE_PHC5535_n4245 (.O(FE_PHN5535_n4245), 
	.I(FE_PHN6275_n4245));
   BUFCHD FE_PHC5534_ram_145__1_ (.O(FE_PHN5534_ram_145__1_), 
	.I(FE_PHN6268_ram_145__1_));
   BUFCKEHD FE_PHC5533_n4003 (.O(FE_PHN5533_n4003), 
	.I(FE_PHN6249_n4003));
   BUFCHD FE_PHC5532_ram_158__11_ (.O(FE_PHN5532_ram_158__11_), 
	.I(FE_PHN6319_ram_158__11_));
   BUFCHD FE_PHC5531_n3940 (.O(FE_PHN5531_n3940), 
	.I(FE_PHN6194_n3940));
   BUFCKEHD FE_PHC5530_n4291 (.O(FE_PHN5530_n4291), 
	.I(FE_PHN6084_n4291));
   BUFCKEHD FE_PHC5529_n3109 (.O(FE_PHN5529_n3109), 
	.I(FE_PHN6435_n3109));
   BUFCKEHD FE_PHC5528_ram_229__3_ (.O(FE_PHN5528_ram_229__3_), 
	.I(FE_PHN3519_ram_229__3_));
   BUFCHD FE_PHC5527_n4269 (.O(FE_PHN5527_n4269), 
	.I(FE_PHN6272_n4269));
   BUFCKEHD FE_PHC5526_ram_229__12_ (.O(FE_PHN5526_ram_229__12_), 
	.I(FE_PHN6115_ram_229__12_));
   BUFCKKHD FE_PHC5525_n2963 (.O(FE_PHN5525_n2963), 
	.I(FE_PHN6388_n2963));
   BUFCHD FE_PHC5524_n4134 (.O(FE_PHN5524_n4134), 
	.I(FE_PHN6270_n4134));
   BUFCHD FE_PHC5523_n3119 (.O(FE_PHN5523_n3119), 
	.I(FE_PHN6428_n3119));
   BUFCHD FE_PHC5522_n3099 (.O(FE_PHN5522_n3099), 
	.I(FE_PHN6308_n3099));
   BUFEHD FE_PHC5521_n3956 (.O(FE_PHN5521_n3956), 
	.I(FE_PHN6113_n3956));
   BUFCKEHD FE_PHC5520_n3003 (.O(FE_PHN5520_n3003), 
	.I(FE_PHN6179_n3003));
   BUFEHD FE_PHC5519_n4262 (.O(FE_PHN5519_n4262), 
	.I(FE_PHN6109_n4262));
   BUFCKEHD FE_PHC5518_n4406 (.O(FE_PHN5518_n4406), 
	.I(FE_PHN6326_n4406));
   BUFCHD FE_PHC5517_n4230 (.O(FE_PHN5517_n4230), 
	.I(FE_PHN6191_n4230));
   BUFCKEHD FE_PHC5516_n2973 (.O(FE_PHN5516_n2973), 
	.I(FE_PHN6159_n2973));
   BUFCHD FE_PHC5515_n4395 (.O(FE_PHN5515_n4395), 
	.I(FE_PHN6370_n4395));
   BUFCHD FE_PHC5514_n918 (.O(FE_PHN5514_n918), 
	.I(FE_PHN6185_n918));
   BUFCHD FE_PHC5513_ram_221__1_ (.O(FE_PHN5513_ram_221__1_), 
	.I(FE_PHN6933_ram_221__1_));
   BUFCKEHD FE_PHC5512_n4367 (.O(FE_PHN5512_n4367), 
	.I(FE_PHN6424_n4367));
   BUFCHD FE_PHC5511_n3080 (.O(FE_PHN5511_n3080), 
	.I(FE_PHN6240_n3080));
   BUFCKIHD FE_PHC5510_n2965 (.O(FE_PHN5510_n2965), 
	.I(FE_PHN6171_n2965));
   BUFCHD FE_PHC5509_n4420 (.O(FE_PHN5509_n4420), 
	.I(FE_PHN6336_n4420));
   BUFCHD FE_PHC5508_n2886 (.O(FE_PHN5508_n2886), 
	.I(FE_PHN6209_n2886));
   BUFCHD FE_PHC5507_n2928 (.O(FE_PHN5507_n2928), 
	.I(FE_PHN6193_n2928));
   BUFCHD FE_PHC5506_n2896 (.O(FE_PHN5506_n2896), 
	.I(FE_PHN6213_n2896));
   BUFCHD FE_PHC5505_n2918 (.O(FE_PHN5505_n2918), 
	.I(FE_PHN6143_n2918));
   BUFCKEHD FE_PHC5504_n4295 (.O(FE_PHN5504_n4295), 
	.I(FE_PHN5950_n4295));
   BUFCHD FE_PHC5503_n3084 (.O(FE_PHN5503_n3084), 
	.I(FE_PHN6244_n3084));
   BUFCHD FE_PHC5502_n3001 (.O(FE_PHN5502_n3001), 
	.I(FE_PHN6211_n3001));
   BUFCKEHD FE_PHC5501_n1896 (.O(FE_PHN5501_n1896), 
	.I(FE_PHN6057_n1896));
   BUFCKEHD FE_PHC5500_n2974 (.O(FE_PHN5500_n2974), 
	.I(FE_PHN6411_n2974));
   BUFCHD FE_PHC5499_n3922 (.O(FE_PHN5499_n3922), 
	.I(FE_PHN6251_n3922));
   BUFCKEHD FE_PHC5498_n3046 (.O(FE_PHN5498_n3046), 
	.I(FE_PHN6402_n3046));
   BUFCHD FE_PHC5497_n3032 (.O(FE_PHN5497_n3032), 
	.I(FE_PHN6263_n3032));
   BUFCHD FE_PHC5496_n4171 (.O(FE_PHN5496_n4171), 
	.I(FE_PHN6311_n4171));
   BUFCHD FE_PHC5495_n4414 (.O(FE_PHN5495_n4414), 
	.I(FE_PHN6325_n4414));
   BUFCHD FE_PHC5494_n845 (.O(FE_PHN5494_n845), 
	.I(FE_PHN6235_n845));
   BUFCHD FE_PHC5493_n3058 (.O(FE_PHN5493_n3058), 
	.I(FE_PHN6323_n3058));
   BUFCHD FE_PHC5492_n4339 (.O(FE_PHN5492_n4339), 
	.I(FE_PHN6247_n4339));
   BUFCHD FE_PHC5491_n3035 (.O(FE_PHN5491_n3035), 
	.I(FE_PHN6255_n3035));
   BUFCHD FE_PHC5490_n1023 (.O(FE_PHN5490_n1023), 
	.I(FE_PHN6405_n1023));
   BUFCHD FE_PHC5489_n854 (.O(FE_PHN5489_n854), 
	.I(FE_PHN6262_n854));
   BUFCHD FE_PHC5488_n4276 (.O(FE_PHN5488_n4276), 
	.I(FE_PHN6366_n4276));
   BUFCHD FE_PHC5487_n3088 (.O(FE_PHN5487_n3088), 
	.I(FE_PHN6154_n3088));
   BUFCHD FE_PHC5486_n3954 (.O(FE_PHN5486_n3954), 
	.I(FE_PHN6168_n3954));
   BUFCHD FE_PHC5485_n2920 (.O(FE_PHN5485_n2920), 
	.I(FE_PHN6150_n2920));
   BUFCHD FE_PHC5484_n4239 (.O(FE_PHN5484_n4239), 
	.I(FE_PHN6160_n4239));
   BUFCHD FE_PHC5483_n843 (.O(FE_PHN5483_n843), 
	.I(FE_PHN6316_n843));
   BUFCHD FE_PHC5482_n3096 (.O(FE_PHN5482_n3096), 
	.I(FE_PHN6173_n3096));
   BUFCHD FE_PHC5481_n3123 (.O(FE_PHN5481_n3123), 
	.I(FE_PHN6409_n3123));
   BUFCKEHD FE_PHC5480_ram_17__14_ (.O(FE_PHN5480_ram_17__14_), 
	.I(FE_PHN6395_ram_17__14_));
   BUFCKEHD FE_PHC5479_n4238 (.O(FE_PHN5479_n4238), 
	.I(FE_PHN6216_n4238));
   BUFCHD FE_PHC5478_n4202 (.O(FE_PHN5478_n4202), 
	.I(FE_PHN6134_n4202));
   BUFCKKHD FE_PHC5477_n968 (.O(FE_PHN5477_n968), 
	.I(FE_PHN6356_n968));
   BUFCHD FE_PHC5476_ram_214__13_ (.O(FE_PHN5476_ram_214__13_), 
	.I(FE_PHN6165_ram_214__13_));
   BUFCHD FE_PHC5475_n3102 (.O(FE_PHN5475_n3102), 
	.I(FE_PHN6218_n3102));
   BUFCHD FE_PHC5474_n3914 (.O(FE_PHN5474_n3914), 
	.I(FE_PHN6878_n3914));
   BUFCHD FE_PHC5473_n3078 (.O(FE_PHN5473_n3078), 
	.I(FE_PHN6226_n3078));
   BUFCHD FE_PHC5472_n2944 (.O(FE_PHN5472_n2944), 
	.I(FE_PHN6091_n2944));
   BUFEHD FE_PHC5471_n1066 (.O(FE_PHN5471_n1066), 
	.I(FE_PHN6037_n1066));
   BUFCKEHD FE_PHC5470_n4195 (.O(FE_PHN5470_n4195), 
	.I(FE_PHN5964_n4195));
   BUFCHD FE_PHC5469_n874 (.O(FE_PHN5469_n874), 
	.I(FE_PHN6144_n874));
   BUFCHD FE_PHC5468_n4388 (.O(FE_PHN5468_n4388), 
	.I(FE_PHN6207_n4388));
   BUFCHD FE_PHC5467_n886 (.O(FE_PHN5467_n886), 
	.I(FE_PHN6278_n886));
   BUFCHD FE_PHC5466_n844 (.O(FE_PHN5466_n844), 
	.I(FE_PHN6195_n844));
   BUFCHD FE_PHC5465_n900 (.O(FE_PHN5465_n900), 
	.I(FE_PHN6136_n900));
   BUFGHD FE_PHC5464_n3044 (.O(FE_PHN5464_n3044), 
	.I(FE_PHN6080_n3044));
   BUFGHD FE_PHC5463_n4228 (.O(FE_PHN5463_n4228), 
	.I(FE_PHN6167_n4228));
   BUFCKKHD FE_PHC5462_n4412 (.O(FE_PHN5462_n4412), 
	.I(FE_PHN6331_n4412));
   BUFCHD FE_PHC5461_n4329 (.O(FE_PHN5461_n4329), 
	.I(FE_PHN6199_n4329));
   BUFCHD FE_PHC5460_n3110 (.O(FE_PHN5460_n3110), 
	.I(FE_PHN6229_n3110));
   BUFCHD FE_PHC5459_n2934 (.O(FE_PHN5459_n2934), 
	.I(FE_PHN6126_n2934));
   BUFCKLHD FE_PHC5458_n4201 (.O(FE_PHN5458_n4201), 
	.I(FE_PHN6379_n4201));
   BUFCHD FE_PHC5457_n2898 (.O(FE_PHN5457_n2898), 
	.I(FE_PHN6313_n2898));
   BUFCKEHD FE_PHC5456_n4219 (.O(FE_PHN5456_n4219), 
	.I(FE_PHN6718_n4219));
   BUFCHD FE_PHC5455_n3139 (.O(FE_PHN5455_n3139), 
	.I(FE_PHN6398_n3139));
   BUFCHD FE_PHC5454_n4169 (.O(FE_PHN5454_n4169), 
	.I(FE_PHN6114_n4169));
   BUFCKEHD FE_PHC5453_n4026 (.O(FE_PHN5453_n4026), 
	.I(FE_PHN6200_n4026));
   BUFCHD FE_PHC5452_n877 (.O(FE_PHN5452_n877), 
	.I(FE_PHN6350_n877));
   BUFCHD FE_PHC5451_n3116 (.O(FE_PHN5451_n3116), 
	.I(FE_PHN6108_n3116));
   BUFCKEHD FE_PHC5450_n3918 (.O(FE_PHN5450_n3918), 
	.I(FE_PHN6300_n3918));
   BUFCHD FE_PHC5449_n902 (.O(FE_PHN5449_n902), 
	.I(FE_PHN6858_n902));
   BUFCKEHD FE_PHC5448_n3094 (.O(FE_PHN5448_n3094), 
	.I(FE_PHN6238_n3094));
   BUFCHD FE_PHC5447_ram_145__7_ (.O(FE_PHN5447_ram_145__7_), 
	.I(FE_PHN6064_ram_145__7_));
   BUFCHD FE_PHC5446_n850 (.O(FE_PHN5446_n850), 
	.I(FE_PHN6310_n850));
   BUFCHD FE_PHC5445_n4183 (.O(FE_PHN5445_n4183), 
	.I(FE_PHN6079_n4183));
   BUFCHD FE_PHC5444_n1042 (.O(FE_PHN5444_n1042), 
	.I(FE_PHN6231_n1042));
   BUFCHD FE_PHC5443_n4240 (.O(FE_PHN5443_n4240), 
	.I(FE_PHN5929_n4240));
   BUFCHD FE_PHC5442_n2943 (.O(FE_PHN5442_n2943), 
	.I(FE_PHN6040_n2943));
   BUFCHD FE_PHC5441_n1005 (.O(FE_PHN5441_n1005), 
	.I(FE_PHN6234_n1005));
   BUFGHD FE_PHC5440_n4215 (.O(FE_PHN5440_n4215), 
	.I(FE_PHN5911_n4215));
   BUFCHD FE_PHC5439_n3141 (.O(FE_PHN5439_n3141), 
	.I(FE_PHN6320_n3141));
   BUFCHD FE_PHC5438_n839 (.O(FE_PHN5438_n839), 
	.I(FE_PHN6107_n839));
   BUFCHD FE_PHC5437_n847 (.O(FE_PHN5437_n847), 
	.I(FE_PHN6287_n847));
   BUFCHD FE_PHC5436_n3210 (.O(FE_PHN5436_n3210), 
	.I(FE_PHN6135_n3210));
   BUFCHD FE_PHC5435_n3126 (.O(FE_PHN5435_n3126), 
	.I(FE_PHN6341_n3126));
   BUFCHD FE_PHC5434_n1000 (.O(FE_PHN5434_n1000), 
	.I(FE_PHN6299_n1000));
   BUFCHD FE_PHC5433_n986 (.O(FE_PHN5433_n986), 
	.I(FE_PHN6279_n986));
   BUFCHD FE_PHC5432_n892 (.O(FE_PHN5432_n892), 
	.I(FE_PHN6023_n892));
   BUFCHD FE_PHC5431_n966 (.O(FE_PHN5431_n966), 
	.I(FE_PHN6346_n966));
   BUFCHD FE_PHC5430_n3972 (.O(FE_PHN5430_n3972), 
	.I(FE_PHN6132_n3972));
   BUFCHD FE_PHC5429_n869 (.O(FE_PHN5429_n869), 
	.I(FE_PHN6276_n869));
   BUFCHD FE_PHC5428_n3134 (.O(FE_PHN5428_n3134), 
	.I(FE_PHN6041_n3134));
   BUFCHD FE_PHC5427_n889 (.O(FE_PHN5427_n889), 
	.I(FE_PHN6027_n889));
   BUFCHD FE_PHC5426_n3011 (.O(FE_PHN5426_n3011), 
	.I(FE_PHN6406_n3011));
   BUFCHD FE_PHC5425_n3959 (.O(FE_PHN5425_n3959), 
	.I(FE_PHN6097_n3959));
   BUFCHD FE_PHC5424_n3112 (.O(FE_PHN5424_n3112), 
	.I(FE_PHN6059_n3112));
   BUFCHD FE_PHC5423_n3108 (.O(FE_PHN5423_n3108), 
	.I(FE_PHN6225_n3108));
   BUFCHD FE_PHC5422_n856 (.O(FE_PHN5422_n856), 
	.I(FE_PHN6048_n856));
   BUFCKGHD FE_PHC5421_n3976 (.O(FE_PHN5421_n3976), 
	.I(FE_PHN5990_n3976));
   BUFCHD FE_PHC5420_n4164 (.O(FE_PHN5420_n4164), 
	.I(FE_PHN5909_n4164));
   BUFCKIHD FE_PHC5419_n1021 (.O(FE_PHN5419_n1021), 
	.I(FE_PHN6044_n1021));
   BUFCHD FE_PHC5418_n4211 (.O(FE_PHN5418_n4211), 
	.I(FE_PHN6038_n4211));
   BUFCHD FE_PHC5417_n3013 (.O(FE_PHN5417_n3013), 
	.I(FE_PHN6161_n3013));
   BUFCHD FE_PHC5416_n2986 (.O(FE_PHN5416_n2986), 
	.I(FE_PHN6258_n2986));
   BUFEHD FE_PHC5415_n3916 (.O(FE_PHN5415_n3916), 
	.I(FE_PHN5967_n3916));
   BUFCHD FE_PHC5414_n991 (.O(FE_PHN5414_n991), 
	.I(FE_PHN6375_n991));
   BUFCHD FE_PHC5413_n3943 (.O(FE_PHN5413_n3943), 
	.I(FE_PHN6077_n3943));
   BUFCHD FE_PHC5412_n3124 (.O(FE_PHN5412_n3124), 
	.I(FE_PHN6217_n3124));
   BUFCHD FE_PHC5411_n4212 (.O(FE_PHN5411_n4212), 
	.I(FE_PHN6303_n4212));
   BUFCHD FE_PHC5410_ram_31__2_ (.O(FE_PHN5410_ram_31__2_), 
	.I(FE_PHN6269_ram_31__2_));
   BUFCHD FE_PHC5409_n3024 (.O(FE_PHN5409_n3024), 
	.I(FE_PHN6112_n3024));
   BUFCHD FE_PHC5408_n1020 (.O(FE_PHN5408_n1020), 
	.I(FE_PHN6098_n1020));
   BUFCHD FE_PHC5407_n993 (.O(FE_PHN5407_n993), 
	.I(FE_PHN6246_n993));
   BUFCHD FE_PHC5406_n3070 (.O(FE_PHN5406_n3070), 
	.I(FE_PHN6141_n3070));
   BUFCHD FE_PHC5405_n2888 (.O(FE_PHN5405_n2888), 
	.I(FE_PHN6085_n2888));
   BUFCHD FE_PHC5404_n3060 (.O(FE_PHN5404_n3060), 
	.I(FE_PHN6033_n3060));
   BUFCHD FE_PHC5403_n3258 (.O(FE_PHN5403_n3258), 
	.I(FE_PHN5922_n3258));
   BUFCHD FE_PHC5402_n3137 (.O(FE_PHN5402_n3137), 
	.I(FE_PHN6369_n3137));
   BUFCHD FE_PHC5401_n3040 (.O(FE_PHN5401_n3040), 
	.I(FE_PHN5833_n3040));
   BUFCHD FE_PHC5400_n882 (.O(FE_PHN5400_n882), 
	.I(FE_PHN6198_n882));
   BUFCKEHD FE_PHC5399_n3028 (.O(FE_PHN5399_n3028), 
	.I(FE_PHN5941_n3028));
   BUFCKLHD FE_PHC5398_n4392 (.O(FE_PHN5398_n4392), 
	.I(FE_PHN3620_n4392));
   BUFCHD FE_PHC5397_n4355 (.O(FE_PHN5397_n4355), 
	.I(FE_PHN5958_n4355));
   BUFCKGHD FE_PHC5396_n969 (.O(FE_PHN5396_n969), 
	.I(FE_PHN6145_n969));
   BUFCHD FE_PHC5395_n4225 (.O(FE_PHN5395_n4225), 
	.I(FE_PHN6009_n4225));
   BUFCKKHD FE_PHC5394_n4364 (.O(FE_PHN5394_n4364), 
	.I(FE_PHN6297_n4364));
   BUFCHD FE_PHC5393_n4188 (.O(FE_PHN5393_n4188), 
	.I(FE_PHN5988_n4188));
   BUFCHD FE_PHC5392_n3993 (.O(FE_PHN5392_n3993), 
	.I(FE_PHN6111_n3993));
   BUFCHD FE_PHC5391_n4209 (.O(FE_PHN5391_n4209), 
	.I(FE_PHN5887_n4209));
   BUFCHD FE_PHC5390_n4222 (.O(FE_PHN5390_n4222), 
	.I(FE_PHN6072_n4222));
   BUFCHD FE_PHC5389_n2995 (.O(FE_PHN5389_n2995), 
	.I(FE_PHN5992_n2995));
   BUFCHD FE_PHC5388_n3989 (.O(FE_PHN5388_n3989), 
	.I(FE_PHN6180_n3989));
   BUFCKEHD FE_PHC5387_n3118 (.O(FE_PHN5387_n3118), 
	.I(FE_PHN6352_n3118));
   BUFCHD FE_PHC5386_ram_133__9_ (.O(FE_PHN5386_ram_133__9_), 
	.I(FE_PHN6021_ram_133__9_));
   BUFCHD FE_PHC5385_n976 (.O(FE_PHN5385_n976), 
	.I(FE_PHN6376_n976));
   BUFCHD FE_PHC5384_n3130 (.O(FE_PHN5384_n3130), 
	.I(FE_PHN6233_n3130));
   BUFCHD FE_PHC5383_n4029 (.O(FE_PHN5383_n4029), 
	.I(FE_PHN5940_n4029));
   BUFMHD FE_PHC5382_n4179 (.O(FE_PHN5382_n4179), 
	.I(n4179));
   BUFCHD FE_PHC5381_n911 (.O(FE_PHN5381_n911), 
	.I(FE_PHN5933_n911));
   BUFCHD FE_PHC5380_n3255 (.O(FE_PHN5380_n3255), 
	.I(FE_PHN6067_n3255));
   BUFCHD FE_PHC5379_n2916 (.O(FE_PHN5379_n2916), 
	.I(FE_PHN6083_n2916));
   BUFCHD FE_PHC5378_n3140 (.O(FE_PHN5378_n3140), 
	.I(FE_PHN6423_n3140));
   BUFCHD FE_PHC5377_n1014 (.O(FE_PHN5377_n1014), 
	.I(FE_PHN6035_n1014));
   BUFCHD FE_PHC5376_n3022 (.O(FE_PHN5376_n3022), 
	.I(FE_PHN6068_n3022));
   BUFCHD FE_PHC5375_n4396 (.O(FE_PHN5375_n4396), 
	.I(FE_PHN6284_n4396));
   BUFCKEHD FE_PHC5374_n3090 (.O(FE_PHN5374_n3090), 
	.I(FE_PHN6397_n3090));
   BUFCHD FE_PHC5373_n4251 (.O(FE_PHN5373_n4251), 
	.I(FE_PHN6074_n4251));
   BUFCHD FE_PHC5372_n4373 (.O(FE_PHN5372_n4373), 
	.I(FE_PHN6283_n4373));
   BUFCHD FE_PHC5371_n1024 (.O(FE_PHN5371_n1024), 
	.I(FE_PHN6307_n1024));
   BUFCHD FE_PHC5370_n3015 (.O(FE_PHN5370_n3015), 
	.I(FE_PHN6301_n3015));
   BUFGHD FE_PHC5369_n4226 (.O(FE_PHN5369_n4226), 
	.I(FE_PHN5893_n4226));
   BUFCHD FE_PHC5368_n3964 (.O(FE_PHN5368_n3964), 
	.I(FE_PHN5915_n3964));
   BUFHHD FE_PHC5367_n4178 (.O(FE_PHN5367_n4178), 
	.I(FE_PHN3665_n4178));
   BUFCHD FE_PHC5366_n4167 (.O(FE_PHN5366_n4167), 
	.I(FE_PHN6230_n4167));
   BUFCHD FE_PHC5365_n1016 (.O(FE_PHN5365_n1016), 
	.I(FE_PHN6343_n1016));
   BUFCHD FE_PHC5364_n4172 (.O(FE_PHN5364_n4172), 
	.I(FE_PHN5969_n4172));
   BUFCHD FE_PHC5363_n2984 (.O(FE_PHN5363_n2984), 
	.I(FE_PHN6131_n2984));
   BUFCHD FE_PHC5362_n4394 (.O(FE_PHN5362_n4394), 
	.I(FE_PHN6125_n4394));
   BUFCHD FE_PHC5361_n2420 (.O(FE_PHN5361_n2420), 
	.I(FE_PHN5894_n2420));
   BUFCHD FE_PHC5360_n4199 (.O(FE_PHN5360_n4199), 
	.I(FE_PHN6222_n4199));
   BUFCHD FE_PHC5359_n4023 (.O(FE_PHN5359_n4023), 
	.I(FE_PHN6294_n4023));
   BUFCKMHD FE_PHC5358_n903 (.O(FE_PHN5358_n903), 
	.I(FE_PHN6210_n903));
   BUFCHD FE_PHC5357_n2564 (.O(FE_PHN5357_n2564), 
	.I(FE_PHN5881_n2564));
   BUFCHD FE_PHC5356_n2959 (.O(FE_PHN5356_n2959), 
	.I(FE_PHN6197_n2959));
   BUFCHD FE_PHC5355_n866 (.O(FE_PHN5355_n866), 
	.I(FE_PHN5996_n866));
   BUFCHD FE_PHC5354_n3910 (.O(FE_PHN5354_n3910), 
	.I(FE_PHN6043_n3910));
   BUFCKJHD FE_PHC5353_n4030 (.O(FE_PHN5353_n4030), 
	.I(FE_PHN5974_n4030));
   BUFCHD FE_PHC5352_n3942 (.O(FE_PHN5352_n3942), 
	.I(FE_PHN6157_n3942));
   BUFCHD FE_PHC5351_n3014 (.O(FE_PHN5351_n3014), 
	.I(FE_PHN6236_n3014));
   BUFCHD FE_PHC5350_n861 (.O(FE_PHN5350_n861), 
	.I(FE_PHN5953_n861));
   BUFCHD FE_PHC5349_n4311 (.O(FE_PHN5349_n4311), 
	.I(FE_PHN6026_n4311));
   BUFEHD FE_PHC5348_n2580 (.O(FE_PHN5348_n2580), 
	.I(FE_PHN5834_n2580));
   BUFCKJHD FE_PHC5347_n2970 (.O(FE_PHN5347_n2970), 
	.I(FE_PHN5985_n2970));
   BUFCHD FE_PHC5346_n858 (.O(FE_PHN5346_n858), 
	.I(FE_PHN5883_n858));
   BUFCHD FE_PHC5345_n4368 (.O(FE_PHN5345_n4368), 
	.I(FE_PHN6315_n4368));
   BUFCHD FE_PHC5344_n4340 (.O(FE_PHN5344_n4340), 
	.I(FE_PHN5956_n4340));
   BUFCHD FE_PHC5343_n2997 (.O(FE_PHN5343_n2997), 
	.I(FE_PHN6122_n2997));
   BUFCHD FE_PHC5342_n849 (.O(FE_PHN5342_n849), 
	.I(FE_PHN6256_n849));
   BUFCHD FE_PHC5341_n997 (.O(FE_PHN5341_n997), 
	.I(FE_PHN6281_n997));
   BUFCHD FE_PHC5340_n2993 (.O(FE_PHN5340_n2993), 
	.I(FE_PHN6174_n2993));
   BUFCHD FE_PHC5339_n4402 (.O(FE_PHN5339_n4402), 
	.I(FE_PHN6105_n4402));
   BUFCHD FE_PHC5338_n3136 (.O(FE_PHN5338_n3136), 
	.I(FE_PHN6182_n3136));
   BUFCHD FE_PHC5337_n4046 (.O(FE_PHN5337_n4046), 
	.I(FE_PHN5856_n4046));
   BUFCHD FE_PHC5336_n4283 (.O(FE_PHN5336_n4283), 
	.I(FE_PHN6302_n4283));
   BUFCHD FE_PHC5335_n2754 (.O(FE_PHN5335_n2754), 
	.I(FE_PHN5897_n2754));
   BUFCHD FE_PHC5334_n4418 (.O(FE_PHN5334_n4418), 
	.I(FE_PHN6025_n4418));
   BUFCHD FE_PHC5333_n2992 (.O(FE_PHN5333_n2992), 
	.I(FE_PHN5993_n2992));
   BUFCHD FE_PHC5332_n4284 (.O(FE_PHN5332_n4284), 
	.I(FE_PHN6106_n4284));
   BUFCHD FE_PHC5331_n2946 (.O(FE_PHN5331_n2946), 
	.I(FE_PHN6116_n2946));
   BUFCHD FE_PHC5330_n959 (.O(FE_PHN5330_n959), 
	.I(FE_PHN5859_n959));
   BUFCHD FE_PHC5329_n3086 (.O(FE_PHN5329_n3086), 
	.I(FE_PHN6152_n3086));
   BUFCHD FE_PHC5328_n3098 (.O(FE_PHN5328_n3098), 
	.I(FE_PHN6051_n3098));
   BUFCHD FE_PHC5327_n3958 (.O(FE_PHN5327_n3958), 
	.I(FE_PHN5998_n3958));
   BUFCKLHD FE_PHC5326_n897 (.O(FE_PHN5326_n897), 
	.I(FE_PHN6237_n897));
   BUFCHD FE_PHC5325_n941 (.O(FE_PHN5325_n941), 
	.I(FE_PHN6052_n941));
   BUFCHD FE_PHC5324_n4252 (.O(FE_PHN5324_n4252), 
	.I(FE_PHN5898_n4252));
   BUFCHD FE_PHC5323_n3067 (.O(FE_PHN5323_n3067), 
	.I(FE_PHN6054_n3067));
   BUFCHD FE_PHC5322_n3131 (.O(FE_PHN5322_n3131), 
	.I(FE_PHN6036_n3131));
   BUFCHD FE_PHC5321_n2998 (.O(FE_PHN5321_n2998), 
	.I(FE_PHN5963_n2998));
   BUFCHD FE_PHC5320_n2950 (.O(FE_PHN5320_n2950), 
	.I(FE_PHN6058_n2950));
   BUFCHD FE_PHC5319_n3089 (.O(FE_PHN5319_n3089), 
	.I(FE_PHN6339_n3089));
   BUFCHD FE_PHC5318_n4281 (.O(FE_PHN5318_n4281), 
	.I(FE_PHN6148_n4281));
   BUFCKLHD FE_PHC5317_n3064 (.O(FE_PHN5317_n3064), 
	.I(FE_PHN6361_n3064));
   BUFCHD FE_PHC5316_n4408 (.O(FE_PHN5316_n4408), 
	.I(FE_PHN6169_n4408));
   BUFCHD FE_PHC5315_n885 (.O(FE_PHN5315_n885), 
	.I(FE_PHN6137_n885));
   BUFCHD FE_PHC5314_n3025 (.O(FE_PHN5314_n3025), 
	.I(FE_PHN6017_n3025));
   BUFCKLHD FE_PHC5313_n4185 (.O(FE_PHN5313_n4185), 
	.I(FE_PHN6289_n4185));
   BUFCHD FE_PHC5312_n3042 (.O(FE_PHN5312_n3042), 
	.I(FE_PHN6264_n3042));
   BUFNHD FE_PHC5311_n2753 (.O(FE_PHN5311_n2753), 
	.I(n2753));
   BUFCHD FE_PHC5310_n4416 (.O(FE_PHN5310_n4416), 
	.I(FE_PHN6176_n4416));
   BUFCKLHD FE_PHC5309_n4166 (.O(FE_PHN5309_n4166), 
	.I(FE_PHN6292_n4166));
   BUFCHD FE_PHC5308_n4204 (.O(FE_PHN5308_n4204), 
	.I(FE_PHN6063_n4204));
   BUFCHD FE_PHC5307_n1013 (.O(FE_PHN5307_n1013), 
	.I(FE_PHN5947_n1013));
   BUFCHD FE_PHC5306_n1006 (.O(FE_PHN5306_n1006), 
	.I(FE_PHN6029_n1006));
   BUFCHD FE_PHC5305_n3125 (.O(FE_PHN5305_n3125), 
	.I(FE_PHN6232_n3125));
   BUFCHD FE_PHC5304_n4415 (.O(FE_PHN5304_n4415), 
	.I(FE_PHN6142_n4415));
   BUFCHD FE_PHC5303_n840 (.O(FE_PHN5303_n840), 
	.I(FE_PHN6019_n840));
   BUFCHD FE_PHC5302_n3963 (.O(FE_PHN5302_n3963), 
	.I(FE_PHN5948_n3963));
   BUFCHD FE_PHC5301_n3087 (.O(FE_PHN5301_n3087), 
	.I(FE_PHN6128_n3087));
   BUFCHD FE_PHC5300_n3105 (.O(FE_PHN5300_n3105), 
	.I(FE_PHN6337_n3105));
   BUFCHD FE_PHC5299_n4299 (.O(FE_PHN5299_n4299), 
	.I(FE_PHN5907_n4299));
   BUFCKKHD FE_PHC5298_n4203 (.O(FE_PHN5298_n4203), 
	.I(FE_PHN6042_n4203));
   BUFCHD FE_PHC5297_n2178 (.O(FE_PHN5297_n2178), 
	.I(FE_PHN5850_n2178));
   BUFCKMHD FE_PHC5296_n2297 (.O(FE_PHN5296_n2297), 
	.I(FE_PHN4009_n2297));
   BUFCHD FE_PHC5295_n3924 (.O(FE_PHN5295_n3924), 
	.I(FE_PHN6066_n3924));
   BUFCHD FE_PHC5294_n3985 (.O(FE_PHN5294_n3985), 
	.I(FE_PHN6186_n3985));
   BUFCHD FE_PHC5293_n876 (.O(FE_PHN5293_n876), 
	.I(FE_PHN5972_n876));
   BUFCHD FE_PHC5292_n4360 (.O(FE_PHN5292_n4360), 
	.I(FE_PHN6003_n4360));
   BUFCHD FE_PHC5291_n4007 (.O(FE_PHN5291_n4007), 
	.I(FE_PHN6093_n4007));
   BUFGHD FE_PHC5290_n2405 (.O(FE_PHN5290_n2405), 
	.I(FE_PHN5839_n2405));
   BUFCHD FE_PHC5289_n3023 (.O(FE_PHN5289_n3023), 
	.I(FE_PHN5989_n3023));
   BUFCHD FE_PHC5288_n4350 (.O(FE_PHN5288_n4350), 
	.I(FE_PHN5852_n4350));
   BUFCHD FE_PHC5287_n913 (.O(FE_PHN5287_n913), 
	.I(FE_PHN5983_n913));
   BUFCHD FE_PHC5286_n3103 (.O(FE_PHN5286_n3103), 
	.I(FE_PHN6092_n3103));
   BUFCHD FE_PHC5285_n4196 (.O(FE_PHN5285_n4196), 
	.I(FE_PHN6163_n4196));
   BUFCHD FE_PHC5284_n3257 (.O(FE_PHN5284_n3257), 
	.I(FE_PHN5923_n3257));
   BUFCHD FE_PHC5283_n975 (.O(FE_PHN5283_n975), 
	.I(FE_PHN5926_n975));
   BUFCHD FE_PHC5282_n2936 (.O(FE_PHN5282_n2936), 
	.I(FE_PHN5903_n2936));
   BUFCHD FE_PHC5281_n943 (.O(FE_PHN5281_n943), 
	.I(FE_PHN6794_n943));
   BUFCHD FE_PHC5280_n957 (.O(FE_PHN5280_n957), 
	.I(FE_PHN5970_n957));
   BUFCHD FE_PHC5279_n3138 (.O(FE_PHN5279_n3138), 
	.I(FE_PHN6305_n3138));
   BUFCHD FE_PHC5278_n2954 (.O(FE_PHN5278_n2954), 
	.I(FE_PHN6088_n2954));
   BUFCHD FE_PHC5277_n1079 (.O(FE_PHN5277_n1079), 
	.I(FE_PHN5954_n1079));
   BUFCHD FE_PHC5276_n1106 (.O(FE_PHN5276_n1106), 
	.I(FE_PHN5867_n1106));
   BUFCHD FE_PHC5275_n2980 (.O(FE_PHN5275_n2980), 
	.I(FE_PHN6120_n2980));
   BUFCHD FE_PHC5274_n4025 (.O(FE_PHN5274_n4025), 
	.I(FE_PHN6318_n4025));
   BUFCHD FE_PHC5273_ram_153__11_ (.O(FE_PHN5273_ram_153__11_), 
	.I(FE_PHN5986_ram_153__11_));
   BUFCHD FE_PHC5272_n1018 (.O(FE_PHN5272_n1018), 
	.I(FE_PHN6214_n1018));
   BUFCHD FE_PHC5271_n881 (.O(FE_PHN5271_n881), 
	.I(FE_PHN6006_n881));
   BUFCHD FE_PHC5270_n2996 (.O(FE_PHN5270_n2996), 
	.I(FE_PHN6095_n2996));
   BUFCHD FE_PHC5269_n3996 (.O(FE_PHN5269_n3996), 
	.I(FE_PHN6055_n3996));
   BUFCHD FE_PHC5268_n905 (.O(FE_PHN5268_n905), 
	.I(FE_PHN5882_n905));
   BUFCHD FE_PHC5267_n4419 (.O(FE_PHN5267_n4419), 
	.I(FE_PHN6013_n4419));
   BUFCKLHD FE_PHC5266_n3065 (.O(FE_PHN5266_n3065), 
	.I(FE_PHN6349_n3065));
   BUFCHD FE_PHC5265_n4217 (.O(FE_PHN5265_n4217), 
	.I(FE_PHN5961_n4217));
   BUFCHD FE_PHC5264_n3006 (.O(FE_PHN5264_n3006), 
	.I(FE_PHN6164_n3006));
   BUFCHD FE_PHC5263_n4049 (.O(FE_PHN5263_n4049), 
	.I(FE_PHN5825_n4049));
   BUFCHD FE_PHC5262_n1920 (.O(FE_PHN5262_n1920), 
	.I(FE_PHN5873_n1920));
   BUFCHD FE_PHC5261_n3207 (.O(FE_PHN5261_n3207), 
	.I(FE_PHN5901_n3207));
   BUFCHD FE_PHC5260_n4220 (.O(FE_PHN5260_n4220), 
	.I(FE_PHN5928_n4220));
   BUFCKKHD FE_PHC5259_n4383 (.O(FE_PHN5259_n4383), 
	.I(FE_PHN6309_n4383));
   BUFCKJHD FE_PHC5258_n4277 (.O(FE_PHN5258_n4277), 
	.I(FE_PHN5858_n4277));
   BUFCHD FE_PHC5257_n4278 (.O(FE_PHN5257_n4278), 
	.I(FE_PHN5824_n4278));
   BUFCHD FE_PHC5256_n2927 (.O(FE_PHN5256_n2927), 
	.I(FE_PHN5880_n2927));
   BUFCHD FE_PHC5255_n972 (.O(FE_PHN5255_n972), 
	.I(FE_PHN5842_n972));
   BUFCKEHD FE_PHC5254_n2384 (.O(FE_PHN5254_n2384), 
	.I(FE_PHN5874_n2384));
   BUFCHD FE_PHC5253_n2897 (.O(FE_PHN5253_n2897), 
	.I(FE_PHN5968_n2897));
   BUFCHD FE_PHC5252_n1037 (.O(FE_PHN5252_n1037), 
	.I(FE_PHN5925_n1037));
   BUFCHD FE_PHC5251_n935 (.O(FE_PHN5251_n935), 
	.I(FE_PHN5884_n935));
   BUFLHD FE_PHC5250_n3069 (.O(FE_PHN5250_n3069), 
	.I(FE_PHN3743_n3069));
   BUFCHD FE_PHC5249_n994 (.O(FE_PHN5249_n994), 
	.I(FE_PHN5991_n994));
   BUFCHD FE_PHC5248_n965 (.O(FE_PHN5248_n965), 
	.I(FE_PHN5919_n965));
   BUFCHD FE_PHC5247_n894 (.O(FE_PHN5247_n894), 
	.I(FE_PHN5865_n894));
   BUFCHD FE_PHC5246_n2574 (.O(FE_PHN5246_n2574), 
	.I(FE_PHN5843_n2574));
   BUFCHD FE_PHC5245_n2987 (.O(FE_PHN5245_n2987), 
	.I(FE_PHN5942_n2987));
   BUFCHD FE_PHC5244_n3082 (.O(FE_PHN5244_n3082), 
	.I(FE_PHN5951_n3082));
   BUFCHD FE_PHC5243_n3969 (.O(FE_PHN5243_n3969), 
	.I(FE_PHN6073_n3969));
   BUFCHD FE_PHC5242_n3002 (.O(FE_PHN5242_n3002), 
	.I(FE_PHN5943_n3002));
   BUFCHD FE_PHC5241_n1870 (.O(FE_PHN5241_n1870), 
	.I(FE_PHN5822_n1870));
   BUFCHD FE_PHC5240_n2722 (.O(FE_PHN5240_n2722), 
	.I(FE_PHN5924_n2722));
   BUFCHD FE_PHC5239_n1002 (.O(FE_PHN5239_n1002), 
	.I(FE_PHN6306_n1002));
   BUFCHD FE_PHC5238_n4232 (.O(FE_PHN5238_n4232), 
	.I(FE_PHN5820_n4232));
   BUFCHD FE_PHC5237_n3029 (.O(FE_PHN5237_n3029), 
	.I(FE_PHN5946_n3029));
   BUFCKMHD FE_PHC5236_n841 (.O(FE_PHN5236_n841), 
	.I(FE_PHN6401_n841));
   BUFCHD FE_PHC5235_n4378 (.O(FE_PHN5235_n4378), 
	.I(FE_PHN5935_n4378));
   BUFCKGHD FE_PHC5234_n2385 (.O(FE_PHN5234_n2385), 
	.I(FE_PHN3939_n2385));
   BUFCHD FE_PHC5233_n3075 (.O(FE_PHN5233_n3075), 
	.I(FE_PHN5960_n3075));
   BUFCKMHD FE_PHC5232_n4316 (.O(FE_PHN5232_n4316), 
	.I(FE_PHN6373_n4316));
   BUFCHD FE_PHC5231_n3026 (.O(FE_PHN5231_n3026), 
	.I(FE_PHN6291_n3026));
   BUFCHD FE_PHC5230_n4174 (.O(FE_PHN5230_n4174), 
	.I(FE_PHN5832_n4174));
   BUFCHD FE_PHC5229_n2930 (.O(FE_PHN5229_n2930), 
	.I(FE_PHN6005_n2930));
   BUFCKMHD FE_PHC5228_n4206 (.O(FE_PHN5228_n4206), 
	.I(FE_PHN3399_n4206));
   BUFCKMHD FE_PHC5227_n4342 (.O(FE_PHN5227_n4342), 
	.I(FE_PHN4415_n4342));
   BUFCHD FE_PHC5226_n3998 (.O(FE_PHN5226_n3998), 
	.I(FE_PHN6069_n3998));
   BUFCHD FE_PHC5225_n2964 (.O(FE_PHN5225_n2964), 
	.I(FE_PHN5904_n2964));
   BUFCHD FE_PHC5224_n4400 (.O(FE_PHN5224_n4400), 
	.I(FE_PHN5932_n4400));
   BUFCHD FE_PHC5223_n929 (.O(FE_PHN5223_n929), 
	.I(FE_PHN5957_n929));
   BUFCHD FE_PHC5222_n4255 (.O(FE_PHN5222_n4255), 
	.I(FE_PHN5808_n4255));
   BUFCHD FE_PHC5221_ram_153__7_ (.O(FE_PHN5221_ram_153__7_), 
	.I(FE_PHN6102_ram_153__7_));
   BUFCHD FE_PHC5220_n3054 (.O(FE_PHN5220_n3054), 
	.I(FE_PHN6239_n3054));
   BUFCHD FE_PHC5219_n4380 (.O(FE_PHN5219_n4380), 
	.I(FE_PHN6123_n4380));
   BUFCHD FE_PHC5218_n3074 (.O(FE_PHN5218_n3074), 
	.I(FE_PHN6189_n3074));
   BUFCHD FE_PHC5217_n3219 (.O(FE_PHN5217_n3219), 
	.I(FE_PHN5807_n3219));
   BUFCHD FE_PHC5216_n4037 (.O(FE_PHN5216_n4037), 
	.I(FE_PHN6071_n4037));
   BUFCKLHD FE_PHC5215_n4286 (.O(FE_PHN5215_n4286), 
	.I(FE_PHN6333_n4286));
   BUFCHD FE_PHC5214_n3987 (.O(FE_PHN5214_n3987), 
	.I(FE_PHN5984_n3987));
   BUFCHD FE_PHC5213_n864 (.O(FE_PHN5213_n864), 
	.I(FE_PHN5920_n864));
   BUFCHD FE_PHC5212_n3048 (.O(FE_PHN5212_n3048), 
	.I(FE_PHN5939_n3048));
   BUFCHD FE_PHC5211_n4377 (.O(FE_PHN5211_n4377), 
	.I(FE_PHN5896_n4377));
   BUFCHD FE_PHC5210_n3020 (.O(FE_PHN5210_n3020), 
	.I(FE_PHN5952_n3020));
   BUFCHD FE_PHC5209_n948 (.O(FE_PHN5209_n948), 
	.I(FE_PHN5806_n948));
   BUFCKEHD FE_PHC5208_n988 (.O(FE_PHN5208_n988), 
	.I(FE_PHN3922_n988));
   BUFCKMHD FE_PHC5207_n2891 (.O(FE_PHN5207_n2891), 
	.I(FE_PHN6422_n2891));
   BUFCHD FE_PHC5206_n3093 (.O(FE_PHN5206_n3093), 
	.I(FE_PHN6001_n3093));
   BUFCHD FE_PHC5205_n4393 (.O(FE_PHN5205_n4393), 
	.I(FE_PHN5860_n4393));
   BUFCHD FE_PHC5204_n890 (.O(FE_PHN5204_n890), 
	.I(FE_PHN6031_n890));
   BUFCHD FE_PHC5203_ram_145__0_ (.O(FE_PHN5203_ram_145__0_), 
	.I(FE_PHN6024_ram_145__0_));
   BUFCHD FE_PHC5202_n982 (.O(FE_PHN5202_n982), 
	.I(FE_PHN6178_n982));
   BUFCHD FE_PHC5201_n3992 (.O(FE_PHN5201_n3992), 
	.I(FE_PHN5877_n3992));
   BUFCHD FE_PHC5200_n2975 (.O(FE_PHN5200_n2975), 
	.I(FE_PHN6086_n2975));
   BUFCHD FE_PHC5199_n4021 (.O(FE_PHN5199_n4021), 
	.I(FE_PHN5945_n4021));
   BUFCHD FE_PHC5198_n3055 (.O(FE_PHN5198_n3055), 
	.I(FE_PHN5930_n3055));
   BUFCHD FE_PHC5197_n2991 (.O(FE_PHN5197_n2991), 
	.I(FE_PHN6151_n2991));
   BUFCHD FE_PHC5196_n910 (.O(FE_PHN5196_n910), 
	.I(FE_PHN5906_n910));
   BUFCHD FE_PHC5195_n2735 (.O(FE_PHN5195_n2735), 
	.I(FE_PHN5936_n2735));
   BUFCHD FE_PHC5194_n2989 (.O(FE_PHN5194_n2989), 
	.I(FE_PHN6012_n2989));
   BUFCHD FE_PHC5193_n3104 (.O(FE_PHN5193_n3104), 
	.I(FE_PHN6220_n3104));
   BUFCHD FE_PHC5192_n887 (.O(FE_PHN5192_n887), 
	.I(FE_PHN6834_n887));
   BUFCHD FE_PHC5191_n1029 (.O(FE_PHN5191_n1029), 
	.I(FE_PHN6293_n1029));
   BUFCHD FE_PHC5190_n3012 (.O(FE_PHN5190_n3012), 
	.I(FE_PHN6266_n3012));
   BUFCHD FE_PHC5189_n3122 (.O(FE_PHN5189_n3122), 
	.I(FE_PHN6183_n3122));
   BUFCHD FE_PHC5188_n878 (.O(FE_PHN5188_n878), 
	.I(FE_PHN5827_n878));
   BUFCHD FE_PHC5187_n1017 (.O(FE_PHN5187_n1017), 
	.I(FE_PHN5851_n1017));
   BUFCHD FE_PHC5186_n936 (.O(FE_PHN5186_n936), 
	.I(FE_PHN5800_n936));
   BUFCHD FE_PHC5185_n3050 (.O(FE_PHN5185_n3050), 
	.I(FE_PHN6121_n3050));
   BUFCHD FE_PHC5184_n3007 (.O(FE_PHN5184_n3007), 
	.I(FE_PHN6075_n3007));
   BUFCKLHD FE_PHC5183_n3063 (.O(FE_PHN5183_n3063), 
	.I(FE_PHN6227_n3063));
   BUFCHD FE_PHC5182_n3919 (.O(FE_PHN5182_n3919), 
	.I(FE_PHN5812_n3919));
   BUFCHD FE_PHC5181_n3921 (.O(FE_PHN5181_n3921), 
	.I(FE_PHN6119_n3921));
   BUFCKLHD FE_PHC5180_n4411 (.O(FE_PHN5180_n4411), 
	.I(FE_PHN3316_n4411));
   BUFCHD FE_PHC5179_n3052 (.O(FE_PHN5179_n3052), 
	.I(FE_PHN5879_n3052));
   BUFCKLHD FE_PHC5178_n4363 (.O(FE_PHN5178_n4363), 
	.I(FE_PHN6419_n4363));
   BUFCHD FE_PHC5177_n4369 (.O(FE_PHN5177_n4369), 
	.I(FE_PHN5937_n4369));
   BUFCKMHD FE_PHC5176_n4285 (.O(FE_PHN5176_n4285), 
	.I(FE_PHN6429_n4285));
   BUFCKMHD FE_PHC5175_n2960 (.O(FE_PHN5175_n2960), 
	.I(FE_PHN6403_n2960));
   BUFCHD FE_PHC5174_n4014 (.O(FE_PHN5174_n4014), 
	.I(FE_PHN5885_n4014));
   BUFJHD FE_PHC5173_n846 (.O(FE_PHN5173_n846), 
	.I(FE_PHN3977_n846));
   BUFLHD FE_PHC5172_n1110 (.O(FE_PHN5172_n1110), 
	.I(FE_PHN3938_n1110));
   BUFCHD FE_PHC5171_n3072 (.O(FE_PHN5171_n3072), 
	.I(FE_PHN5841_n3072));
   BUFCHD FE_PHC5170_n999 (.O(FE_PHN5170_n999), 
	.I(FE_PHN6050_n999));
   BUFCHD FE_PHC5169_n4361 (.O(FE_PHN5169_n4361), 
	.I(FE_PHN5913_n4361));
   BUFNHD FE_PHC5168_n4333 (.O(FE_PHN5168_n4333), 
	.I(FE_PHN6190_n4333));
   BUFCHD FE_PHC5167_n4334 (.O(FE_PHN5167_n4334), 
	.I(FE_PHN5831_n4334));
   BUFCHD FE_PHC5166_n848 (.O(FE_PHN5166_n848), 
	.I(FE_PHN5999_n848));
   BUFCHD FE_PHC5165_n893 (.O(FE_PHN5165_n893), 
	.I(FE_PHN6000_n893));
   BUFCHD FE_PHC5164_n4229 (.O(FE_PHN5164_n4229), 
	.I(FE_PHN5787_n4229));
   BUFCHD FE_PHC5163_n3975 (.O(FE_PHN5163_n3975), 
	.I(FE_PHN6089_n3975));
   BUFCHD FE_PHC5162_n3053 (.O(FE_PHN5162_n3053), 
	.I(FE_PHN6028_n3053));
   BUFCHD FE_PHC5161_n3027 (.O(FE_PHN5161_n3027), 
	.I(FE_PHN5978_n3027));
   BUFCKKHD FE_PHC5160_n2983 (.O(FE_PHN5160_n2983), 
	.I(FE_PHN6096_n2983));
   BUFCHD FE_PHC5159_n4180 (.O(FE_PHN5159_n4180), 
	.I(FE_PHN6727_n4180));
   BUFCHD FE_PHC5158_n3974 (.O(FE_PHN5158_n3974), 
	.I(FE_PHN6181_n3974));
   BUFCHD FE_PHC5157_n4028 (.O(FE_PHN5157_n4028), 
	.I(FE_PHN5917_n4028));
   BUFCHD FE_PHC5156_n3977 (.O(FE_PHN5156_n3977), 
	.I(FE_PHN6094_n3977));
   BUFCHD FE_PHC5155_n3984 (.O(FE_PHN5155_n3984), 
	.I(FE_PHN5979_n3984));
   BUFCKMHD FE_PHC5154_n4241 (.O(FE_PHN5154_n4241), 
	.I(FE_PHN6383_n4241));
   BUFCKMHD FE_PHC5153_n2933 (.O(FE_PHN5153_n2933), 
	.I(FE_PHN6184_n2933));
   BUFCHD FE_PHC5152_n2932 (.O(FE_PHN5152_n2932), 
	.I(FE_PHN5849_n2932));
   BUFCKLHD FE_PHC5151_n865 (.O(FE_PHN5151_n865), 
	.I(FE_PHN6162_n865));
   BUFCHD FE_PHC5150_n3018 (.O(FE_PHN5150_n3018), 
	.I(FE_PHN5976_n3018));
   BUFCHD FE_PHC5149_n1077 (.O(FE_PHN5149_n1077), 
	.I(FE_PHN6078_n1077));
   BUFCHD FE_PHC5148_n925 (.O(FE_PHN5148_n925), 
	.I(FE_PHN5891_n925));
   BUFCHD FE_PHC5147_n870 (.O(FE_PHN5147_n870), 
	.I(FE_PHN5997_n870));
   BUFCHD FE_PHC5146_n4260 (.O(FE_PHN5146_n4260), 
	.I(FE_PHN6053_n4260));
   BUFCHD FE_PHC5145_n3076 (.O(FE_PHN5145_n3076), 
	.I(FE_PHN6020_n3076));
   BUFCKMHD FE_PHC5144_n4300 (.O(FE_PHN5144_n4300), 
	.I(FE_PHN6118_n4300));
   BUFCHD FE_PHC5143_n1038 (.O(FE_PHN5143_n1038), 
	.I(FE_PHN5803_n1038));
   BUFCHD FE_PHC5142_n4194 (.O(FE_PHN5142_n4194), 
	.I(FE_PHN5857_n4194));
   BUFCHD FE_PHC5141_n3263 (.O(FE_PHN5141_n3263), 
	.I(FE_PHN5802_n3263));
   BUFCKLHD FE_PHC5140_n3079 (.O(FE_PHN5140_n3079), 
	.I(FE_PHN6196_n3079));
   BUFCKLHD FE_PHC5139_n4327 (.O(FE_PHN5139_n4327), 
	.I(FE_PHN6208_n4327));
   BUFCKIHD FE_PHC5138_n1030 (.O(FE_PHN5138_n1030), 
	.I(FE_PHN5916_n1030));
   BUFCHD FE_PHC5137_n1072 (.O(FE_PHN5137_n1072), 
	.I(FE_PHN6061_n1072));
   BUFCKMHD FE_PHC5136_n2982 (.O(FE_PHN5136_n2982), 
	.I(FE_PHN6253_n2982));
   BUFCHD FE_PHC5135_n842 (.O(FE_PHN5135_n842), 
	.I(FE_PHN5862_n842));
   BUFCHD FE_PHC5134_n978 (.O(FE_PHN5134_n978), 
	.I(FE_PHN6271_n978));
   BUFCHD FE_PHC5133_n2951 (.O(FE_PHN5133_n2951), 
	.I(FE_PHN5845_n2951));
   BUFCHD FE_PHC5132_n3982 (.O(FE_PHN5132_n3982), 
	.I(FE_PHN6047_n3982));
   BUFCHD FE_PHC5131_n852 (.O(FE_PHN5131_n852), 
	.I(FE_PHN5864_n852));
   BUFCHD FE_PHC5130_n4243 (.O(FE_PHN5130_n4243), 
	.I(FE_PHN5938_n4243));
   BUFCHD FE_PHC5129_n3915 (.O(FE_PHN5129_n3915), 
	.I(FE_PHN5910_n3915));
   BUFCHD FE_PHC5128_n4214 (.O(FE_PHN5128_n4214), 
	.I(FE_PHN5823_n4214));
   BUFCHD FE_PHC5127_n4401 (.O(FE_PHN5127_n4401), 
	.I(FE_PHN5971_n4401));
   BUFCHD FE_PHC5126_n3948 (.O(FE_PHN5126_n3948), 
	.I(FE_PHN5890_n3948));
   BUFCHD FE_PHC5125_n1082 (.O(FE_PHN5125_n1082), 
	.I(FE_PHN5811_n1082));
   BUFCKIHD FE_PHC5124_n989 (.O(FE_PHN5124_n989), 
	.I(FE_PHN6030_n989));
   BUFCHD FE_PHC5123_n4279 (.O(FE_PHN5123_n4279), 
	.I(FE_PHN6049_n4279));
   BUFCHD FE_PHC5122_n879 (.O(FE_PHN5122_n879), 
	.I(FE_PHN6022_n879));
   BUFCKMHD FE_PHC5121_n4218 (.O(FE_PHN5121_n4218), 
	.I(FE_PHN3753_n4218));
   BUFCKJHD FE_PHC5120_n2971 (.O(FE_PHN5120_n2971), 
	.I(FE_PHN5840_n2971));
   BUFCKMHD FE_PHC5119_n4266 (.O(FE_PHN5119_n4266), 
	.I(FE_PHN6382_n4266));
   DELAKHD FE_PHC5118_n4338 (.O(FE_PHN5118_n4338), 
	.I(FE_PHN4403_n4338));
   BUFCHD FE_PHC5117_n3961 (.O(FE_PHN5117_n3961), 
	.I(FE_PHN6153_n3961));
   BUFCHD FE_PHC5116_n3929 (.O(FE_PHN5116_n3929), 
	.I(FE_PHN6010_n3929));
   BUFCHD FE_PHC5115_n3009 (.O(FE_PHN5115_n3009), 
	.I(FE_PHN6124_n3009));
   BUFCHD FE_PHC5114_n1069 (.O(FE_PHN5114_n1069), 
	.I(FE_PHN5836_n1069));
   BUFCKMHD FE_PHC5113_n1911 (.O(FE_PHN5113_n1911), 
	.I(FE_PHN6360_n1911));
   BUFCKLHD FE_PHC5112_n2988 (.O(FE_PHN5112_n2988), 
	.I(FE_PHN3315_n2988));
   BUFCKMHD FE_PHC5111_n1864 (.O(FE_PHN5111_n1864), 
	.I(FE_PHN6335_n1864));
   BUFCKMHD FE_PHC5110_n2621 (.O(FE_PHN5110_n2621), 
	.I(FE_PHN6101_n2621));
   BUFCHD FE_PHC5109_n2400 (.O(FE_PHN5109_n2400), 
	.I(FE_PHN5804_n2400));
   BUFCHD FE_PHC5108_n853 (.O(FE_PHN5108_n853), 
	.I(FE_PHN6117_n853));
   BUFCHD FE_PHC5107_n3926 (.O(FE_PHN5107_n3926), 
	.I(FE_PHN5899_n3926));
   BUFCHD FE_PHC5106_n945 (.O(FE_PHN5106_n945), 
	.I(FE_PHN5866_n945));
   BUFCKMHD FE_PHC5105_n3262 (.O(FE_PHN5105_n3262), 
	.I(FE_PHN6257_n3262));
   BUFCHD FE_PHC5104_n3092 (.O(FE_PHN5104_n3092), 
	.I(FE_PHN6228_n3092));
   BUFCHD FE_PHC5103_n3043 (.O(FE_PHN5103_n3043), 
	.I(FE_PHN5921_n3043));
   BUFCHD FE_PHC5102_n4248 (.O(FE_PHN5102_n4248), 
	.I(FE_PHN5805_n4248));
   BUFCHD FE_PHC5101_n2599 (.O(FE_PHN5101_n2599), 
	.I(FE_PHN5794_n2599));
   BUFCHD FE_PHC5100_n2945 (.O(FE_PHN5100_n2945), 
	.I(FE_PHN5838_n2945));
   BUFCHD FE_PHC5099_n1074 (.O(FE_PHN5099_n1074), 
	.I(FE_PHN6104_n1074));
   BUFCHD FE_PHC5098_n1902 (.O(FE_PHN5098_n1902), 
	.I(FE_PHN5791_n1902));
   BUFCHD FE_PHC5097_n3937 (.O(FE_PHN5097_n3937), 
	.I(FE_PHN5905_n3937));
   BUFCHD FE_PHC5096_n2976 (.O(FE_PHN5096_n2976), 
	.I(FE_PHN6018_n2976));
   BUFCHD FE_PHC5095_n946 (.O(FE_PHN5095_n946), 
	.I(FE_PHN5786_n946));
   BUFCHD FE_PHC5094_n1009 (.O(FE_PHN5094_n1009), 
	.I(FE_PHN6087_n1009));
   BUFCHD FE_PHC5093_n1064 (.O(FE_PHN5093_n1064), 
	.I(FE_PHN6175_n1064));
   BUFCHD FE_PHC5092_n992 (.O(FE_PHN5092_n992), 
	.I(FE_PHN6149_n992));
   BUFCHD FE_PHC5091_n3107 (.O(FE_PHN5091_n3107), 
	.I(FE_PHN6129_n3107));
   BUFCKKHD FE_PHC5090_n4386 (.O(FE_PHN5090_n4386), 
	.I(FE_PHN6076_n4386));
   BUFCHD FE_PHC5089_n1040 (.O(FE_PHN5089_n1040), 
	.I(FE_PHN5982_n1040));
   BUFCKMHD FE_PHC5088_n922 (.O(FE_PHN5088_n922), 
	.I(FE_PHN6344_n922));
   BUFCKGHD FE_PHC5087_n974 (.O(FE_PHN5087_n974), 
	.I(FE_PHN5792_n974));
   BUFCHD FE_PHC5086_n4405 (.O(FE_PHN5086_n4405), 
	.I(FE_PHN6015_n4405));
   BUFCHD FE_PHC5085_n2623 (.O(FE_PHN5085_n2623), 
	.I(FE_PHN5788_n2623));
   BUFCHD FE_PHC5084_n3049 (.O(FE_PHN5084_n3049), 
	.I(FE_PHN5888_n3049));
   BUFCKMHD FE_PHC5083_n3217 (.O(FE_PHN5083_n3217), 
	.I(FE_PHN4179_n3217));
   BUFCHD FE_PHC5082_n4263 (.O(FE_PHN5082_n4263), 
	.I(FE_PHN5944_n4263));
   BUFCKEHD FE_PHC5081_n954 (.O(FE_PHN5081_n954), 
	.I(FE_PHN5782_n954));
   BUFCHD FE_PHC5080_n3056 (.O(FE_PHN5080_n3056), 
	.I(FE_PHN6014_n3056));
   BUFCKMHD FE_PHC5079_n1886 (.O(FE_PHN5079_n1886), 
	.I(FE_PHN3437_n1886));
   BUFCHD FE_PHC5078_n1034 (.O(FE_PHN5078_n1034), 
	.I(FE_PHN5872_n1034));
   BUFCHD FE_PHC5077_n1026 (.O(FE_PHN5077_n1026), 
	.I(FE_PHN6133_n1026));
   BUFCHD FE_PHC5076_n891 (.O(FE_PHN5076_n891), 
	.I(FE_PHN5797_n891));
   BUFCHD FE_PHC5075_n4006 (.O(FE_PHN5075_n4006), 
	.I(FE_PHN6056_n4006));
   BUFCHD FE_PHC5074_ram_145__10_ (.O(FE_PHN5074_ram_145__10_), 
	.I(FE_PHN6034_ram_145__10_));
   BUFCKEHD FE_PHC5073_n1873 (.O(FE_PHN5073_n1873), 
	.I(FE_PHN5784_n1873));
   BUFCHD FE_PHC5072_n3071 (.O(FE_PHN5072_n3071), 
	.I(FE_PHN5846_n3071));
   BUFCHD FE_PHC5071_n3988 (.O(FE_PHN5071_n3988), 
	.I(FE_PHN5844_n3988));
   BUFCKMHD FE_PHC5070_n4289 (.O(FE_PHN5070_n4289), 
	.I(FE_PHN6224_n4289));
   BUFCKGHD FE_PHC5069_n1022 (.O(FE_PHN5069_n1022), 
	.I(FE_PHN5853_n1022));
   BUFCKIHD FE_PHC5068_n1051 (.O(FE_PHN5068_n1051), 
	.I(FE_PHN3686_n1051));
   BUFCHD FE_PHC5067_n2956 (.O(FE_PHN5067_n2956), 
	.I(FE_PHN5848_n2956));
   BUFCHD FE_PHC5066_n855 (.O(FE_PHN5066_n855), 
	.I(FE_PHN5902_n855));
   BUFCHD FE_PHC5065_n4010 (.O(FE_PHN5065_n4010), 
	.I(FE_PHN6007_n4010));
   BUFCKEHD FE_PHC5064_n2421 (.O(FE_PHN5064_n2421), 
	.I(FE_PHN5819_n2421));
   BUFCHD FE_PHC5063_n2383 (.O(FE_PHN5063_n2383), 
	.I(FE_PHN5816_n2383));
   BUFCHD FE_PHC5062_n2900 (.O(FE_PHN5062_n2900), 
	.I(FE_PHN5828_n2900));
   BUFCHD FE_PHC5061_n4385 (.O(FE_PHN5061_n4385), 
	.I(FE_PHN5875_n4385));
   BUFCKMHD FE_PHC5060_n4111 (.O(FE_PHN5060_n4111), 
	.I(FE_PHN6099_n4111));
   BUFCKLHD FE_PHC5059_n2430 (.O(FE_PHN5059_n2430), 
	.I(FE_PHN5973_n2430));
   BUFCHD FE_PHC5058_n4407 (.O(FE_PHN5058_n4407), 
	.I(FE_PHN5813_n4407));
   BUFCKMHD FE_PHC5057_n947 (.O(FE_PHN5057_n947), 
	.I(FE_PHN6245_n947));
   BUFCHD FE_PHC5056_n1905 (.O(FE_PHN5056_n1905), 
	.I(FE_PHN5795_n1905));
   BUFCKMHD FE_PHC5055_n1904 (.O(FE_PHN5055_n1904), 
	.I(FE_PHN6437_n1904));
   BUFCKMHD FE_PHC5054_n919 (.O(FE_PHN5054_n919), 
	.I(FE_PHN6241_n919));
   BUFCKMHD FE_PHC5053_n952 (.O(FE_PHN5053_n952), 
	.I(FE_PHN6365_n952));
   BUFCHD FE_PHC5052_n2955 (.O(FE_PHN5052_n2955), 
	.I(FE_PHN5854_n2955));
   BUFCKMHD FE_PHC5051_n4271 (.O(FE_PHN5051_n4271), 
	.I(FE_PHN6146_n4271));
   BUFCHD FE_PHC5050_n4410 (.O(FE_PHN5050_n4410), 
	.I(FE_PHN5821_n4410));
   BUFCKMHD FE_PHC5049_n4356 (.O(FE_PHN5049_n4356), 
	.I(FE_PHN6338_n4356));
   BUFCHD FE_PHC5048_n4359 (.O(FE_PHN5048_n4359), 
	.I(FE_PHN5818_n4359));
   BUFCHD FE_PHC5047_n2958 (.O(FE_PHN5047_n2958), 
	.I(FE_PHN5886_n2958));
   BUFCHD FE_PHC5046_ram_144__8_ (.O(FE_PHN5046_ram_144__8_), 
	.I(FE_PHN5878_ram_144__8_));
   BUFCHD FE_PHC5045_n1088 (.O(FE_PHN5045_n1088), 
	.I(FE_PHN6158_n1088));
   BUFCHD FE_PHC5044_n2437 (.O(FE_PHN5044_n2437), 
	.I(FE_PHN5814_n2437));
   BUFCHD FE_PHC5043_n857 (.O(FE_PHN5043_n857), 
	.I(FE_PHN5912_n857));
   BUFCHD FE_PHC5042_n4421 (.O(FE_PHN5042_n4421), 
	.I(FE_PHN5927_n4421));
   BUFCKMHD FE_PHC5041_n951 (.O(FE_PHN5041_n951), 
	.I(FE_PHN6394_n951));
   BUFCHD FE_PHC5040_n920 (.O(FE_PHN5040_n920), 
	.I(FE_PHN5779_n920));
   BUFCHD FE_PHC5039_n3930 (.O(FE_PHN5039_n3930), 
	.I(FE_PHN5847_n3930));
   BUFCHD FE_PHC5038_n1025 (.O(FE_PHN5038_n1025), 
	.I(FE_PHN6046_n1025));
   BUFCHD FE_PHC5037_n2433 (.O(FE_PHN5037_n2433), 
	.I(FE_PHN5798_n2433));
   BUFCHD FE_PHC5036_n3077 (.O(FE_PHN5036_n3077), 
	.I(FE_PHN5780_n3077));
   BUFCHD FE_PHC5035_n2399 (.O(FE_PHN5035_n2399), 
	.I(FE_PHN5801_n2399));
   BUFCHD FE_PHC5034_n872 (.O(FE_PHN5034_n872), 
	.I(FE_PHN5810_n872));
   BUFCKMHD FE_PHC5033_n904 (.O(FE_PHN5033_n904), 
	.I(FE_PHN6436_n904));
   BUFCHD FE_PHC5032_n4324 (.O(FE_PHN5032_n4324), 
	.I(FE_PHN5914_n4324));
   BUFCHD FE_PHC5031_n1056 (.O(FE_PHN5031_n1056), 
	.I(FE_PHN5900_n1056));
   BUFCKKHD FE_PHC5030_n4372 (.O(FE_PHN5030_n4372), 
	.I(FE_PHN6277_n4372));
   BUFCHD FE_PHC5029_n4036 (.O(FE_PHN5029_n4036), 
	.I(FE_PHN5817_n4036));
   BUFCKMHD FE_PHC5028_n1916 (.O(FE_PHN5028_n1916), 
	.I(FE_PHN6267_n1916));
   BUFCHD FE_PHC5027_n3978 (.O(FE_PHN5027_n3978), 
	.I(FE_PHN5965_n3978));
   BUFCHD FE_PHC5026_n4001 (.O(FE_PHN5026_n4001), 
	.I(FE_PHN5826_n4001));
   BUFCHD FE_PHC5025_n4017 (.O(FE_PHN5025_n4017), 
	.I(FE_PHN5892_n4017));
   BUFCHD FE_PHC5024_n3010 (.O(FE_PHN5024_n3010), 
	.I(FE_PHN5987_n3010));
   BUFCKEHD FE_PHC5023_n2431 (.O(FE_PHN5023_n2431), 
	.I(FE_PHN5785_n2431));
   BUFCHD FE_PHC5022_n851 (.O(FE_PHN5022_n851), 
	.I(FE_PHN5869_n851));
   BUFCHD FE_PHC5021_n4362 (.O(FE_PHN5021_n4362), 
	.I(FE_PHN5815_n4362));
   BUFCHD FE_PHC5020_n998 (.O(FE_PHN5020_n998), 
	.I(FE_PHN6032_n998));
   BUFCKMHD FE_PHC5019_n2703 (.O(FE_PHN5019_n2703), 
	.I(FE_PHN6347_n2703));
   BUFCHD FE_PHC5018_n1008 (.O(FE_PHN5018_n1008), 
	.I(FE_PHN6254_n1008));
   BUFCHD FE_PHC5017_n3128 (.O(FE_PHN5017_n3128), 
	.I(FE_PHN5966_n3128));
   BUFCKLHD FE_PHC5016_n2374 (.O(FE_PHN5016_n2374), 
	.I(FE_PHN3486_n2374));
   BUFCHD FE_PHC5015_n2389 (.O(FE_PHN5015_n2389), 
	.I(FE_PHN5799_n2389));
   BUFCHD FE_PHC5014_n4399 (.O(FE_PHN5014_n4399), 
	.I(FE_PHN5949_n4399));
   BUFCKMHD FE_PHC5013_n2952 (.O(FE_PHN5013_n2952), 
	.I(FE_PHN6242_n2952));
   BUFCKMHD FE_PHC5012_n3223 (.O(FE_PHN5012_n3223), 
	.I(FE_PHN6322_n3223));
   BUFCKLHD FE_PHC5011_n4375 (.O(FE_PHN5011_n4375), 
	.I(FE_PHN6354_n4375));
   BUFCHD FE_PHC5010_n4387 (.O(FE_PHN5010_n4387), 
	.I(FE_PHN5855_n4387));
   BUFCHD FE_PHC5009_n3927 (.O(FE_PHN5009_n3927), 
	.I(FE_PHN5870_n3927));
   BUFCHD FE_PHC5008_n4307 (.O(FE_PHN5008_n4307), 
	.I(FE_PHN5876_n4307));
   BUFCHD FE_PHC5007_n4033 (.O(FE_PHN5007_n4033), 
	.I(FE_PHN5934_n4033));
   BUFCHD FE_PHC5006_n1032 (.O(FE_PHN5006_n1032), 
	.I(FE_PHN6082_n1032));
   BUFCHD FE_PHC5005_n2967 (.O(FE_PHN5005_n2967), 
	.I(FE_PHN5783_n2967));
   BUFCHD FE_PHC5004_n1045 (.O(FE_PHN5004_n1045), 
	.I(FE_PHN6002_n1045));
   BUFCKMHD FE_PHC5003_n4146 (.O(FE_PHN5003_n4146), 
	.I(FE_PHN6421_n4146));
   BUFCKMHD FE_PHC5002_n4332 (.O(FE_PHN5002_n4332), 
	.I(FE_PHN6039_n4332));
   BUFCKKHD FE_PHC5001_n4379 (.O(FE_PHN5001_n4379), 
	.I(FE_PHN6004_n4379));
   BUFCHD FE_PHC5000_n984 (.O(FE_PHN5000_n984), 
	.I(FE_PHN6100_n984));
   BUFCHD FE_PHC4999_n2977 (.O(FE_PHN4999_n2977), 
	.I(FE_PHN6130_n2977));
   BUFCHD FE_PHC4998_n2994 (.O(FE_PHN4998_n2994), 
	.I(FE_PHN6008_n2994));
   BUFCHD FE_PHC4997_n3994 (.O(FE_PHN4997_n3994), 
	.I(FE_PHN5889_n3994));
   BUFCHD FE_PHC4996_n4005 (.O(FE_PHN4996_n4005), 
	.I(FE_PHN5830_n4005));
   BUFCHD FE_PHC4995_n4371 (.O(FE_PHN4995_n4371), 
	.I(FE_PHN5809_n4371));
   BUFCHD FE_PHC4994_n2981 (.O(FE_PHN4994_n2981), 
	.I(FE_PHN6103_n2981));
   BUFCHD FE_PHC4993_n4000 (.O(FE_PHN4993_n4000), 
	.I(FE_PHN5789_n4000));
   BUFCHD FE_PHC4992_n4343 (.O(FE_PHN4992_n4343), 
	.I(FE_PHN5793_n4343));
   BUFCKMHD FE_PHC4991_n3947 (.O(FE_PHN4991_n3947), 
	.I(FE_PHN6353_n3947));
   BUFCKKHD FE_PHC4990_n2953 (.O(FE_PHN4990_n2953), 
	.I(FE_PHN6065_n2953));
   BUFCHD FE_PHC4989_n3073 (.O(FE_PHN4989_n3073), 
	.I(FE_PHN5835_n3073));
   BUFCHD FE_PHC4988_n1087 (.O(FE_PHN4988_n1087), 
	.I(FE_PHN5837_n1087));
   BUFCHD FE_PHC4987_n2415 (.O(FE_PHN4987_n2415), 
	.I(FE_PHN5781_n2415));
   BUFCHD FE_PHC4986_n2978 (.O(FE_PHN4986_n2978), 
	.I(FE_PHN5977_n2978));
   BUFCHD FE_PHC4985_n4022 (.O(FE_PHN4985_n4022), 
	.I(FE_PHN6090_n4022));
   BUFCKMHD FE_PHC4984_n2966 (.O(FE_PHN4984_n2966), 
	.I(FE_PHN6327_n2966));
   BUFCHD FE_PHC4983_n2979 (.O(FE_PHN4983_n2979), 
	.I(FE_PHN6127_n2979));
   BUFCKMHD FE_PHC4982_n958 (.O(FE_PHN4982_n958), 
	.I(FE_PHN6314_n958));
   BUFCHD FE_PHC4981_n4389 (.O(FE_PHN4981_n4389), 
	.I(FE_PHN5959_n4389));
   BUFCKGHD FE_PHC4980_n2408 (.O(FE_PHN4980_n2408), 
	.I(FE_PHN5790_n2408));
   BUFCKMHD FE_PHC4979_n961 (.O(FE_PHN4979_n961), 
	.I(FE_PHN6081_n961));
   BUFCKEHD FE_PHC4978_n928 (.O(FE_PHN4978_n928), 
	.I(FE_PHN5778_n928));
   BUFCHD FE_PHC4977_n1093 (.O(FE_PHN4977_n1093), 
	.I(FE_PHN5863_n1093));
   BUFCKMHD FE_PHC4976_n960 (.O(FE_PHN4976_n960), 
	.I(FE_PHN6274_n960));
   BUFCKMHD FE_PHC4975_n2906 (.O(FE_PHN4975_n2906), 
	.I(FE_PHN6408_n2906));
   BUFCKMHD FE_PHC4974_n1921 (.O(FE_PHN4974_n1921), 
	.I(FE_PHN6265_n1921));
   BUFCKMHD FE_PHC4973_n3931 (.O(FE_PHN4973_n3931), 
	.I(FE_PHN6374_n3931));
   BUFCHD FE_PHC4972_n2961 (.O(FE_PHN4972_n2961), 
	.I(FE_PHN5981_n2961));
   BUFCKMHD FE_PHC4971_ram_98__3_ (.O(FE_PHN4971_ram_98__3_), 
	.I(FE_PHN6427_ram_98__3_));
   BUFCHD FE_PHC4970_n2962 (.O(FE_PHN4970_n2962), 
	.I(FE_PHN5931_n2962));
   BUFCHD FE_PHC4969_n1090 (.O(FE_PHN4969_n1090), 
	.I(FE_PHN5918_n1090));
   BUFCKMHD FE_PHC4968_n3265 (.O(FE_PHN4968_n3265), 
	.I(FE_PHN6400_n3265));
   BUFCKMHD FE_PHC4967_n3999 (.O(FE_PHN4967_n3999), 
	.I(FE_PHN6407_n3999));
   BUFCHD FE_PHC4966_n970 (.O(FE_PHN4966_n970), 
	.I(FE_PHN6070_n970));
   BUFCHD FE_PHC4965_n1048 (.O(FE_PHN4965_n1048), 
	.I(FE_PHN6060_n1048));
   BUFCHD FE_PHC4964_n4009 (.O(FE_PHN4964_n4009), 
	.I(FE_PHN5995_n4009));
   BUFCKMHD FE_PHC4963_n899 (.O(FE_PHN4963_n899), 
	.I(FE_PHN3487_n899));
   BUFCHD FE_PHC4962_n1078 (.O(FE_PHN4962_n1078), 
	.I(FE_PHN5796_n1078));
   BUFCHD FE_PHC4961_n4323 (.O(FE_PHN4961_n4323), 
	.I(FE_PHN5829_n4323));
   BUFEHD FE_PHC4960_n3150 (.O(FE_PHN4960_n3150), 
	.I(n3150));
   BUFCKMHD FE_PHC4959_n1913 (.O(FE_PHN4959_n1913), 
	.I(n1913));
   BUFEHD FE_PHC4958_n4002 (.O(FE_PHN4958_n4002), 
	.I(n4002));
   BUFIHD FE_PHC4957_n1019 (.O(FE_PHN4957_n1019), 
	.I(n1019));
   BUFEHD FE_PHC4956_n2155 (.O(FE_PHN4956_n2155), 
	.I(n2155));
   BUFCKEHD FE_PHC4955_n2154 (.O(FE_PHN4955_n2154), 
	.I(n2154));
   BUFCKEHD FE_PHC4954_n2257 (.O(FE_PHN4954_n2257), 
	.I(n2257));
   BUFCKMHD FE_PHC4953_n2577 (.O(FE_PHN4953_n2577), 
	.I(FE_PHN5775_n2577));
   BUFEHD FE_PHC4952_n2740 (.O(FE_PHN4952_n2740), 
	.I(n2740));
   BUFCKEHD FE_PHC4951_n1086 (.O(FE_PHN4951_n1086), 
	.I(n1086));
   BUFEHD FE_PHC4950_n2126 (.O(FE_PHN4950_n2126), 
	.I(n2126));
   BUFCKMHD FE_PHC4949_n1865 (.O(FE_PHN4949_n1865), 
	.I(n1865));
   BUFKHD FE_PHC4948_n2172 (.O(FE_PHN4948_n2172), 
	.I(n2172));
   BUFNHD FE_PHC4947_n2406 (.O(FE_PHN4947_n2406), 
	.I(FE_PHN5773_n2406));
   BUFCKMHD FE_PHC4946_n921 (.O(FE_PHN4946_n921), 
	.I(n921));
   BUFKHD FE_PHC4945_n2251 (.O(FE_PHN4945_n2251), 
	.I(n2251));
   BUFCKMHD FE_PHC4944_n3017 (.O(FE_PHN4944_n3017), 
	.I(FE_PHN5776_n3017));
   BUFNHD FE_PHC4943_n1012 (.O(FE_PHN4943_n1012), 
	.I(n1012));
   BUFEHD FE_PHC4942_n4102 (.O(FE_PHN4942_n4102), 
	.I(n4102));
   BUFJHD FE_PHC4941_n2747 (.O(FE_PHN4941_n2747), 
	.I(n2747));
   BUFHHD FE_PHC4940_n2615 (.O(FE_PHN4940_n2615), 
	.I(n2615));
   BUFEHD FE_PHC4939_n1178 (.O(FE_PHN4939_n1178), 
	.I(n1178));
   BUFEHD FE_PHC4938_n2133 (.O(FE_PHN4938_n2133), 
	.I(n2133));
   BUFCHD FE_PHC4937_n3021 (.O(FE_PHN4937_n3021), 
	.I(FE_PHN6584_n3021));
   BUFNHD FE_PHC4936_n2414 (.O(FE_PHN4936_n2414), 
	.I(n2414));
   BUFLHD FE_PHC4935_n973 (.O(FE_PHN4935_n973), 
	.I(n973));
   BUFEHD FE_PHC4934_n1190 (.O(FE_PHN4934_n1190), 
	.I(n1190));
   BUFCKMHD FE_PHC4933_n1908 (.O(FE_PHN4933_n1908), 
	.I(n1908));
   BUFKHD FE_PHC4932_n2181 (.O(FE_PHN4932_n2181), 
	.I(n2181));
   BUFHHD FE_PHC4931_n2622 (.O(FE_PHN4931_n2622), 
	.I(n2622));
   BUFCHD FE_PHC4930_n2610 (.O(FE_PHN4930_n2610), 
	.I(FE_PHN7263_n2610));
   BUFLHD FE_PHC4929_n1028 (.O(FE_PHN4929_n1028), 
	.I(n1028));
   BUFEHD FE_PHC4928_n967 (.O(FE_PHN4928_n967), 
	.I(n967));
   BUFEHD FE_PHC4927_n2625 (.O(FE_PHN4927_n2625), 
	.I(n2625));
   BUFEHD FE_PHC4926_n2177 (.O(FE_PHN4926_n2177), 
	.I(n2177));
   BUFEHD FE_PHC4925_n1286 (.O(FE_PHN4925_n1286), 
	.I(n1286));
   BUFCKEHD FE_PHC4924_n2743 (.O(FE_PHN4924_n2743), 
	.I(n2743));
   BUFEHD FE_PHC4923_n2696 (.O(FE_PHN4923_n2696), 
	.I(n2696));
   BUFCHD FE_PHC4922_n2180 (.O(FE_PHN4922_n2180), 
	.I(FE_PHN6709_n2180));
   BUFCHD FE_PHC4921_n2175 (.O(FE_PHN4921_n2175), 
	.I(n2175));
   BUFHHD FE_PHC4920_n977 (.O(FE_PHN4920_n977), 
	.I(n977));
   BUFEHD FE_PHC4919_n1863 (.O(FE_PHN4919_n1863), 
	.I(n1863));
   BUFEHD FE_PHC4918_n2750 (.O(FE_PHN4918_n2750), 
	.I(n2750));
   BUFNHD FE_PHC4917_n2397 (.O(FE_PHN4917_n2397), 
	.I(n2397));
   BUFCKEHD FE_PHC4916_n2876 (.O(FE_PHN4916_n2876), 
	.I(n2876));
   BUFEHD FE_PHC4915_n2566 (.O(FE_PHN4915_n2566), 
	.I(n2566));
   BUFIHD FE_PHC4914_n2125 (.O(FE_PHN4914_n2125), 
	.I(n2125));
   BUFCHD FE_PHC4913_n2873 (.O(FE_PHN4913_n2873), 
	.I(n2873));
   BUFLHD FE_PHC4912_n2611 (.O(FE_PHN4912_n2611), 
	.I(n2611));
   BUFEHD FE_PHC4911_n2857 (.O(FE_PHN4911_n2857), 
	.I(n2857));
   BUFEHD FE_PHC4910_n2590 (.O(FE_PHN4910_n2590), 
	.I(n2590));
   BUFCKEHD FE_PHC4909_n2119 (.O(FE_PHN4909_n2119), 
	.I(n2119));
   BUFEHD FE_PHC4908_n2378 (.O(FE_PHN4908_n2378), 
	.I(n2378));
   BUFNHD FE_PHC4907_n1003 (.O(FE_PHN4907_n1003), 
	.I(n1003));
   BUFNHD FE_PHC4906_n2624 (.O(FE_PHN4906_n2624), 
	.I(n2624));
   BUFMHD FE_PHC4905_n2381 (.O(FE_PHN4905_n2381), 
	.I(n2381));
   BUFCHD FE_PHC4904_n981 (.O(FE_PHN4904_n981), 
	.I(FE_PHN6581_n981));
   BUFCKEHD FE_PHC4903_n4147 (.O(FE_PHN4903_n4147), 
	.I(n4147));
   BUFIHD FE_PHC4902_n1031 (.O(FE_PHN4902_n1031), 
	.I(n1031));
   BUFNHD FE_PHC4901_n2619 (.O(FE_PHN4901_n2619), 
	.I(FE_PHN5767_n2619));
   BUFCHD FE_PHC4900_n2123 (.O(FE_PHN4900_n2123), 
	.I(n2123));
   BUFNHD FE_PHC4899_n2921 (.O(FE_PHN4899_n2921), 
	.I(n2921));
   BUFEHD FE_PHC4898_n979 (.O(FE_PHN4898_n979), 
	.I(n979));
   BUFLHD FE_PHC4897_n2919 (.O(FE_PHN4897_n2919), 
	.I(n2919));
   BUFCKEHD FE_PHC4896_n2749 (.O(FE_PHN4896_n2749), 
	.I(n2749));
   BUFEHD FE_PHC4895_n2434 (.O(FE_PHN4895_n2434), 
	.I(n2434));
   BUFCHD FE_PHC4894_n996 (.O(FE_PHN4894_n996), 
	.I(FE_PHN6559_n996));
   BUFCKEHD FE_PHC4893_n1054 (.O(FE_PHN4893_n1054), 
	.I(n1054));
   BUFJHD FE_PHC4892_n2594 (.O(FE_PHN4892_n2594), 
	.I(n2594));
   BUFCHD FE_PHC4891_n1007 (.O(FE_PHN4891_n1007), 
	.I(FE_PHN5743_n1007));
   BUFCHD FE_PHC4890_n2603 (.O(FE_PHN4890_n2603), 
	.I(n2603));
   BUFHHD FE_PHC4889_n2614 (.O(FE_PHN4889_n2614), 
	.I(n2614));
   BUFCHD FE_PHC4888_n2890 (.O(FE_PHN4888_n2890), 
	.I(FE_PHN6706_n2890));
   BUFCKEHD FE_PHC4887_n2589 (.O(FE_PHN4887_n2589), 
	.I(n2589));
   BUFCKEHD FE_PHC4886_n2159 (.O(FE_PHN4886_n2159), 
	.I(n2159));
   BUFIHD FE_PHC4885_n2572 (.O(FE_PHN4885_n2572), 
	.I(n2572));
   BUFEHD FE_PHC4884_n2161 (.O(FE_PHN4884_n2161), 
	.I(n2161));
   BUFKHD FE_PHC4883_n2576 (.O(FE_PHN4883_n2576), 
	.I(n2576));
   BUFCKEHD FE_PHC4882_n1001 (.O(FE_PHN4882_n1001), 
	.I(FE_PHN5712_n1001));
   BUFIHD FE_PHC4881_n2423 (.O(FE_PHN4881_n2423), 
	.I(n2423));
   BUFEHD FE_PHC4880_n2570 (.O(FE_PHN4880_n2570), 
	.I(n2570));
   BUFNHD FE_PHC4879_n2697 (.O(FE_PHN4879_n2697), 
	.I(n2697));
   BUFCHD FE_PHC4878_n4107 (.O(FE_PHN4878_n4107), 
	.I(n4107));
   BUFCHD FE_PHC4877_n4013 (.O(FE_PHN4877_n4013), 
	.I(FE_PHN6702_n4013));
   BUFEHD FE_PHC4876_n1015 (.O(FE_PHN4876_n1015), 
	.I(n1015));
   BUFNHD FE_PHC4875_n3047 (.O(FE_PHN4875_n3047), 
	.I(FE_PHN5772_n3047));
   BUFEHD FE_PHC4874_n2169 (.O(FE_PHN4874_n2169), 
	.I(n2169));
   BUFHHD FE_PHC4873_n3230 (.O(FE_PHN4873_n3230), 
	.I(n3230));
   BUFCKMHD FE_PHC4872_n1375 (.O(FE_PHN4872_n1375), 
	.I(n1375));
   BUFLHD FE_PHC4871_n1142 (.O(FE_PHN4871_n1142), 
	.I(n1142));
   BUFCHD FE_PHC4870_n2592 (.O(FE_PHN4870_n2592), 
	.I(FE_PHN7220_n2592));
   BUFNHD FE_PHC4869_n2422 (.O(FE_PHN4869_n2422), 
	.I(FE_PHN5769_n2422));
   BUFEHD FE_PHC4868_n2892 (.O(FE_PHN4868_n2892), 
	.I(n2892));
   BUFCHD FE_PHC4867_n985 (.O(FE_PHN4867_n985), 
	.I(FE_PHN5726_n985));
   BUFCHD FE_PHC4866_n2118 (.O(FE_PHN4866_n2118), 
	.I(n2118));
   BUFJHD FE_PHC4865_n2695 (.O(FE_PHN4865_n2695), 
	.I(n2695));
   BUFCKMHD FE_PHC4864_n2889 (.O(FE_PHN4864_n2889), 
	.I(FE_PHN5766_n2889));
   BUFEHD FE_PHC4863_n1154 (.O(FE_PHN4863_n1154), 
	.I(n1154));
   BUFCHD FE_PHC4862_n2604 (.O(FE_PHN4862_n2604), 
	.I(n2604));
   BUFEHD FE_PHC4861_n4139 (.O(FE_PHN4861_n4139), 
	.I(n4139));
   BUFIHD FE_PHC4860_n2166 (.O(FE_PHN4860_n2166), 
	.I(n2166));
   BUFEHD FE_PHC4859_n2628 (.O(FE_PHN4859_n2628), 
	.I(n2628));
   BUFEHD FE_PHC4858_n2616 (.O(FE_PHN4858_n2616), 
	.I(n2616));
   BUFCHD FE_PHC4857_n4114 (.O(FE_PHN4857_n4114), 
	.I(n4114));
   BUFEHD FE_PHC4856_n2701 (.O(FE_PHN4856_n2701), 
	.I(n2701));
   BUFCHD FE_PHC4855_n2609 (.O(FE_PHN4855_n2609), 
	.I(n2609));
   BUFJHD FE_PHC4854_n2376 (.O(FE_PHN4854_n2376), 
	.I(n2376));
   BUFCHD FE_PHC4853_n2402 (.O(FE_PHN4853_n2402), 
	.I(n2402));
   BUFHHD FE_PHC4852_n2612 (.O(FE_PHN4852_n2612), 
	.I(n2612));
   BUFHHD FE_PHC4851_n2120 (.O(FE_PHN4851_n2120), 
	.I(n2120));
   BUFCHD FE_PHC4850_n2379 (.O(FE_PHN4850_n2379), 
	.I(n2379));
   BUFNHD FE_PHC4849_n2626 (.O(FE_PHN4849_n2626), 
	.I(n2626));
   BUFNHD FE_PHC4848_n2386 (.O(FE_PHN4848_n2386), 
	.I(n2386));
   BUFCHD FE_PHC4847_n2582 (.O(FE_PHN4847_n2582), 
	.I(FE_PHN6673_n2582));
   BUFCKEHD FE_PHC4846_n4155 (.O(FE_PHN4846_n4155), 
	.I(n4155));
   BUFCHD FE_PHC4845_n2132 (.O(FE_PHN4845_n2132), 
	.I(n2132));
   BUFLHD FE_PHC4844_n1094 (.O(FE_PHN4844_n1094), 
	.I(n1094));
   BUFEHD FE_PHC4843_n2578 (.O(FE_PHN4843_n2578), 
	.I(n2578));
   BUFCHD FE_PHC4842_n2144 (.O(FE_PHN4842_n2144), 
	.I(FE_PHN6552_n2144));
   BUFLHD FE_PHC4841_n2893 (.O(FE_PHN4841_n2893), 
	.I(n2893));
   BUFCKEHD FE_PHC4840_n2165 (.O(FE_PHN4840_n2165), 
	.I(n2165));
   BUFCKEHD FE_PHC4839_n2426 (.O(FE_PHN4839_n2426), 
	.I(n2426));
   BUFIHD FE_PHC4838_n953 (.O(FE_PHN4838_n953), 
	.I(n953));
   BUFEHD FE_PHC4837_n2375 (.O(FE_PHN4837_n2375), 
	.I(n2375));
   BUFCHD FE_PHC4836_n1158 (.O(FE_PHN4836_n1158), 
	.I(FE_PHN5697_n1158));
   BUFCKMHD FE_PHC4835_n4135 (.O(FE_PHN4835_n4135), 
	.I(n4135));
   BUFIHD FE_PHC4834_n980 (.O(FE_PHN4834_n980), 
	.I(n980));
   BUFJHD FE_PHC4833_n2424 (.O(FE_PHN4833_n2424), 
	.I(n2424));
   BUFCHD FE_PHC4832_n4137 (.O(FE_PHN4832_n4137), 
	.I(FE_PHN6701_n4137));
   BUFIHD FE_PHC4831_n3981 (.O(FE_PHN4831_n3981), 
	.I(n3981));
   BUFEHD FE_PHC4830_n2382 (.O(FE_PHN4830_n2382), 
	.I(n2382));
   BUFEHD FE_PHC4829_n2427 (.O(FE_PHN4829_n2427), 
	.I(n2427));
   BUFHHD FE_PHC4828_n2124 (.O(FE_PHN4828_n2124), 
	.I(n2124));
   BUFCHD FE_PHC4827_n2377 (.O(FE_PHN4827_n2377), 
	.I(n2377));
   BUFCKEHD FE_PHC4826_n2122 (.O(FE_PHN4826_n2122), 
	.I(n2122));
   BUFIHD FE_PHC4825_n2138 (.O(FE_PHN4825_n2138), 
	.I(n2138));
   BUFEHD FE_PHC4824_n2152 (.O(FE_PHN4824_n2152), 
	.I(n2152));
   BUFEHD FE_PHC4823_n2137 (.O(FE_PHN4823_n2137), 
	.I(n2137));
   BUFEHD FE_PHC4822_n2121 (.O(FE_PHN4822_n2121), 
	.I(n2121));
   BUFJHD FE_PHC4821_n2156 (.O(FE_PHN4821_n2156), 
	.I(n2156));
   BUFNHD FE_PHC4820_n2587 (.O(FE_PHN4820_n2587), 
	.I(n2587));
   BUFEHD FE_PHC4819_n2571 (.O(FE_PHN4819_n2571), 
	.I(n2571));
   BUFNHD FE_PHC4818_n4150 (.O(FE_PHN4818_n4150), 
	.I(n4150));
   BUFCKMHD FE_PHC4817_n3033 (.O(FE_PHN4817_n3033), 
	.I(FE_PHN5774_n3033));
   BUFEHD FE_PHC4816_n2135 (.O(FE_PHN4816_n2135), 
	.I(n2135));
   BUFMHD FE_PHC4815_n2618 (.O(FE_PHN4815_n2618), 
	.I(n2618));
   BUFNHD FE_PHC4814_n2390 (.O(FE_PHN4814_n2390), 
	.I(n2390));
   BUFEHD FE_PHC4813_n2171 (.O(FE_PHN4813_n2171), 
	.I(n2171));
   BUFCHD FE_PHC4812_n2429 (.O(FE_PHN4812_n2429), 
	.I(n2429));
   BUFNHD FE_PHC4811_n2398 (.O(FE_PHN4811_n2398), 
	.I(n2398));
   BUFCKMHD FE_PHC4810_n2938 (.O(FE_PHN4810_n2938), 
	.I(FE_PHN5768_n2938));
   BUFCKEHD FE_PHC4809_n2170 (.O(FE_PHN4809_n2170), 
	.I(n2170));
   BUFNHD FE_PHC4808_n2908 (.O(FE_PHN4808_n2908), 
	.I(n2908));
   BUFEHD FE_PHC4807_n2407 (.O(FE_PHN4807_n2407), 
	.I(n2407));
   BUFJHD FE_PHC4806_n2148 (.O(FE_PHN4806_n2148), 
	.I(n2148));
   BUFCKMHD FE_PHC4805_n4151 (.O(FE_PHN4805_n4151), 
	.I(n4151));
   BUFCHD FE_PHC4804_n2887 (.O(FE_PHN4804_n2887), 
	.I(FE_PHN6704_n2887));
   BUFCHD FE_PHC4803_n2410 (.O(FE_PHN4803_n2410), 
	.I(n2410));
   BUFEHD FE_PHC4802_n2393 (.O(FE_PHN4802_n2393), 
	.I(n2393));
   BUFCHD FE_PHC4801_n2417 (.O(FE_PHN4801_n2417), 
	.I(FE_PHN6665_n2417));
   BUFEHD FE_PHC4800_n2411 (.O(FE_PHN4800_n2411), 
	.I(n2411));
   BUFLHD FE_PHC4799_n2907 (.O(FE_PHN4799_n2907), 
	.I(n2907));
   BUFEHD FE_PHC4798_n2401 (.O(FE_PHN4798_n2401), 
	.I(n2401));
   BUFJHD FE_PHC4797_n2380 (.O(FE_PHN4797_n2380), 
	.I(n2380));
   BUFCKEHD FE_PHC4796_n2176 (.O(FE_PHN4796_n2176), 
	.I(n2176));
   BUFIHD FE_PHC4795_n2167 (.O(FE_PHN4795_n2167), 
	.I(n2167));
   BUFLHD FE_PHC4794_n983 (.O(FE_PHN4794_n983), 
	.I(n983));
   BUFLHD FE_PHC4793_n2602 (.O(FE_PHN4793_n2602), 
	.I(n2602));
   BUFHHD FE_PHC4792_n2394 (.O(FE_PHN4792_n2394), 
	.I(n2394));
   BUFCKEHD FE_PHC4791_n2151 (.O(FE_PHN4791_n2151), 
	.I(n2151));
   BUFCKEHD FE_PHC4790_n2425 (.O(FE_PHN4790_n2425), 
	.I(n2425));
   BUFCKEHD FE_PHC4789_n2164 (.O(FE_PHN4789_n2164), 
	.I(n2164));
   BUFIHD FE_PHC4788_n2149 (.O(FE_PHN4788_n2149), 
	.I(n2149));
   BUFCKEHD FE_PHC4787_n4011 (.O(FE_PHN4787_n4011), 
	.I(n4011));
   BUFLHD FE_PHC4786_n2941 (.O(FE_PHN4786_n2941), 
	.I(n2941));
   BUFCHD FE_PHC4785_n2179 (.O(FE_PHN4785_n2179), 
	.I(FE_PHN6695_n2179));
   BUFMHD FE_PHC4784_n4012 (.O(FE_PHN4784_n4012), 
	.I(n4012));
   BUFMHD FE_PHC4783_n2925 (.O(FE_PHN4783_n2925), 
	.I(n2925));
   BUFCKEHD FE_PHC4782_n4163 (.O(FE_PHN4782_n4163), 
	.I(n4163));
   BUFJHD FE_PHC4781_n2412 (.O(FE_PHN4781_n2412), 
	.I(n2412));
   BUFCKEHD FE_PHC4780_n4153 (.O(FE_PHN4780_n4153), 
	.I(n4153));
   BUFCHD FE_PHC4779_n2130 (.O(FE_PHN4779_n2130), 
	.I(FE_PHN7214_n2130));
   BUFCKEHD FE_PHC4778_n2395 (.O(FE_PHN4778_n2395), 
	.I(n2395));
   BUFCKEHD FE_PHC4777_n4121 (.O(FE_PHN4777_n4121), 
	.I(n4121));
   BUFJHD FE_PHC4776_n4018 (.O(FE_PHN4776_n4018), 
	.I(n4018));
   BUFCKEHD FE_PHC4775_n2168 (.O(FE_PHN4775_n2168), 
	.I(n2168));
   BUFCKEHD FE_PHC4774_n2428 (.O(FE_PHN4774_n2428), 
	.I(n2428));
   BUFCKEHD FE_PHC4773_n1027 (.O(FE_PHN4773_n1027), 
	.I(FE_PHN5644_n1027));
   BUFCKEHD FE_PHC4772_n2413 (.O(FE_PHN4772_n2413), 
	.I(FE_PHN5621_n2413));
   BUFCKEHD FE_PHC4771_n1062 (.O(FE_PHN4771_n1062), 
	.I(FE_PHN5619_n1062));
   BUFCKEHD FE_PHC4770_n4123 (.O(FE_PHN4770_n4123), 
	.I(FE_PHN5635_n4123));
   BUFCKEHD FE_PHC4769_n2262 (.O(FE_PHN4769_n2262), 
	.I(FE_PHN6425_n2262));
   BUFCKEHD FE_PHC4768_n2127 (.O(FE_PHN4768_n2127), 
	.I(FE_PHN5605_n2127));
   BUFCKEHD FE_PHC4767_n1068 (.O(FE_PHN4767_n1068), 
	.I(FE_PHN5609_n1068));
   BUFCKEHD FE_PHC4766_n2926 (.O(FE_PHN4766_n2926), 
	.I(FE_PHN5618_n2926));
   BUFCKEHD FE_PHC4765_n2258 (.O(FE_PHN4765_n2258), 
	.I(FE_PHN5608_n2258));
   BUFCKEHD FE_PHC4764_n971 (.O(FE_PHN4764_n971), 
	.I(FE_PHN5626_n971));
   BUFCKEHD FE_PHC4763_n2158 (.O(FE_PHN4763_n2158), 
	.I(FE_PHN5604_n2158));
   BUFCKEHD FE_PHC4762_n2923 (.O(FE_PHN4762_n2923), 
	.I(FE_PHN5646_n2923));
   BUFCKEHD FE_PHC4761_n2396 (.O(FE_PHN4761_n2396), 
	.I(FE_PHN5603_n2396));
   BUFCKEHD FE_PHC4760_n2141 (.O(FE_PHN4760_n2141), 
	.I(FE_PHN5597_n2141));
   BUFCKEHD FE_PHC4759_n2733 (.O(FE_PHN4759_n2733), 
	.I(FE_PHN5643_n2733));
   BUFCKEHD FE_PHC4758_n2605 (.O(FE_PHN4758_n2605), 
	.I(FE_PHN5640_n2605));
   BUFCKEHD FE_PHC4757_n2732 (.O(FE_PHN4757_n2732), 
	.I(FE_PHN5642_n2732));
   BUFCKEHD FE_PHC4756_n2727 (.O(FE_PHN4756_n2727), 
	.I(FE_PHN5645_n2727));
   BUFCKEHD FE_PHC4755_n3241 (.O(FE_PHN4755_n3241), 
	.I(FE_PHN6417_n3241));
   BUFCHD FE_PHC4754_n1206 (.O(FE_PHN4754_n1206), 
	.I(FE_PHN6399_n1206));
   BUFCKEHD FE_PHC4753_n4175 (.O(FE_PHN4753_n4175), 
	.I(FE_PHN5630_n4175));
   BUFCKEHD FE_PHC4752_n2600 (.O(FE_PHN4752_n2600), 
	.I(FE_PHN5631_n2600));
   BUFCHD FE_PHC4751_n4170 (.O(FE_PHN4751_n4170), 
	.I(FE_PHN6393_n4170));
   BUFCKEHD FE_PHC4750_n1046 (.O(FE_PHN4750_n1046), 
	.I(FE_PHN5629_n1046));
   BUFCHD FE_PHC4749_n2391 (.O(FE_PHN4749_n2391), 
	.I(FE_PHN5623_n2391));
   BUFCHD FE_PHC4748_n3920 (.O(FE_PHN4748_n3920), 
	.I(FE_PHN6364_n3920));
   BUFCHD FE_PHC4747_n2910 (.O(FE_PHN4747_n2910), 
	.I(FE_PHN5613_n2910));
   BUFCHD FE_PHC4746_n4015 (.O(FE_PHN4746_n4015), 
	.I(FE_PHN5627_n4015));
   BUFCHD FE_PHC4745_n4094 (.O(FE_PHN4745_n4094), 
	.I(FE_PHN6304_n4094));
   BUFCHD FE_PHC4744_n4097 (.O(FE_PHN4744_n4097), 
	.I(FE_PHN5598_n4097));
   BUFCHD FE_PHC4743_n3950 (.O(FE_PHN4743_n3950), 
	.I(FE_PHN5600_n3950));
   BUFCHD FE_PHC4742_n2990 (.O(FE_PHN4742_n2990), 
	.I(FE_PHN5592_n2990));
   BUFCHD FE_PHC4741_n3917 (.O(FE_PHN4741_n3917), 
	.I(FE_PHN5594_n3917));
   BUFCHD FE_PHC4740_n4265 (.O(FE_PHN4740_n4265), 
	.I(FE_PHN5586_n4265));
   BUFCHD FE_PHC4739_n4076 (.O(FE_PHN4739_n4076), 
	.I(FE_PHN5591_n4076));
   BUFCHD FE_PHC4738_n3951 (.O(FE_PHN4738_n3951), 
	.I(FE_PHN5576_n3951));
   BUFCHD FE_PHC4737_n3936 (.O(FE_PHN4737_n3936), 
	.I(FE_PHN5567_n3936));
   BUFCHD FE_PHC4736_n4236 (.O(FE_PHN4736_n4236), 
	.I(FE_PHN5564_n4236));
   BUFCHD FE_PHC4735_n3952 (.O(FE_PHN4735_n3952), 
	.I(FE_PHN5577_n3952));
   BUFCHD FE_PHC4734_n873 (.O(FE_PHN4734_n873), 
	.I(FE_PHN5566_n873));
   BUFCHD FE_PHC4733_n4366 (.O(FE_PHN4733_n4366), 
	.I(FE_PHN5556_n4366));
   BUFCHD FE_PHC4732_n4395 (.O(FE_PHN4732_n4395), 
	.I(FE_PHN5515_n4395));
   BUFCHD FE_PHC4731_n3135 (.O(FE_PHN4731_n3135), 
	.I(FE_PHN5572_n3135));
   BUFCHD FE_PHC4730_n4267 (.O(FE_PHN4730_n4267), 
	.I(FE_PHN5589_n4267));
   BUFCHD FE_PHC4729_n4420 (.O(FE_PHN4729_n4420), 
	.I(FE_PHN5509_n4420));
   BUFCHD FE_PHC4728_n2974 (.O(FE_PHN4728_n2974), 
	.I(FE_PHN5500_n2974));
   DELAKHD FE_PHC4727_n4087 (.O(FE_PHN4727_n4087), 
	.I(FE_PHN3499_n4087));
   DELCKHD FE_PHC4726_n4207 (.O(FE_PHN4726_n4207), 
	.I(FE_PHN3773_n4207));
   BUFCHD FE_PHC4725_n3008 (.O(FE_PHN4725_n3008), 
	.I(FE_PHN5539_n3008));
   BUFCHD FE_PHC4724_n3940 (.O(FE_PHN4724_n3940), 
	.I(FE_PHN5531_n3940));
   BUFCHD FE_PHC4723_n3062 (.O(FE_PHN4723_n3062), 
	.I(FE_PHN5548_n3062));
   BUFCHD FE_PHC4722_n838 (.O(FE_PHN4722_n838), 
	.I(FE_PHN5553_n838));
   BUFCHD FE_PHC4721_n4235 (.O(FE_PHN4721_n4235), 
	.I(FE_PHN5580_n4235));
   BUFCHD FE_PHC4720_n2957 (.O(FE_PHN4720_n2957), 
	.I(FE_PHN5542_n2957));
   BUFCHD FE_PHC4719_n4262 (.O(FE_PHN4719_n4262), 
	.I(FE_PHN5519_n4262));
   BUFCHD FE_PHC4718_n4233 (.O(FE_PHN4718_n4233), 
	.I(FE_PHN5536_n4233));
   BUFCHD FE_PHC4717_n3038 (.O(FE_PHN4717_n3038), 
	.I(FE_PHN5565_n3038));
   BUFCHD FE_PHC4716_n4171 (.O(FE_PHN4716_n4171), 
	.I(FE_PHN5496_n4171));
   BUFCHD FE_PHC4715_n3956 (.O(FE_PHN4715_n3956), 
	.I(FE_PHN5521_n3956));
   BUFCHD FE_PHC4714_n4202 (.O(FE_PHN4714_n4202), 
	.I(FE_PHN5478_n4202));
   BUFCHD FE_PHC4713_n4414 (.O(FE_PHN4713_n4414), 
	.I(FE_PHN5495_n4414));
   BUFCHD FE_PHC4712_n2928 (.O(FE_PHN4712_n2928), 
	.I(FE_PHN5507_n2928));
   BUFCHD FE_PHC4711_n863 (.O(FE_PHN4711_n863), 
	.I(FE_PHN5550_n863));
   BUFCHD FE_PHC4710_n2918 (.O(FE_PHN4710_n2918), 
	.I(FE_PHN5505_n2918));
   BUFCHD FE_PHC4709_n2886 (.O(FE_PHN4709_n2886), 
	.I(FE_PHN5508_n2886));
   BUFCHD FE_PHC4708_n3210 (.O(FE_PHN4708_n3210), 
	.I(FE_PHN5436_n3210));
   BUFCHD FE_PHC4707_n895 (.O(FE_PHN4707_n895), 
	.I(FE_PHN5540_n895));
   BUFCHD FE_PHC4706_n4329 (.O(FE_PHN4706_n4329), 
	.I(FE_PHN5461_n4329));
   BUFCHD FE_PHC4705_n1066 (.O(FE_PHN4705_n1066), 
	.I(FE_PHN5471_n1066));
   BUFCHD FE_PHC4704_n4215 (.O(FE_PHN4704_n4215), 
	.I(FE_PHN5440_n4215));
   BUFCHD FE_PHC4703_n4240 (.O(FE_PHN4703_n4240), 
	.I(FE_PHN5443_n4240));
   BUFCHD FE_PHC4702_n2943 (.O(FE_PHN4702_n2943), 
	.I(FE_PHN5442_n2943));
   BUFCHD FE_PHC4701_n2920 (.O(FE_PHN4701_n2920), 
	.I(FE_PHN5485_n2920));
   BUFCHD FE_PHC4700_n4209 (.O(FE_PHN4700_n4209), 
	.I(FE_PHN5391_n4209));
   BUFCHD FE_PHC4699_n892 (.O(FE_PHN4699_n892), 
	.I(FE_PHN5432_n892));
   BUFCHD FE_PHC4698_n839 (.O(FE_PHN4698_n839), 
	.I(FE_PHN5438_n839));
   BUFCHD FE_PHC4697_n854 (.O(FE_PHN4697_n854), 
	.I(FE_PHN5489_n854));
   BUFCHD FE_PHC4696_n843 (.O(FE_PHN4696_n843), 
	.I(FE_PHN5483_n843));
   BUFCHD FE_PHC4695_n4402 (.O(FE_PHN4695_n4402), 
	.I(FE_PHN5339_n4402));
   BUFCHD FE_PHC4694_n2564 (.O(FE_PHN4694_n2564), 
	.I(FE_PHN5357_n2564));
   BUFCHD FE_PHC4693_n2888 (.O(FE_PHN4693_n2888), 
	.I(FE_PHN5405_n2888));
   BUFCHD FE_PHC4692_n3126 (.O(FE_PHN4692_n3126), 
	.I(FE_PHN5435_n3126));
   BUFCHD FE_PHC4691_n3916 (.O(FE_PHN4691_n3916), 
	.I(FE_PHN5415_n3916));
   BUFCHD FE_PHC4690_n4276 (.O(FE_PHN4690_n4276), 
	.I(FE_PHN5488_n4276));
   BUFCHD FE_PHC4689_n4164 (.O(FE_PHN4689_n4164), 
	.I(FE_PHN5420_n4164));
   BUFCHD FE_PHC4688_n880 (.O(FE_PHN4688_n880), 
	.I(FE_PHN6545_n880));
   BUFCHD FE_PHC4687_n896 (.O(FE_PHN4687_n896), 
	.I(FE_PHN6568_n896));
   BUFCHD FE_PHC4686_n3258 (.O(FE_PHN4686_n3258), 
	.I(FE_PHN5403_n3258));
   BUFCHD FE_PHC4685_n4178 (.O(FE_PHN4685_n4178), 
	.I(FE_PHN5868_n4178));
   BUFCHD FE_PHC4684_n4226 (.O(FE_PHN4684_n4226), 
	.I(FE_PHN5369_n4226));
   BUFCHD FE_PHC4683_n4311 (.O(FE_PHN4683_n4311), 
	.I(FE_PHN5349_n4311));
   BUFCHD FE_PHC4682_n4222 (.O(FE_PHN4682_n4222), 
	.I(FE_PHN5390_n4222));
   BUFCHD FE_PHC4681_n911 (.O(FE_PHN4681_n911), 
	.I(FE_PHN5381_n911));
   BUFCHD FE_PHC4680_n4210 (.O(FE_PHN4680_n4210), 
	.I(FE_PHN6542_n4210));
   BUFCHD FE_PHC4679_n886 (.O(FE_PHN4679_n886), 
	.I(FE_PHN5467_n886));
   BUFCHD FE_PHC4678_n3109 (.O(FE_PHN4678_n3109), 
	.I(FE_PHN5529_n3109));
   BUFCHD FE_PHC4677_n4046 (.O(FE_PHN4677_n4046), 
	.I(FE_PHN5337_n4046));
   BUFCKEHD FE_PHC4676_n966 (.O(FE_PHN4676_n966), 
	.I(n966));
   BUFCHD FE_PHC4675_n2970 (.O(FE_PHN4675_n2970), 
	.I(FE_PHN5347_n2970));
   BUFCHD FE_PHC4674_n3980 (.O(FE_PHN4674_n3980), 
	.I(FE_PHN6531_n3980));
   BUFCHD FE_PHC4673_n874 (.O(FE_PHN4673_n874), 
	.I(FE_PHN5469_n874));
   BUFCHD FE_PHC4672_n2297 (.O(FE_PHN4672_n2297), 
	.I(FE_PHN6252_n2297));
   BUFCHD FE_PHC4671_n2580 (.O(FE_PHN4671_n2580), 
	.I(FE_PHN5348_n2580));
   BUFCKEHD FE_PHC4670_n3932 (.O(FE_PHN4670_n3932), 
	.I(FE_PHN6521_n3932));
   BUFCHD FE_PHC4669_n3924 (.O(FE_PHN4669_n3924), 
	.I(FE_PHN5295_n3924));
   BUFCHD FE_PHC4668_n4029 (.O(FE_PHN4668_n4029), 
	.I(FE_PHN5383_n4029));
   BUFCHD FE_PHC4667_n903 (.O(FE_PHN4667_n903), 
	.I(FE_PHN5358_n903));
   BUFCHD FE_PHC4666_n2916 (.O(FE_PHN4666_n2916), 
	.I(FE_PHN5379_n2916));
   BUFCHD FE_PHC4665_n4412 (.O(FE_PHN4665_n4412), 
	.I(FE_PHN5462_n4412));
   BUFCHD FE_PHC4664_n1920 (.O(FE_PHN4664_n1920), 
	.I(FE_PHN5262_n1920));
   BUFCHD FE_PHC4663_n962 (.O(FE_PHN4663_n962), 
	.I(FE_PHN6525_n962));
   BUFCHD FE_PHC4662_n3976 (.O(FE_PHN4662_n3976), 
	.I(FE_PHN5421_n3976));
   BUFCHD FE_PHC4661_n4299 (.O(FE_PHN4661_n4299), 
	.I(FE_PHN5299_n4299));
   BUFCHD FE_PHC4660_n4364 (.O(FE_PHN4660_n4364), 
	.I(FE_PHN5394_n4364));
   BUFCHD FE_PHC4659_n3086 (.O(FE_PHN4659_n3086), 
	.I(FE_PHN5329_n3086));
   BUFCHD FE_PHC4658_n3131 (.O(FE_PHN4658_n3131), 
	.I(FE_PHN5322_n3131));
   BUFCHD FE_PHC4657_n3945 (.O(FE_PHN4657_n3945), 
	.I(FE_PHN6543_n3945));
   BUFCHD FE_PHC4656_n3044 (.O(FE_PHN4656_n3044), 
	.I(FE_PHN5464_n3044));
   BUFCHD FE_PHC4655_n2420 (.O(FE_PHN4655_n2420), 
	.I(FE_PHN5361_n2420));
   BUFCHD FE_PHC4654_n2984 (.O(FE_PHN4654_n2984), 
	.I(FE_PHN5363_n2984));
   BUFCHD FE_PHC4653_n3964 (.O(FE_PHN4653_n3964), 
	.I(FE_PHN5368_n3964));
   BUFCHD FE_PHC4652_n3255 (.O(FE_PHN4652_n3255), 
	.I(FE_PHN5380_n3255));
   BUFCHD FE_PHC4651_n2936 (.O(FE_PHN4651_n2936), 
	.I(FE_PHN5282_n2936));
   BUFCHD FE_PHC4650_n4392 (.O(FE_PHN4650_n4392), 
	.I(FE_PHN5398_n4392));
   BUFCHD FE_PHC4649_n4281 (.O(FE_PHN4649_n4281), 
	.I(FE_PHN5318_n4281));
   BUFCHD FE_PHC4648_n2963 (.O(FE_PHN4648_n2963), 
	.I(FE_PHN5525_n2963));
   BUFCHD FE_PHC4647_n850 (.O(FE_PHN4647_n850), 
	.I(FE_PHN5446_n850));
   BUFCHD FE_PHC4646_n3028 (.O(FE_PHN4646_n3028), 
	.I(FE_PHN5399_n3028));
   BUFCHD FE_PHC4645_n2965 (.O(FE_PHN4645_n2965), 
	.I(FE_PHN5510_n2965));
   BUFCHD FE_PHC4644_n2950 (.O(FE_PHN4644_n2950), 
	.I(FE_PHN5320_n2950));
   BUFMHD FE_PHC4643_n4227 (.O(FE_PHN4643_n4227), 
	.I(n4227));
   BUFCHD FE_PHC4642_n4284 (.O(FE_PHN4642_n4284), 
	.I(FE_PHN5332_n4284));
   BUFCHD FE_PHC4641_n3098 (.O(FE_PHN4641_n3098), 
	.I(FE_PHN5328_n3098));
   BUFCHD FE_PHC4640_n4368 (.O(FE_PHN4640_n4368), 
	.I(FE_PHN5345_n4368));
   BUFCHD FE_PHC4639_n3020 (.O(FE_PHN4639_n3020), 
	.I(FE_PHN5210_n3020));
   BUFCHD FE_PHC4638_n4396 (.O(FE_PHN4638_n4396), 
	.I(FE_PHN5375_n4396));
   BUFMHD FE_PHC4637_n4187 (.O(FE_PHN4637_n4187), 
	.I(n4187));
   BUFCHD FE_PHC4636_n1106 (.O(FE_PHN4636_n1106), 
	.I(n1106));
   BUFCKLHD FE_PHC4635_n4268 (.O(FE_PHN4635_n4268), 
	.I(FE_PHN5617_n4268));
   BUFLHD FE_PHC4634_n2944 (.O(FE_PHN4634_n2944), 
	.I(n2944));
   BUFCHD FE_PHC4633_n4212 (.O(FE_PHN4633_n4212), 
	.I(FE_PHN5411_n4212));
   BUFCHD FE_PHC4632_n3130 (.O(FE_PHN4632_n3130), 
	.I(FE_PHN5384_n3130));
   BUFCHD FE_PHC4631_n4252 (.O(FE_PHN4631_n4252), 
	.I(FE_PHN5324_n4252));
   BUFCHD FE_PHC4630_n2987 (.O(FE_PHN4630_n2987), 
	.I(FE_PHN5245_n2987));
   BUFCHD FE_PHC4629_n3040 (.O(FE_PHN4629_n3040), 
	.I(FE_PHN5401_n3040));
   BUFCKEHD FE_PHC4628_n898 (.O(FE_PHN4628_n898), 
	.I(FE_PHN6533_n898));
   BUFCHD FE_PHC4627_n3136 (.O(FE_PHN4627_n3136), 
	.I(FE_PHN5338_n3136));
   BUFCHD FE_PHC4626_n1870 (.O(FE_PHN4626_n1870), 
	.I(FE_PHN5241_n1870));
   BUFIHD FE_PHC4625_n1042 (.O(FE_PHN4625_n1042), 
	.I(FE_PHN3999_n1042));
   BUFCHD FE_PHC4624_n1014 (.O(FE_PHN4624_n1014), 
	.I(FE_PHN5377_n1014));
   BUFCHD FE_PHC4623_n4049 (.O(FE_PHN4623_n4049), 
	.I(FE_PHN5263_n4049));
   BUFCHD FE_PHC4622_n969 (.O(FE_PHN4622_n969), 
	.I(FE_PHN5396_n969));
   BUFCHD FE_PHC4621_n1023 (.O(FE_PHN4621_n1023), 
	.I(FE_PHN5490_n1023));
   BUFCHD FE_PHC4620_n4278 (.O(FE_PHN4620_n4278), 
	.I(FE_PHN5257_n4278));
   BUFCHD FE_PHC4619_n4241 (.O(FE_PHN4619_n4241), 
	.I(FE_PHN5154_n4241));
   BUFGHD FE_PHC4618_n4172 (.O(FE_PHN4618_n4172), 
	.I(FE_PHN5364_n4172));
   BUFCHD FE_PHC4617_n2927 (.O(FE_PHN4617_n2927), 
	.I(FE_PHN5256_n2927));
   BUFEHD FE_PHC4616_n4416 (.O(FE_PHN4616_n4416), 
	.I(FE_PHN5310_n4416));
   BUFCHD FE_PHC4615_n4016 (.O(FE_PHN4615_n4016), 
	.I(FE_PHN6526_n4016));
   BUFCKEHD FE_PHC4614_n1922 (.O(FE_PHN4614_n1922), 
	.I(n1922));
   BUFCHD FE_PHC4613_n3958 (.O(FE_PHN4613_n3958), 
	.I(FE_PHN5327_n3958));
   BUFCHD FE_PHC4612_n2983 (.O(FE_PHN4612_n2983), 
	.I(FE_PHN5160_n2983));
   BUFCHD FE_PHC4611_n935 (.O(FE_PHN4611_n935), 
	.I(FE_PHN5251_n935));
   BUFCHD FE_PHC4610_n4179 (.O(FE_PHN4610_n4179), 
	.I(FE_PHN6202_n4179));
   BUFCHD FE_PHC4609_n1874 (.O(FE_PHN4609_n1874), 
	.I(FE_PHN7063_n1874));
   BUFCKGHD FE_PHC4608_n2986 (.O(FE_PHN4608_n2986), 
	.I(FE_PHN5416_n2986));
   BUFCHD FE_PHC4607_n993 (.O(FE_PHN4607_n993), 
	.I(FE_PHN5407_n993));
   BUFCHD FE_PHC4606_n1021 (.O(FE_PHN4606_n1021), 
	.I(FE_PHN5419_n1021));
   BUFCHD FE_PHC4605_n841 (.O(FE_PHN4605_n841), 
	.I(FE_PHN5236_n841));
   BUFCKLHD FE_PHC4604_n4219 (.O(FE_PHN4604_n4219), 
	.I(FE_PHN5456_n4219));
   BUFCHD FE_PHC4603_n2722 (.O(FE_PHN4603_n2722), 
	.I(FE_PHN5240_n2722));
   BUFCHD FE_PHC4602_n2384 (.O(FE_PHN4602_n2384), 
	.I(FE_PHN5254_n2384));
   BUFCHD FE_PHC4601_n877 (.O(FE_PHN4601_n877), 
	.I(FE_PHN5452_n877));
   BUFCHD FE_PHC4600_n2405 (.O(FE_PHN4600_n2405), 
	.I(FE_PHN5290_n2405));
   BUFIHD FE_PHC4599_n3058 (.O(FE_PHN4599_n3058), 
	.I(FE_PHN3873_n3058));
   BUFCHD FE_PHC4598_n3015 (.O(FE_PHN4598_n3015), 
	.I(FE_PHN5370_n3015));
   BUFCHD FE_PHC4597_n4232 (.O(FE_PHN4597_n4232), 
	.I(FE_PHN5238_n4232));
   BUFCHD FE_PHC4596_n2891 (.O(FE_PHN4596_n2891), 
	.I(FE_PHN5207_n2891));
   BUFNHD FE_PHC4595_n1020 (.O(FE_PHN4595_n1020), 
	.I(n1020));
   BUFCHD FE_PHC4594_n3962 (.O(FE_PHN4594_n3962), 
	.I(FE_PHN6515_n3962));
   BUFCHD FE_PHC4593_n910 (.O(FE_PHN4593_n910), 
	.I(FE_PHN5196_n910));
   BUFCHD FE_PHC4592_n878 (.O(FE_PHN4592_n878), 
	.I(FE_PHN5188_n878));
   BUFCHD FE_PHC4591_n3139 (.O(FE_PHN4591_n3139), 
	.I(FE_PHN5455_n3139));
   BUFCKLHD FE_PHC4590_n889 (.O(FE_PHN4590_n889), 
	.I(n889));
   BUFCKLHD FE_PHC4589_n4231 (.O(FE_PHN4589_n4231), 
	.I(FE_PHN5599_n4231));
   BUFCHD FE_PHC4588_n847 (.O(FE_PHN4588_n847), 
	.I(FE_PHN5437_n847));
   BUFCHD FE_PHC4587_n858 (.O(FE_PHN4587_n858), 
	.I(FE_PHN5346_n858));
   BUFCHD FE_PHC4586_n1110 (.O(FE_PHN4586_n1110), 
	.I(FE_PHN5994_n1110));
   BUFCHD FE_PHC4585_n975 (.O(FE_PHN4585_n975), 
	.I(FE_PHN5283_n975));
   BUFCHD FE_PHC4584_n3082 (.O(FE_PHN4584_n3082), 
	.I(FE_PHN5244_n3082));
   BUFCHD FE_PHC4583_n4021 (.O(FE_PHN4583_n4021), 
	.I(FE_PHN5199_n4021));
   BUFCHD FE_PHC4582_n2574 (.O(FE_PHN4582_n2574), 
	.I(FE_PHN5246_n2574));
   BUFCHD FE_PHC4581_n948 (.O(FE_PHN4581_n948), 
	.I(FE_PHN5209_n948));
   BUFCHD FE_PHC4580_n3257 (.O(FE_PHN4580_n3257), 
	.I(FE_PHN5284_n3257));
   BUFCHD FE_PHC4579_n2989 (.O(FE_PHN4579_n2989), 
	.I(FE_PHN5194_n2989));
   BUFCKEHD FE_PHC4578_n3052 (.O(FE_PHN4578_n3052), 
	.I(FE_PHN5179_n3052));
   BUFCKGHD FE_PHC4577_n991 (.O(FE_PHN4577_n991), 
	.I(FE_PHN5414_n991));
   BUFCHD FE_PHC4576_n4316 (.O(FE_PHN4576_n4316), 
	.I(FE_PHN5232_n4316));
   BUFCHD FE_PHC4575_n882 (.O(FE_PHN4575_n882), 
	.I(FE_PHN5400_n882));
   BUFCHD FE_PHC4574_n4228 (.O(FE_PHN4574_n4228), 
	.I(FE_PHN5463_n4228));
   BUFCKMHD FE_PHC4573_n4181 (.O(FE_PHN4573_n4181), 
	.I(FE_PHN5633_n4181));
   BUFCHD FE_PHC4572_n4259 (.O(FE_PHN4572_n4259), 
	.I(FE_PHN6519_n4259));
   BUFCKEHD FE_PHC4571_n2388 (.O(FE_PHN4571_n2388), 
	.I(FE_PHN6494_n2388));
   BUFCHD FE_PHC4570_n4169 (.O(FE_PHN4570_n4169), 
	.I(FE_PHN5454_n4169));
   BUFCHD FE_PHC4569_n4211 (.O(FE_PHN4569_n4211), 
	.I(FE_PHN5418_n4211));
   BUFCHD FE_PHC4568_n4277 (.O(FE_PHN4568_n4277), 
	.I(FE_PHN5258_n4277));
   BUFCKEHD FE_PHC4567_n4401 (.O(FE_PHN4567_n4401), 
	.I(FE_PHN5127_n4401));
   BUFCKEHD FE_PHC4566_n1018 (.O(FE_PHN4566_n1018), 
	.I(n1018));
   BUFCHD FE_PHC4565_n986 (.O(FE_PHN4565_n986), 
	.I(FE_PHN5433_n986));
   BUFCKNHD FE_PHC4564_n2554 (.O(FE_PHN4564_n2554), 
	.I(FE_PHN5636_n2554));
   BUFCKJHD FE_PHC4563_n2992 (.O(FE_PHN4563_n2992), 
	.I(n2992));
   BUFCHD FE_PHC4562_n4203 (.O(FE_PHN4562_n4203), 
	.I(FE_PHN5298_n4203));
   BUFCHD FE_PHC4561_n4243 (.O(FE_PHN4561_n4243), 
	.I(FE_PHN5130_n4243));
   BUFCHD FE_PHC4560_n913 (.O(FE_PHN4560_n913), 
	.I(FE_PHN5287_n913));
   BUFHHD FE_PHC4559_n3219 (.O(FE_PHN4559_n3219), 
	.I(FE_PHN3916_n3219));
   BUFHHD FE_PHC4558_n4183 (.O(FE_PHN4558_n4183), 
	.I(FE_PHN3898_n4183));
   BUFCHD FE_PHC4557_n905 (.O(FE_PHN4557_n905), 
	.I(FE_PHN5268_n905));
   DELBKHD FE_PHC4556_n1143 (.O(FE_PHN4556_n1143), 
	.I(FE_PHN4002_n1143));
   BUFNHD FE_PHC4555_n3918 (.O(FE_PHN4555_n3918), 
	.I(n3918));
   BUFMHD FE_PHC4554_n4382 (.O(FE_PHN4554_n4382), 
	.I(n4382));
   BUFNHD FE_PHC4553_n869 (.O(FE_PHN4553_n869), 
	.I(n869));
   BUFCHD FE_PHC4552_n4418 (.O(FE_PHN4552_n4418), 
	.I(FE_PHN5334_n4418));
   BUFNHD FE_PHC4551_n3066 (.O(FE_PHN4551_n3066), 
	.I(FE_PHN5616_n3066));
   BUFHHD FE_PHC4550_n3024 (.O(FE_PHN4550_n3024), 
	.I(n3024));
   BUFCHD FE_PHC4549_n1013 (.O(FE_PHN4549_n1013), 
	.I(FE_PHN5307_n1013));
   BUFCHD FE_PHC4548_n4026 (.O(FE_PHN4548_n4026), 
	.I(FE_PHN5453_n4026));
   BUFCHD FE_PHC4547_n4148 (.O(FE_PHN4547_n4148), 
	.I(FE_PHN6458_n4148));
   BUFCHD FE_PHC4546_n3989 (.O(FE_PHN4546_n3989), 
	.I(FE_PHN5388_n3989));
   BUFCHD FE_PHC4545_n968 (.O(FE_PHN4545_n968), 
	.I(FE_PHN5477_n968));
   BUFCHD FE_PHC4544_n2995 (.O(FE_PHN4544_n2995), 
	.I(FE_PHN5389_n2995));
   BUFCKMHD FE_PHC4543_n4168 (.O(FE_PHN4543_n4168), 
	.I(n4168));
   BUFCHD FE_PHC4542_n972 (.O(FE_PHN4542_n972), 
	.I(FE_PHN5255_n972));
   BUFCHD FE_PHC4541_n3119 (.O(FE_PHN4541_n3119), 
	.I(FE_PHN5523_n3119));
   BUFHHD FE_PHC4540_n4255 (.O(FE_PHN4540_n4255), 
	.I(FE_PHN3735_n4255));
   BUFCHD FE_PHC4539_n2971 (.O(FE_PHN4539_n2971), 
	.I(FE_PHN5120_n2971));
   BUFCHD FE_PHC4538_n1872 (.O(FE_PHN4538_n1872), 
	.I(FE_PHN6497_n1872));
   BUFCHD FE_PHC4537_n1037 (.O(FE_PHN4537_n1037), 
	.I(FE_PHN5252_n1037));
   BUFCKGHD FE_PHC4536_n4415 (.O(FE_PHN4536_n4415), 
	.I(n4415));
   BUFCKEHD FE_PHC4535_n3207 (.O(FE_PHN4535_n3207), 
	.I(FE_PHN5261_n3207));
   BUFEHD FE_PHC4534_n2933 (.O(FE_PHN4534_n2933), 
	.I(FE_PHN5153_n2933));
   BUFCKEHD FE_PHC4533_n1082 (.O(FE_PHN4533_n1082), 
	.I(FE_PHN5125_n1082));
   BUFCKJHD FE_PHC4532_n3088 (.O(FE_PHN4532_n3088), 
	.I(FE_PHN5487_n3088));
   BUFCKLHD FE_PHC4531_n3091 (.O(FE_PHN4531_n3091), 
	.I(FE_PHN3576_n3091));
   BUFCHD FE_PHC4530_n4037 (.O(FE_PHN4530_n4037), 
	.I(FE_PHN5216_n4037));
   BUFCHD FE_PHC4529_n2898 (.O(FE_PHN4529_n2898), 
	.I(FE_PHN5457_n2898));
   BUFLHD FE_PHC4528_n2896 (.O(FE_PHN4528_n2896), 
	.I(FE_PHN3858_n2896));
   BUFCHD FE_PHC4527_ram_158__11_ (.O(FE_PHN4527_ram_158__11_), 
	.I(FE_PHN5532_ram_158__11_));
   BUFCHD FE_PHC4526_n4116 (.O(FE_PHN4526_n4116), 
	.I(FE_PHN6464_n4116));
   BUFHHD FE_PHC4525_n3140 (.O(FE_PHN4525_n3140), 
	.I(FE_PHN5378_n3140));
   BUFCHD FE_PHC4524_n3018 (.O(FE_PHN4524_n3018), 
	.I(FE_PHN5150_n3018));
   BUFCKEHD FE_PHC4523_n2954 (.O(FE_PHN4523_n2954), 
	.I(FE_PHN5278_n2954));
   BUFCHD FE_PHC4522_n3942 (.O(FE_PHN4522_n3942), 
	.I(FE_PHN5352_n3942));
   BUFCKEHD FE_PHC4521_n3029 (.O(FE_PHN4521_n3029), 
	.I(FE_PHN3837_n3029));
   BUFLHD FE_PHC4520_n844 (.O(FE_PHN4520_n844), 
	.I(n844));
   BUFCHD FE_PHC4519_n3212 (.O(FE_PHN4519_n3212), 
	.I(FE_PHN6502_n3212));
   BUFCHD FE_PHC4518_n4403 (.O(FE_PHN4518_n4403), 
	.I(FE_PHN6532_n4403));
   BUFCKEHD FE_PHC4517_n999 (.O(FE_PHN4517_n999), 
	.I(FE_PHN5170_n999));
   BUFCHD FE_PHC4516_n4294 (.O(FE_PHN4516_n4294), 
	.I(FE_PHN6507_n4294));
   BUFCHD FE_PHC4515_n4030 (.O(FE_PHN4515_n4030), 
	.I(FE_PHN5353_n4030));
   BUFCHD FE_PHC4514_n3970 (.O(FE_PHN4514_n3970), 
	.I(FE_PHN6493_n3970));
   BUFCHD FE_PHC4513_n2753 (.O(FE_PHN4513_n2753), 
	.I(FE_PHN6201_n2753));
   BUFCHD FE_PHC4512_n3069 (.O(FE_PHN4512_n3069), 
	.I(FE_PHN6138_n3069));
   BUFCKIHD FE_PHC4511_ram_133__9_ (.O(FE_PHN4511_ram_133__9_), 
	.I(FE_PHN3571_ram_133__9_));
   BUFCHD FE_PHC4510_n4394 (.O(FE_PHN4510_n4394), 
	.I(FE_PHN5362_n4394));
   BUFCHD FE_PHC4509_n3065 (.O(FE_PHN4509_n3065), 
	.I(FE_PHN5266_n3065));
   BUFCHD FE_PHC4508_n917 (.O(FE_PHN4508_n917), 
	.I(FE_PHN6516_n917));
   BUFCHD FE_PHC4507_n3137 (.O(FE_PHN4507_n3137), 
	.I(FE_PHN5402_n3137));
   BUFCHD FE_PHC4506_n2385 (.O(FE_PHN4506_n2385), 
	.I(FE_PHN5861_n2385));
   BUFCHD FE_PHC4505_n2996 (.O(FE_PHN4505_n2996), 
	.I(FE_PHN5270_n2996));
   BUFHHD FE_PHC4504_n870 (.O(FE_PHN4504_n870), 
	.I(FE_PHN5147_n870));
   BUFCHD FE_PHC4503_n4229 (.O(FE_PHN4503_n4229), 
	.I(FE_PHN5164_n4229));
   BUFCKMHD FE_PHC4502_n3913 (.O(FE_PHN4502_n3913), 
	.I(FE_PHN5634_n3913));
   BUFCHD FE_PHC4501_n3971 (.O(FE_PHN4501_n3971), 
	.I(FE_PHN6513_n3971));
   BUFCHD FE_PHC4500_n4400 (.O(FE_PHN4500_n4400), 
	.I(FE_PHN5224_n4400));
   BUFCHD FE_PHC4499_n4373 (.O(FE_PHN4499_n4373), 
	.I(FE_PHN5372_n4373));
   BUFCHD FE_PHC4498_n4355 (.O(FE_PHN4498_n4355), 
	.I(FE_PHN5397_n4355));
   BUFCHD FE_PHC4497_n2951 (.O(FE_PHN4497_n2951), 
	.I(FE_PHN5133_n2951));
   BUFCKEHD FE_PHC4496_n4285 (.O(FE_PHN4496_n4285), 
	.I(n4285));
   BUFCHD FE_PHC4495_n4201 (.O(FE_PHN4495_n4201), 
	.I(FE_PHN5458_n4201));
   BUFCHD FE_PHC4494_n1017 (.O(FE_PHN4494_n1017), 
	.I(FE_PHN5187_n1017));
   BUFCKEHD FE_PHC4493_n3072 (.O(FE_PHN4493_n3072), 
	.I(FE_PHN5171_n3072));
   BUFCHD FE_PHC4492_n4308 (.O(FE_PHN4492_n4308), 
	.I(FE_PHN6496_n4308));
   BUFCHD FE_PHC4491_n849 (.O(FE_PHN4491_n849), 
	.I(FE_PHN5342_n849));
   BUFCKIHD FE_PHC4490_n900 (.O(FE_PHN4490_n900), 
	.I(FE_PHN3894_n900));
   BUFCHD FE_PHC4489_n4174 (.O(FE_PHN4489_n4174), 
	.I(FE_PHN5230_n4174));
   BUFCHD FE_PHC4488_n888 (.O(FE_PHN4488_n888), 
	.I(FE_PHN6508_n888));
   BUFCHD FE_PHC4487_n4350 (.O(FE_PHN4487_n4350), 
	.I(FE_PHN5288_n4350));
   BUFCHD FE_PHC4486_n2623 (.O(FE_PHN4486_n2623), 
	.I(FE_PHN5085_n2623));
   BUFCHD FE_PHC4485_n4199 (.O(FE_PHN4485_n4199), 
	.I(FE_PHN5360_n4199));
   BUFCHD FE_PHC4484_n4391 (.O(FE_PHN4484_n4391), 
	.I(FE_PHN6504_n4391));
   BUFCKEHD FE_PHC4483_n2946 (.O(FE_PHN4483_n2946), 
	.I(FE_PHN5331_n2946));
   BUFCHD FE_PHC4482_n3013 (.O(FE_PHN4482_n3013), 
	.I(FE_PHN5417_n3013));
   BUFCHD FE_PHC4481_n4393 (.O(FE_PHN4481_n4393), 
	.I(FE_PHN5205_n4393));
   BUFHHD FE_PHC4480_n879 (.O(FE_PHN4480_n879), 
	.I(n879));
   BUFCKEHD FE_PHC4479_n4360 (.O(FE_PHN4479_n4360), 
	.I(n4360));
   BUFCHD FE_PHC4478_n3076 (.O(FE_PHN4478_n3076), 
	.I(FE_PHN5145_n3076));
   BUFCHD FE_PHC4477_n4188 (.O(FE_PHN4477_n4188), 
	.I(FE_PHN5393_n4188));
   BUFCKEHD FE_PHC4476_n1918 (.O(FE_PHN4476_n1918), 
	.I(FE_PHN6480_n1918));
   BUFNHD FE_PHC4475_n3036 (.O(FE_PHN4475_n3036), 
	.I(FE_PHN5614_n3036));
   BUFCKEHD FE_PHC4474_n944 (.O(FE_PHN4474_n944), 
	.I(FE_PHN6470_n944));
   BUFCHD FE_PHC4473_n4334 (.O(FE_PHN4473_n4334), 
	.I(FE_PHN5167_n4334));
   BUFNHD FE_PHC4472_n4261 (.O(FE_PHN4472_n4261), 
	.I(FE_PHN3699_n4261));
   BUFCHD FE_PHC4471_n2131 (.O(FE_PHN4471_n2131), 
	.I(FE_PHN6498_n2131));
   BUFCKEHD FE_PHC4470_n941 (.O(FE_PHN4470_n941), 
	.I(FE_PHN5325_n941));
   BUFCKMHD FE_PHC4469_n3016 (.O(FE_PHN4469_n3016), 
	.I(FE_PHN5625_n3016));
   BUFCKEHD FE_PHC4468_n936 (.O(FE_PHN4468_n936), 
	.I(FE_PHN3919_n936));
   BUFCHD FE_PHC4467_n897 (.O(FE_PHN4467_n897), 
	.I(FE_PHN5326_n897));
   BUFCHD FE_PHC4466_n2998 (.O(FE_PHN4466_n2998), 
	.I(FE_PHN5321_n2998));
   BUFCHD FE_PHC4465_n3141 (.O(FE_PHN4465_n3141), 
	.I(FE_PHN5439_n3141));
   BUFCHD FE_PHC4464_n4273 (.O(FE_PHN4464_n4273), 
	.I(FE_PHN6488_n4273));
   BUFCKEHD FE_PHC4463_n4419 (.O(FE_PHN4463_n4419), 
	.I(FE_PHN5267_n4419));
   BUFHHD FE_PHC4462_n4300 (.O(FE_PHN4462_n4300), 
	.I(FE_PHN3380_n4300));
   BUFCHD FE_PHC4461_n3963 (.O(FE_PHN4461_n3963), 
	.I(FE_PHN5302_n3963));
   BUFCKEHD FE_PHC4460_n3064 (.O(FE_PHN4460_n3064), 
	.I(n3064));
   BUFCKMHD FE_PHC4459_ram_20__10_ (.O(FE_PHN4459_ram_20__10_), 
	.I(FE_PHN5596_ram_20__10_));
   BUFCKEHD FE_PHC4458_n938 (.O(FE_PHN4458_n938), 
	.I(FE_PHN6479_n938));
   BUFCHD FE_PHC4457_n881 (.O(FE_PHN4457_n881), 
	.I(FE_PHN5271_n881));
   BUFCKMHD FE_PHC4456_n4270 (.O(FE_PHN4456_n4270), 
	.I(FE_PHN5638_n4270));
   BUFCKEHD FE_PHC4455_n1000 (.O(FE_PHN4455_n1000), 
	.I(FE_PHN5434_n1000));
   BUFCHD FE_PHC4454_n965 (.O(FE_PHN4454_n965), 
	.I(FE_PHN5248_n965));
   BUFCHD FE_PHC4453_n4404 (.O(FE_PHN4453_n4404), 
	.I(FE_PHN6489_n4404));
   BUFCHD FE_PHC4452_n997 (.O(FE_PHN4452_n997), 
	.I(FE_PHN5341_n997));
   BUFNHD FE_PHC4451_n4213 (.O(FE_PHN4451_n4213), 
	.I(n4213));
   BUFCKJHD FE_PHC4450_n894 (.O(FE_PHN4450_n894), 
	.I(n894));
   BUFCKEHD FE_PHC4449_n4032 (.O(FE_PHN4449_n4032), 
	.I(FE_PHN4003_n4032));
   BUFCHD FE_PHC4448_n2930 (.O(FE_PHN4448_n2930), 
	.I(FE_PHN5229_n2930));
   BUFCHD FE_PHC4447_n2735 (.O(FE_PHN4447_n2735), 
	.I(FE_PHN5195_n2735));
   BUFCKEHD FE_PHC4446_n3262 (.O(FE_PHN4446_n3262), 
	.I(FE_PHN5105_n3262));
   BUFCKEHD FE_PHC4445_n1034 (.O(FE_PHN4445_n1034), 
	.I(FE_PHN3935_n1034));
   BUFCKGHD FE_PHC4444_n861 (.O(FE_PHN4444_n861), 
	.I(FE_PHN5350_n861));
   BUFCHD FE_PHC4443_n988 (.O(FE_PHN4443_n988), 
	.I(FE_PHN5871_n988));
   BUFCKEHD FE_PHC4442_n2906 (.O(FE_PHN4442_n2906), 
	.I(n2906));
   BUFCKLHD FE_PHC4441_ram_214__13_ (.O(FE_PHN4441_ram_214__13_), 
	.I(FE_PHN3691_ram_214__13_));
   BUFNHD FE_PHC4440_n909 (.O(FE_PHN4440_n909), 
	.I(FE_PHN3619_n909));
   BUFCKLHD FE_PHC4439_n3120 (.O(FE_PHN4439_n3120), 
	.I(FE_PHN5575_n3120));
   BUFCHD FE_PHC4438_n2598 (.O(FE_PHN4438_n2598), 
	.I(FE_PHN6474_n2598));
   BUFCHD FE_PHC4437_n4218 (.O(FE_PHN4437_n4218), 
	.I(FE_PHN6312_n4218));
   BUFCKEHD FE_PHC4436_n2897 (.O(FE_PHN4436_n2897), 
	.I(FE_PHN3766_n2897));
   BUFCKGHD FE_PHC4435_n957 (.O(FE_PHN4435_n957), 
	.I(n957));
   BUFCHD FE_PHC4434_n3985 (.O(FE_PHN4434_n3985), 
	.I(FE_PHN5294_n3985));
   BUFCHD FE_PHC4433_n4166 (.O(FE_PHN4433_n4166), 
	.I(FE_PHN5309_n4166));
   BUFHHD FE_PHC4432_n3919 (.O(FE_PHN4432_n3919), 
	.I(FE_PHN3293_n3919));
   BUFCHD FE_PHC4431_n4185 (.O(FE_PHN4431_n4185), 
	.I(FE_PHN5313_n4185));
   BUFCHD FE_PHC4430_n3910 (.O(FE_PHN4430_n3910), 
	.I(FE_PHN5354_n3910));
   BUFCHD FE_PHC4429_n4180 (.O(FE_PHN4429_n4180), 
	.I(FE_PHN5159_n4180));
   BUFCHD FE_PHC4428_n1030 (.O(FE_PHN4428_n1030), 
	.I(FE_PHN5138_n1030));
   BUFCHD FE_PHC4427_n4194 (.O(FE_PHN4427_n4194), 
	.I(FE_PHN5142_n4194));
   BUFCHD FE_PHC4426_n2599 (.O(FE_PHN4426_n2599), 
	.I(FE_PHN5101_n2599));
   BUFCHD FE_PHC4425_n3969 (.O(FE_PHN4425_n3969), 
	.I(FE_PHN5243_n3969));
   BUFCKEHD FE_PHC4424_n2975 (.O(FE_PHN4424_n2975), 
	.I(FE_PHN5200_n2975));
   BUFCHD FE_PHC4423_n4378 (.O(FE_PHN4423_n4378), 
	.I(FE_PHN5235_n4378));
   BUFCKEHD FE_PHC4422_n2430 (.O(FE_PHN4422_n2430), 
	.I(FE_PHN5059_n2430));
   BUFCKEHD FE_PHC4421_n3075 (.O(FE_PHN4421_n3075), 
	.I(FE_PHN5233_n3075));
   BUFCKEHD FE_PHC4420_n3011 (.O(FE_PHN4420_n3011), 
	.I(FE_PHN5426_n3011));
   BUFCKIHD FE_PHC4419_n3002 (.O(FE_PHN4419_n3002), 
	.I(n3002));
   BUFCKEHD FE_PHC4418_n2403 (.O(FE_PHN4418_n2403), 
	.I(n2403));
   BUFCHD FE_PHC4417_n4206 (.O(FE_PHN4417_n4206), 
	.I(FE_PHN5228_n4206));
   BUFCHD FE_PHC4416_n4017 (.O(FE_PHN4416_n4017), 
	.I(FE_PHN5025_n4017));
   BUFCKEHD FE_PHC4415_n4342 (.O(FE_PHN4415_n4342), 
	.I(n4342));
   BUFCKHHD FE_PHC4414_ram_31__2_ (.O(FE_PHN4414_ram_31__2_), 
	.I(FE_PHN3862_ram_31__2_));
   BUFHHD FE_PHC4413_n3996 (.O(FE_PHN4413_n3996), 
	.I(FE_PHN3259_n3996));
   BUFCHD FE_PHC4412_n4035 (.O(FE_PHN4412_n4035), 
	.I(FE_PHN6500_n4035));
   BUFCHD FE_PHC4411_n1016 (.O(FE_PHN4411_n1016), 
	.I(FE_PHN5365_n1016));
   BUFCKEHD FE_PHC4410_n4370 (.O(FE_PHN4410_n4370), 
	.I(FE_PHN6478_n4370));
   BUFCHD FE_PHC4409_n2997 (.O(FE_PHN4409_n2997), 
	.I(FE_PHN5343_n2997));
   BUFCHD FE_PHC4408_n2959 (.O(FE_PHN4408_n2959), 
	.I(FE_PHN5356_n2959));
   BUFCHD FE_PHC4407_n4266 (.O(FE_PHN4407_n4266), 
	.I(FE_PHN5119_n4266));
   BUFCHD FE_PHC4406_ram_153__11_ (.O(FE_PHN4406_ram_153__11_), 
	.I(FE_PHN5273_ram_153__11_));
   BUFCHD FE_PHC4405_n2993 (.O(FE_PHN4405_n2993), 
	.I(FE_PHN5340_n2993));
   BUFCHD FE_PHC4404_n3006 (.O(FE_PHN4404_n3006), 
	.I(FE_PHN5264_n3006));
   BUFHHD FE_PHC4403_n4338 (.O(FE_PHN4403_n4338), 
	.I(FE_PHN3896_n4338));
   BUFCKEHD FE_PHC4402_n4242 (.O(FE_PHN4402_n4242), 
	.I(FE_PHN6482_n4242));
   BUFCKEHD FE_PHC4401_n2922 (.O(FE_PHN4401_n2922), 
	.I(FE_PHN6452_n2922));
   BUFCHD FE_PHC4400_n1906 (.O(FE_PHN4400_n1906), 
	.I(FE_PHN6481_n1906));
   BUFCKEHD FE_PHC4399_n976 (.O(FE_PHN4399_n976), 
	.I(FE_PHN5385_n976));
   BUFCKMHD FE_PHC4398_n4134 (.O(FE_PHN4398_n4134), 
	.I(n4134));
   BUFCHD FE_PHC4397_n1074 (.O(FE_PHN4397_n1074), 
	.I(FE_PHN5099_n1074));
   BUFCHD FE_PHC4396_n3055 (.O(FE_PHN4396_n3055), 
	.I(FE_PHN5198_n3055));
   BUFCHD FE_PHC4395_n2960 (.O(FE_PHN4395_n2960), 
	.I(FE_PHN5175_n2960));
   BUFCHD FE_PHC4394_n1002 (.O(FE_PHN4394_n1002), 
	.I(FE_PHN5239_n1002));
   BUFCHD FE_PHC4393_n885 (.O(FE_PHN4393_n885), 
	.I(FE_PHN5315_n885));
   BUFCHD FE_PHC4392_n1051 (.O(FE_PHN4392_n1051), 
	.I(FE_PHN5895_n1051));
   BUFCKEHD FE_PHC4391_n4027 (.O(FE_PHN4391_n4027), 
	.I(FE_PHN3742_n4027));
   BUFCHD FE_PHC4390_n4283 (.O(FE_PHN4390_n4283), 
	.I(FE_PHN5336_n4283));
   BUFLHD FE_PHC4389_n2934 (.O(FE_PHN4389_n2934), 
	.I(FE_PHN3253_n2934));
   BUFCHD FE_PHC4388_n3063 (.O(FE_PHN4388_n3063), 
	.I(FE_PHN5183_n3063));
   BUFCKEHD FE_PHC4387_n4271 (.O(FE_PHN4387_n4271), 
	.I(FE_PHN5051_n4271));
   BUFCKLHD FE_PHC4386_n4397 (.O(FE_PHN4386_n4397), 
	.I(FE_PHN5581_n4397));
   BUFCKEHD FE_PHC4385_n3074 (.O(FE_PHN4385_n3074), 
	.I(FE_PHN5218_n3074));
   BUFCHD FE_PHC4384_n3994 (.O(FE_PHN4384_n3994), 
	.I(FE_PHN4997_n3994));
   BUFCHD FE_PHC4383_n3974 (.O(FE_PHN4383_n3974), 
	.I(FE_PHN5158_n3974));
   BUFCHD FE_PHC4382_n3050 (.O(FE_PHN4382_n3050), 
	.I(FE_PHN5185_n3050));
   BUFHHD FE_PHC4381_n3025 (.O(FE_PHN4381_n3025), 
	.I(FE_PHN3891_n3025));
   BUFCKEHD FE_PHC4380_n964 (.O(FE_PHN4380_n964), 
	.I(FE_PHN6477_n964));
   BUFLHD FE_PHC4379_n3080 (.O(FE_PHN4379_n3080), 
	.I(FE_PHN5511_n3080));
   BUFCHD FE_PHC4378_n3992 (.O(FE_PHN4378_n3992), 
	.I(FE_PHN5201_n3992));
   BUFCHD FE_PHC4377_n4358 (.O(FE_PHN4377_n4358), 
	.I(FE_PHN6520_n4358));
   BUFCHD FE_PHC4376_n2945 (.O(FE_PHN4376_n2945), 
	.I(FE_PHN5100_n2945));
   BUFHHD FE_PHC4375_n3927 (.O(FE_PHN4375_n3927), 
	.I(n3927));
   BUFCHD FE_PHC4374_n890 (.O(FE_PHN4374_n890), 
	.I(FE_PHN5204_n890));
   BUFCKHHD FE_PHC4373_n1022 (.O(FE_PHN4373_n1022), 
	.I(n1022));
   BUFCHD FE_PHC4372_n3014 (.O(FE_PHN4372_n3014), 
	.I(FE_PHN5351_n3014));
   BUFCKEHD FE_PHC4371_n1024 (.O(FE_PHN4371_n1024), 
	.I(FE_PHN5371_n1024));
   BUFCKEHD FE_PHC4370_n1880 (.O(FE_PHN4370_n1880), 
	.I(FE_PHN6463_n1880));
   BUFCHD FE_PHC4369_n3263 (.O(FE_PHN4369_n3263), 
	.I(FE_PHN5141_n3263));
   BUFCHD FE_PHC4368_n1009 (.O(FE_PHN4368_n1009), 
	.I(FE_PHN3603_n1009));
   BUFCHD FE_PHC4367_n3921 (.O(FE_PHN4367_n3921), 
	.I(FE_PHN5181_n3921));
   BUFCHD FE_PHC4366_n4411 (.O(FE_PHN4366_n4411), 
	.I(FE_PHN5180_n4411));
   BUFCHD FE_PHC4365_n3961 (.O(FE_PHN4365_n3961), 
	.I(FE_PHN5117_n3961));
   BUFCHD FE_PHC4364_n4217 (.O(FE_PHN4364_n4217), 
	.I(FE_PHN5265_n4217));
   BUFCKEHD FE_PHC4363_n1916 (.O(FE_PHN4363_n1916), 
	.I(FE_PHN5028_n1916));
   BUFCKEHD FE_PHC4362_n4407 (.O(FE_PHN4362_n4407), 
	.I(FE_PHN5058_n4407));
   BUFCKEHD FE_PHC4361_n906 (.O(FE_PHN4361_n906), 
	.I(FE_PHN6476_n906));
   BUFCHD FE_PHC4360_n3122 (.O(FE_PHN4360_n3122), 
	.I(FE_PHN5189_n3122));
   BUFCKEHD FE_PHC4359_n2935 (.O(FE_PHN4359_n2935), 
	.I(FE_PHN3600_n2935));
   BUFCKMHD FE_PHC4358_ram_154__5_ (.O(FE_PHN4358_ram_154__5_), 
	.I(FE_PHN5606_ram_154__5_));
   BUFCKEHD FE_PHC4357_n3049 (.O(FE_PHN4357_n3049), 
	.I(n3049));
   BUFCKMHD FE_PHC4356_n1899 (.O(FE_PHN4356_n1899), 
	.I(FE_PHN5543_n1899));
   BUFCHD FE_PHC4355_n974 (.O(FE_PHN4355_n974), 
	.I(FE_PHN5087_n974));
   BUFCHD FE_PHC4354_n949 (.O(FE_PHN4354_n949), 
	.I(FE_PHN6505_n949));
   BUFCKEHD FE_PHC4353_n2621 (.O(FE_PHN4353_n2621), 
	.I(FE_PHN5110_n2621));
   BUFCKEHD FE_PHC4352_n4333 (.O(FE_PHN4352_n4333), 
	.I(FE_PHN5168_n4333));
   BUFCHD FE_PHC4351_n3093 (.O(FE_PHN4351_n3093), 
	.I(FE_PHN5206_n3093));
   BUFCKEHD FE_PHC4350_n998 (.O(FE_PHN4350_n998), 
	.I(n998));
   BUFCKEHD FE_PHC4349_n3079 (.O(FE_PHN4349_n3079), 
	.I(n3079));
   BUFCKMHD FE_PHC4348_n3129 (.O(FE_PHN4348_n3129), 
	.I(FE_PHN5541_n3129));
   BUFCHD FE_PHC4347_n2421 (.O(FE_PHN4347_n2421), 
	.I(FE_PHN5064_n2421));
   BUFCHD FE_PHC4346_n1029 (.O(FE_PHN4346_n1029), 
	.I(FE_PHN5191_n1029));
   BUFCKEHD FE_PHC4345_n2399 (.O(FE_PHN4345_n2399), 
	.I(FE_PHN3635_n2399));
   BUFCHD FE_PHC4344_n4025 (.O(FE_PHN4344_n4025), 
	.I(FE_PHN5274_n4025));
   BUFCKEHD FE_PHC4343_n2419 (.O(FE_PHN4343_n2419), 
	.I(FE_PHN6467_n2419));
   BUFIHD FE_PHC4342_n1079 (.O(FE_PHN4342_n1079), 
	.I(FE_PHN3842_n1079));
   BUFCKEHD FE_PHC4341_n3975 (.O(FE_PHN4341_n3975), 
	.I(FE_PHN3928_n3975));
   BUFCHD FE_PHC4340_n933 (.O(FE_PHN4340_n933), 
	.I(FE_PHN6468_n933));
   BUFCKEHD FE_PHC4339_n891 (.O(FE_PHN4339_n891), 
	.I(FE_PHN5076_n891));
   BUFCKEHD FE_PHC4338_n904 (.O(FE_PHN4338_n904), 
	.I(FE_PHN3870_n904));
   BUFCKEHD FE_PHC4337_n4036 (.O(FE_PHN4337_n4036), 
	.I(FE_PHN5029_n4036));
   BUFLHD FE_PHC4336_n1006 (.O(FE_PHN4336_n1006), 
	.I(n1006));
   BUFCKJHD FE_PHC4335_n3067 (.O(FE_PHN4335_n3067), 
	.I(n3067));
   BUFHHD FE_PHC4334_n4369 (.O(FE_PHN4334_n4369), 
	.I(FE_PHN3514_n4369));
   BUFCHD FE_PHC4333_n851 (.O(FE_PHN4333_n851), 
	.I(FE_PHN5022_n851));
   BUFCKGHD FE_PHC4332_n3090 (.O(FE_PHN4332_n3090), 
	.I(FE_PHN5374_n3090));
   BUFCHD FE_PHC4331_n853 (.O(FE_PHN4331_n853), 
	.I(FE_PHN5108_n853));
   BUFLHD FE_PHC4330_n845 (.O(FE_PHN4330_n845), 
	.I(FE_PHN3806_n845));
   BUFCKMHD FE_PHC4329_n902 (.O(FE_PHN4329_n902), 
	.I(n902));
   BUFCHD FE_PHC4328_n4374 (.O(FE_PHN4328_n4374), 
	.I(FE_PHN6485_n4374));
   BUFCKEHD FE_PHC4327_n3955 (.O(FE_PHN4327_n3955), 
	.I(FE_PHN6490_n3955));
   BUFCHD FE_PHC4326_n982 (.O(FE_PHN4326_n982), 
	.I(FE_PHN5202_n982));
   BUFCKEHD FE_PHC4325_n4248 (.O(FE_PHN4325_n4248), 
	.I(FE_PHN5102_n4248));
   BUFCHD FE_PHC4324_n840 (.O(FE_PHN4324_n840), 
	.I(FE_PHN5303_n840));
   BUFCHD FE_PHC4323_n3054 (.O(FE_PHN4323_n3054), 
	.I(FE_PHN5220_n3054));
   BUFCHD FE_PHC4322_n3988 (.O(FE_PHN4322_n3988), 
	.I(FE_PHN5071_n3988));
   BUFCHD FE_PHC4321_n2432 (.O(FE_PHN4321_n2432), 
	.I(FE_PHN6444_n2432));
   BUFCHD FE_PHC4320_n3984 (.O(FE_PHN4320_n3984), 
	.I(FE_PHN5155_n3984));
   BUFCKEHD FE_PHC4319_n2163 (.O(FE_PHN4319_n2163), 
	.I(FE_PHN6475_n2163));
   BUFCKMHD FE_PHC4318_n3085 (.O(FE_PHN4318_n3085), 
	.I(FE_PHN5601_n3085));
   BUFCKEHD FE_PHC4317_n2437 (.O(FE_PHN4317_n2437), 
	.I(FE_PHN5044_n2437));
   BUFCHD FE_PHC4316_n4386 (.O(FE_PHN4316_n4386), 
	.I(FE_PHN5090_n4386));
   BUFHHD FE_PHC4315_n994 (.O(FE_PHN4315_n994), 
	.I(FE_PHN3440_n994));
   BUFCKEHD FE_PHC4314_n2904 (.O(FE_PHN4314_n2904), 
	.I(n2904));
   BUFCHD FE_PHC4313_n1026 (.O(FE_PHN4313_n1026), 
	.I(FE_PHN5077_n1026));
   BUFCHD FE_PHC4312_n2988 (.O(FE_PHN4312_n2988), 
	.I(FE_PHN5112_n2988));
   BUFCHD FE_PHC4311_n929 (.O(FE_PHN4311_n929), 
	.I(FE_PHN5223_n929));
   BUFCKEHD FE_PHC4310_n3977 (.O(FE_PHN4310_n3977), 
	.I(FE_PHN5156_n3977));
   BUFCKEHD FE_PHC4309_n954 (.O(FE_PHN4309_n954), 
	.I(FE_PHN5081_n954));
   BUFCHD FE_PHC4308_n4332 (.O(FE_PHN4308_n4332), 
	.I(FE_PHN5002_n4332));
   BUFCKIHD FE_PHC4307_n2754 (.O(FE_PHN4307_n2754), 
	.I(n2754));
   BUFNHD FE_PHC4306_n3005 (.O(FE_PHN4306_n3005), 
	.I(n3005));
   BUFCKEHD FE_PHC4305_n1038 (.O(FE_PHN4305_n1038), 
	.I(FE_PHN3802_n1038));
   BUFCKEHD FE_PHC4304_n2383 (.O(FE_PHN4304_n2383), 
	.I(n2383));
   BUFKHD FE_PHC4303_n3060 (.O(FE_PHN4303_n3060), 
	.I(FE_PHN3841_n3060));
   BUFCHD FE_PHC4302_n2964 (.O(FE_PHN4302_n2964), 
	.I(FE_PHN5225_n2964));
   BUFMHD FE_PHC4301_n4244 (.O(FE_PHN4301_n4244), 
	.I(FE_PHN5546_n4244));
   BUFCKLHD FE_PHC4300_n4291 (.O(FE_PHN4300_n4291), 
	.I(FE_PHN5530_n4291));
   BUFLHD FE_PHC4299_n3046 (.O(FE_PHN4299_n3046), 
	.I(FE_PHN5498_n3046));
   BUFNHD FE_PHC4298_n3946 (.O(FE_PHN4298_n3946), 
	.I(FE_PHN5571_n3946));
   BUFCHD FE_PHC4297_n2967 (.O(FE_PHN4297_n2967), 
	.I(FE_PHN5005_n2967));
   BUFCHD FE_PHC4296_n4034 (.O(FE_PHN4296_n4034), 
	.I(FE_PHN6492_n4034));
   BUFCKMHD FE_PHC4295_n4103 (.O(FE_PHN4295_n4103), 
	.I(n4103));
   BUFCKLHD FE_PHC4294_n3030 (.O(FE_PHN4294_n3030), 
	.I(FE_PHN5560_n3030));
   BUFCHD FE_PHC4293_n4286 (.O(FE_PHN4293_n4286), 
	.I(FE_PHN5215_n4286));
   BUFCHD FE_PHC4292_n3983 (.O(FE_PHN4292_n3983), 
	.I(FE_PHN6466_n3983));
   BUFCKEHD FE_PHC4291_n951 (.O(FE_PHN4291_n951), 
	.I(FE_PHN3909_n951));
   BUFCKEHD FE_PHC4290_n1902 (.O(FE_PHN4290_n1902), 
	.I(FE_PHN5098_n1902));
   BUFCKEHD FE_PHC4289_n1069 (.O(FE_PHN4289_n1069), 
	.I(FE_PHN5114_n1069));
   BUFCKMHD FE_PHC4288_n1896 (.O(FE_PHN4288_n1896), 
	.I(FE_PHN5501_n1896));
   BUFCHD FE_PHC4287_n3087 (.O(FE_PHN4287_n3087), 
	.I(FE_PHN5301_n3087));
   BUFCHD FE_PHC4286_n1025 (.O(FE_PHN4286_n1025), 
	.I(FE_PHN5038_n1025));
   BUFCKEHD FE_PHC4285_n992 (.O(FE_PHN4285_n992), 
	.I(FE_PHN3647_n992));
   BUFCHD FE_PHC4284_n2968 (.O(FE_PHN4284_n2968), 
	.I(FE_PHN6486_n2968));
   BUFNHD FE_PHC4283_n934 (.O(FE_PHN4283_n934), 
	.I(FE_PHN3847_n934));
   BUFCHD FE_PHC4282_n1064 (.O(FE_PHN4282_n1064), 
	.I(FE_PHN5093_n1064));
   BUFCHD FE_PHC4281_n3929 (.O(FE_PHN4281_n3929), 
	.I(FE_PHN5116_n3929));
   BUFCKEHD FE_PHC4280_n2433 (.O(FE_PHN4280_n2433), 
	.I(FE_PHN5037_n2433));
   BUFCHD FE_PHC4279_n4408 (.O(FE_PHN4279_n4408), 
	.I(FE_PHN5316_n4408));
   BUFCKEHD FE_PHC4278_n4361 (.O(FE_PHN4278_n4361), 
	.I(FE_PHN5169_n4361));
   BUFCKEHD FE_PHC4277_n4362 (.O(FE_PHN4277_n4362), 
	.I(FE_PHN5021_n4362));
   BUFHHD FE_PHC4276_n3071 (.O(FE_PHN4276_n3071), 
	.I(FE_PHN5072_n3071));
   BUFCHD FE_PHC4275_n4260 (.O(FE_PHN4275_n4260), 
	.I(FE_PHN5146_n4260));
   BUFCKEHD FE_PHC4274_n2703 (.O(FE_PHN4274_n2703), 
	.I(n2703));
   BUFCKLHD FE_PHC4273_n4398 (.O(FE_PHN4273_n4398), 
	.I(FE_PHN5593_n4398));
   BUFCHD FE_PHC4272_n4220 (.O(FE_PHN4272_n4220), 
	.I(FE_PHN5260_n4220));
   BUFEHD FE_PHC4271_n1032 (.O(FE_PHN4271_n1032), 
	.I(FE_PHN5006_n1032));
   BUFCKMHD FE_PHC4270_n3132 (.O(FE_PHN4270_n3132), 
	.I(FE_PHN5641_n3132));
   BUFCKEHD FE_PHC4269_n2900 (.O(FE_PHN4269_n2900), 
	.I(FE_PHN5062_n2900));
   BUFCKMHD FE_PHC4268_n3117 (.O(FE_PHN4268_n3117), 
	.I(FE_PHN5639_n3117));
   BUFCHD FE_PHC4267_n846 (.O(FE_PHN4267_n846), 
	.I(FE_PHN6011_n846));
   BUFCHD FE_PHC4266_n887 (.O(FE_PHN4266_n887), 
	.I(FE_PHN5192_n887));
   BUFCKEHD FE_PHC4265_n2953 (.O(FE_PHN4265_n2953), 
	.I(FE_PHN4990_n2953));
   BUFCHD FE_PHC4264_n4307 (.O(FE_PHN4264_n4307), 
	.I(FE_PHN5008_n4307));
   BUFCKGHD FE_PHC4263_n4167 (.O(FE_PHN4263_n4167), 
	.I(FE_PHN5366_n4167));
   BUFCKIHD FE_PHC4262_n4023 (.O(FE_PHN4262_n4023), 
	.I(FE_PHN5359_n4023));
   BUFCKEHD FE_PHC4261_n852 (.O(FE_PHN4261_n852), 
	.I(FE_PHN5131_n852));
   BUFCHD FE_PHC4260_n3042 (.O(FE_PHN4260_n3042), 
	.I(FE_PHN5312_n3042));
   BUFCHD FE_PHC4259_n2985 (.O(FE_PHN4259_n2985), 
	.I(FE_PHN6449_n2985));
   BUFNHD FE_PHC4258_n3031 (.O(FE_PHN4258_n3031), 
	.I(FE_PHN5607_n3031));
   BUFCHD FE_PHC4257_ram_153__7_ (.O(FE_PHN4257_ram_153__7_), 
	.I(FE_PHN5221_ram_153__7_));
   BUFCHD FE_PHC4256_n4274 (.O(FE_PHN4256_n4274), 
	.I(FE_PHN6511_n4274));
   BUFCHD FE_PHC4255_n4010 (.O(FE_PHN4255_n4010), 
	.I(FE_PHN5065_n4010));
   BUFNHD FE_PHC4254_n3114 (.O(FE_PHN4254_n3114), 
	.I(FE_PHN5582_n3114));
   BUFCKEHD FE_PHC4253_n3966 (.O(FE_PHN4253_n3966), 
	.I(FE_PHN6461_n3966));
   BUFNHD FE_PHC4252_n3083 (.O(FE_PHN4252_n3083), 
	.I(FE_PHN5602_n3083));
   BUFCKEHD FE_PHC4251_n1873 (.O(FE_PHN4251_n1873), 
	.I(FE_PHN5073_n1873));
   BUFCKEHD FE_PHC4250_n1919 (.O(FE_PHN4250_n1919), 
	.I(FE_PHN6456_n1919));
   BUFCKEHD FE_PHC4249_n872 (.O(FE_PHN4249_n872), 
	.I(FE_PHN5034_n872));
   BUFCKGHD FE_PHC4248_n864 (.O(FE_PHN4248_n864), 
	.I(n864));
   BUFCKEHD FE_PHC4247_n2932 (.O(FE_PHN4247_n2932), 
	.I(FE_PHN3542_n2932));
   BUFCHD FE_PHC4246_n1886 (.O(FE_PHN4246_n1886), 
	.I(FE_PHN5079_n1886));
   BUFNHD FE_PHC4245_n2969 (.O(FE_PHN4245_n2969), 
	.I(FE_PHN5551_n2969));
   BUFCKMHD FE_PHC4244_n3095 (.O(FE_PHN4244_n3095), 
	.I(FE_PHN5624_n3095));
   BUFCKEHD FE_PHC4243_n3223 (.O(FE_PHN4243_n3223), 
	.I(FE_PHN5012_n3223));
   BUFCKEHD FE_PHC4242_n947 (.O(FE_PHN4242_n947), 
	.I(FE_PHN5057_n947));
   BUFCKEHD FE_PHC4241_n978 (.O(FE_PHN4241_n978), 
	.I(FE_PHN5134_n978));
   BUFCKMHD FE_PHC4240_n3911 (.O(FE_PHN4240_n3911), 
	.I(FE_PHN5610_n3911));
   BUFCHD FE_PHC4239_n1911 (.O(FE_PHN4239_n1911), 
	.I(FE_PHN5113_n1911));
   BUFHHD FE_PHC4238_n2980 (.O(FE_PHN4238_n2980), 
	.I(FE_PHN3518_n2980));
   BUFCKMHD FE_PHC4237_n4290 (.O(FE_PHN4237_n4290), 
	.I(FE_PHN5615_n4290));
   BUFCKEHD FE_PHC4236_n1904 (.O(FE_PHN4236_n1904), 
	.I(n1904));
   BUFJHD FE_PHC4235_n959 (.O(FE_PHN4235_n959), 
	.I(FE_PHN3827_n959));
   BUFNHD FE_PHC4234_n871 (.O(FE_PHN4234_n871), 
	.I(FE_PHN3684_n871));
   BUFCKEHD FE_PHC4233_n950 (.O(FE_PHN4233_n950), 
	.I(FE_PHN3670_n950));
   BUFCKEHD FE_PHC4232_n920 (.O(FE_PHN4232_n920), 
	.I(FE_PHN3876_n920));
   BUFLHD FE_PHC4231_n3110 (.O(FE_PHN4231_n3110), 
	.I(FE_PHN3772_n3110));
   BUFCKEHD FE_PHC4230_n1072 (.O(FE_PHN4230_n1072), 
	.I(FE_PHN5137_n1072));
   BUFCHD FE_PHC4229_n4327 (.O(FE_PHN4229_n4327), 
	.I(FE_PHN5139_n4327));
   BUFCKEHD FE_PHC4228_n945 (.O(FE_PHN4228_n945), 
	.I(FE_PHN5106_n945));
   BUFCKEHD FE_PHC4227_n3073 (.O(FE_PHN4227_n3073), 
	.I(FE_PHN4989_n3073));
   BUFCHD FE_PHC4226_n4363 (.O(FE_PHN4226_n4363), 
	.I(FE_PHN5178_n4363));
   BUFCKEHD FE_PHC4225_n989 (.O(FE_PHN4225_n989), 
	.I(n989));
   BUFCKLHD FE_PHC4224_ram_238__0_ (.O(FE_PHN4224_ram_238__0_), 
	.I(FE_PHN5552_ram_238__0_));
   BUFCKJHD FE_PHC4223_n3123 (.O(FE_PHN4223_n3123), 
	.I(FE_PHN5481_n3123));
   BUFCHD FE_PHC4222_n4110 (.O(FE_PHN4222_n4110), 
	.I(FE_PHN6442_n4110));
   BUFCHD FE_PHC4221_n848 (.O(FE_PHN4221_n848), 
	.I(FE_PHN5166_n848));
   BUFCKEHD FE_PHC4220_n4289 (.O(FE_PHN4220_n4289), 
	.I(FE_PHN5070_n4289));
   BUFHHD FE_PHC4219_n3987 (.O(FE_PHN4219_n3987), 
	.I(FE_PHN3238_n3987));
   BUFCKEHD FE_PHC4218_n1864 (.O(FE_PHN4218_n1864), 
	.I(FE_PHN5111_n1864));
   BUFCKEHD FE_PHC4217_n842 (.O(FE_PHN4217_n842), 
	.I(FE_PHN5135_n842));
   BUFCKEHD FE_PHC4216_n1087 (.O(FE_PHN4216_n1087), 
	.I(FE_PHN3658_n1087));
   BUFCKEHD FE_PHC4215_n2958 (.O(FE_PHN4215_n2958), 
	.I(FE_PHN5047_n2958));
   BUFCKEHD FE_PHC4214_n3007 (.O(FE_PHN4214_n3007), 
	.I(FE_PHN5184_n3007));
   BUFCHD FE_PHC4213_n4379 (.O(FE_PHN4213_n4379), 
	.I(FE_PHN5001_n4379));
   BUFCHD FE_PHC4212_n1077 (.O(FE_PHN4212_n1077), 
	.I(FE_PHN5149_n1077));
   BUFCKEHD FE_PHC4211_n2952 (.O(FE_PHN4211_n2952), 
	.I(FE_PHN5013_n2952));
   BUFCHD FE_PHC4210_n3138 (.O(FE_PHN4210_n3138), 
	.I(FE_PHN5279_n3138));
   BUFCKEHD FE_PHC4209_n2408 (.O(FE_PHN4209_n2408), 
	.I(FE_PHN4980_n2408));
   BUFCKEHD FE_PHC4208_n927 (.O(FE_PHN4208_n927), 
	.I(FE_PHN6455_n927));
   BUFCKEHD FE_PHC4207_n4000 (.O(FE_PHN4207_n4000), 
	.I(FE_PHN3650_n4000));
   BUFCHD FE_PHC4206_n3089 (.O(FE_PHN4206_n3089), 
	.I(FE_PHN5319_n3089));
   BUFCKEHD FE_PHC4205_n2415 (.O(FE_PHN4205_n2415), 
	.I(FE_PHN4987_n2415));
   BUFCKIHD FE_PHC4204_n3043 (.O(FE_PHN4204_n3043), 
	.I(n3043));
   BUFCHD FE_PHC4203_n4375 (.O(FE_PHN4203_n4375), 
	.I(FE_PHN5011_n4375));
   BUFCKJHD FE_PHC4202_n3070 (.O(FE_PHN4202_n3070), 
	.I(FE_PHN5406_n3070));
   BUFCKLHD FE_PHC4201_n4417 (.O(FE_PHN4201_n4417), 
	.I(FE_PHN5587_n4417));
   BUFCKEHD FE_PHC4200_n2982 (.O(FE_PHN4200_n2982), 
	.I(FE_PHN5136_n2982));
   BUFCKLHD FE_PHC4199_n4292 (.O(FE_PHN4199_n4292), 
	.I(FE_PHN5590_n4292));
   BUFCKEHD FE_PHC4198_n952 (.O(FE_PHN4198_n952), 
	.I(FE_PHN5053_n952));
   BUFLHD FE_PHC4197_n3972 (.O(FE_PHN4197_n3972), 
	.I(FE_PHN3526_n3972));
   BUFCKEHD FE_PHC4196_n3077 (.O(FE_PHN4196_n3077), 
	.I(FE_PHN5036_n3077));
   BUFCHD FE_PHC4195_n3012 (.O(FE_PHN4195_n3012), 
	.I(FE_PHN5190_n3012));
   BUFCKEHD FE_PHC4194_n893 (.O(FE_PHN4194_n893), 
	.I(FE_PHN5165_n893));
   BUFCHD FE_PHC4193_n1905 (.O(FE_PHN4193_n1905), 
	.I(FE_PHN5056_n1905));
   BUFCKEHD FE_PHC4192_n922 (.O(FE_PHN4192_n922), 
	.I(FE_PHN5088_n922));
   BUFCHD FE_PHC4191_n4001 (.O(FE_PHN4191_n4001), 
	.I(FE_PHN5026_n4001));
   BUFCKGHD FE_PHC4190_n4383 (.O(FE_PHN4190_n4383), 
	.I(FE_PHN5259_n4383));
   BUFCKMHD FE_PHC4189_n3111 (.O(FE_PHN4189_n3111), 
	.I(FE_PHN5622_n3111));
   BUFCHD FE_PHC4188_n4331 (.O(FE_PHN4188_n4331), 
	.I(FE_PHN6446_n4331));
   BUFCKEHD FE_PHC4187_n3027 (.O(FE_PHN4187_n3027), 
	.I(FE_PHN5161_n3027));
   BUFCKEHD FE_PHC4186_n1921 (.O(FE_PHN4186_n1921), 
	.I(FE_PHN4974_n1921));
   BUFCHD FE_PHC4185_ram_144__8_ (.O(FE_PHN4185_ram_144__8_), 
	.I(FE_PHN5046_ram_144__8_));
   BUFCKMHD FE_PHC4184_n3133 (.O(FE_PHN4184_n3133), 
	.I(FE_PHN5568_n3133));
   BUFCKEHD FE_PHC4183_n961 (.O(FE_PHN4183_n961), 
	.I(FE_PHN4979_n961));
   BUFCKEHD FE_PHC4182_n1040 (.O(FE_PHN4182_n1040), 
	.I(FE_PHN5089_n1040));
   BUFCHD FE_PHC4181_n4033 (.O(FE_PHN4181_n4033), 
	.I(FE_PHN5007_n4033));
   BUFMHD FE_PHC4180_n3959 (.O(FE_PHN4180_n3959), 
	.I(n3959));
   BUFCKEHD FE_PHC4179_n3217 (.O(FE_PHN4179_n3217), 
	.I(FE_PHN3905_n3217));
   BUFCKEHD FE_PHC4178_n4410 (.O(FE_PHN4178_n4410), 
	.I(FE_PHN5050_n4410));
   BUFLHD FE_PHC4177_n3078 (.O(FE_PHN4177_n3078), 
	.I(FE_PHN3481_n3078));
   BUFCKGHD FE_PHC4176_n4007 (.O(FE_PHN4176_n4007), 
	.I(FE_PHN5291_n4007));
   BUFCKMHD FE_PHC4175_n2999 (.O(FE_PHN4175_n2999), 
	.I(FE_PHN5569_n2999));
   BUFCKEHD FE_PHC4174_n3000 (.O(FE_PHN4174_n3000), 
	.I(FE_PHN6451_n3000));
   BUFCHD FE_PHC4173_n3026 (.O(FE_PHN4173_n3026), 
	.I(FE_PHN5231_n3026));
   BUFCKLHD FE_PHC4172_ram_237__7_ (.O(FE_PHN4172_ram_237__7_), 
	.I(FE_PHN5562_ram_237__7_));
   BUFNHD FE_PHC4171_n4269 (.O(FE_PHN4171_n4269), 
	.I(FE_PHN3687_n4269));
   BUFCHD FE_PHC4170_n3103 (.O(FE_PHN4170_n3103), 
	.I(FE_PHN5286_n3103));
   BUFCKEHD FE_PHC4169_n3978 (.O(FE_PHN4169_n3978), 
	.I(FE_PHN5027_n3978));
   BUFCHD FE_PHC4168_n943 (.O(FE_PHN4168_n943), 
	.I(FE_PHN5281_n943));
   BUFHHD FE_PHC4167_n3023 (.O(FE_PHN4167_n3023), 
	.I(FE_PHN3640_n3023));
   BUFCKEHD FE_PHC4166_n4111 (.O(FE_PHN4166_n4111), 
	.I(FE_PHN5060_n4111));
   BUFCKMHD FE_PHC4165_n884 (.O(FE_PHN4165_n884), 
	.I(FE_PHN5559_n884));
   BUFHHD FE_PHC4164_n946 (.O(FE_PHN4164_n946), 
	.I(FE_PHN3439_n946));
   BUFLHD FE_PHC4163_n4225 (.O(FE_PHN4163_n4225), 
	.I(FE_PHN3937_n4225));
   BUFCHD FE_PHC4162_n3056 (.O(FE_PHN4162_n3056), 
	.I(FE_PHN5080_n3056));
   BUFCHD FE_PHC4161_ram_145__0_ (.O(FE_PHN4161_ram_145__0_), 
	.I(FE_PHN5203_ram_145__0_));
   BUFCHD FE_PHC4160_n4028 (.O(FE_PHN4160_n4028), 
	.I(FE_PHN5157_n4028));
   BUFCKLHD FE_PHC4159_n4413 (.O(FE_PHN4159_n4413), 
	.I(FE_PHN5579_n4413));
   BUFCKMHD FE_PHC4158_n3003 (.O(FE_PHN4158_n3003), 
	.I(FE_PHN5520_n3003));
   BUFCHD FE_PHC4157_n4022 (.O(FE_PHN4157_n4022), 
	.I(FE_PHN4985_n4022));
   BUFCKLHD FE_PHC4156_n4254 (.O(FE_PHN4156_n4254), 
	.I(FE_PHN5574_n4254));
   BUFCKLHD FE_PHC4155_ram_229__3_ (.O(FE_PHN4155_ram_229__3_), 
	.I(FE_PHN5528_ram_229__3_));
   BUFCHD FE_PHC4154_n901 (.O(FE_PHN4154_n901), 
	.I(FE_PHN6472_n901));
   BUFMHD FE_PHC4153_n4239 (.O(FE_PHN4153_n4239), 
	.I(FE_PHN3624_n4239));
   BUFCHD FE_PHC4152_n1088 (.O(FE_PHN4152_n1088), 
	.I(FE_PHN5045_n1088));
   BUFCHD FE_PHC4151_n3053 (.O(FE_PHN4151_n3053), 
	.I(FE_PHN5162_n3053));
   BUFCHD FE_PHC4150_n930 (.O(FE_PHN4150_n930), 
	.I(FE_PHN6441_n930));
   BUFCHD FE_PHC4149_n4031 (.O(FE_PHN4149_n4031), 
	.I(FE_PHN6439_n4031));
   BUFEHD FE_PHC4148_n1078 (.O(FE_PHN4148_n1078), 
	.I(FE_PHN3476_n1078));
   BUFCKEHD FE_PHC4147_n928 (.O(FE_PHN4147_n928), 
	.I(FE_PHN4978_n928));
   BUFCHD FE_PHC4146_n3979 (.O(FE_PHN4146_n3979), 
	.I(FE_PHN6459_n3979));
   BUFHHD FE_PHC4145_n4214 (.O(FE_PHN4145_n4214), 
	.I(n4214));
   BUFCHD FE_PHC4144_n919 (.O(FE_PHN4144_n919), 
	.I(FE_PHN5054_n919));
   BUFLHD FE_PHC4143_n3943 (.O(FE_PHN4143_n3943), 
	.I(FE_PHN3963_n3943));
   BUFCHD FE_PHC4142_n4380 (.O(FE_PHN4142_n4380), 
	.I(FE_PHN5219_n4380));
   BUFCKMHD FE_PHC4141_n3115 (.O(FE_PHN4141_n3115), 
	.I(FE_PHN5588_n3115));
   BUFHHD FE_PHC4140_n4014 (.O(FE_PHN4140_n4014), 
	.I(FE_PHN3284_n4014));
   BUFCKEHD FE_PHC4139_n4009 (.O(FE_PHN4139_n4009), 
	.I(FE_PHN4964_n4009));
   BUFCKEHD FE_PHC4138_n2389 (.O(FE_PHN4138_n2389), 
	.I(FE_PHN5015_n2389));
   BUFCHD FE_PHC4137_n3982 (.O(FE_PHN4137_n3982), 
	.I(FE_PHN5132_n3982));
   BUFNHD FE_PHC4136_n4245 (.O(FE_PHN4136_n4245), 
	.I(FE_PHN3627_n4245));
   BUFCKEHD FE_PHC4135_n3265 (.O(FE_PHN4135_n3265), 
	.I(FE_PHN3688_n3265));
   BUFCKMHD FE_PHC4134_ram_145__1_ (.O(FE_PHN4134_ram_145__1_), 
	.I(FE_PHN3502_ram_145__1_));
   BUFCHD FE_PHC4133_n4008 (.O(FE_PHN4133_n4008), 
	.I(FE_PHN6454_n4008));
   BUFCKEHD FE_PHC4132_n4279 (.O(FE_PHN4132_n4279), 
	.I(FE_PHN5123_n4279));
   BUFCHD FE_PHC4131_n1008 (.O(FE_PHN4131_n1008), 
	.I(FE_PHN5018_n1008));
   BUFCKEHD FE_PHC4130_n1056 (.O(FE_PHN4130_n1056), 
	.I(FE_PHN5031_n1056));
   BUFCKMHD FE_PHC4129_ram_229__12_ (.O(FE_PHN4129_ram_229__12_), 
	.I(FE_PHN5526_ram_229__12_));
   BUFCHD FE_PHC4128_n865 (.O(FE_PHN4128_n865), 
	.I(FE_PHN5151_n865));
   BUFNHD FE_PHC4127_n3019 (.O(FE_PHN4127_n3019), 
	.I(FE_PHN5538_n3019));
   BUFCKEHD FE_PHC4126_n3009 (.O(FE_PHN4126_n3009), 
	.I(FE_PHN5115_n3009));
   BUFCKEHD FE_PHC4125_n4421 (.O(FE_PHN4125_n4421), 
	.I(FE_PHN3385_n4421));
   BUFCKIHD FE_PHC4124_n866 (.O(FE_PHN4124_n866), 
	.I(n866));
   BUFCKLHD FE_PHC4123_ram_145__7_ (.O(FE_PHN4123_ram_145__7_), 
	.I(FE_PHN3593_ram_145__7_));
   BUFCHD FE_PHC4122_n4196 (.O(FE_PHN4122_n4196), 
	.I(FE_PHN5285_n4196));
   BUFCKEHD FE_PHC4121_n857 (.O(FE_PHN4121_n857), 
	.I(FE_PHN5043_n857));
   BUFCKMHD FE_PHC4120_n3081 (.O(FE_PHN4120_n3081), 
	.I(FE_PHN5578_n3081));
   BUFCKLHD FE_PHC4119_n4295 (.O(FE_PHN4119_n4295), 
	.I(FE_PHN5504_n4295));
   BUFCHD FE_PHC4118_n925 (.O(FE_PHN4118_n925), 
	.I(FE_PHN5148_n925));
   BUFCHD FE_PHC4117_n2374 (.O(FE_PHN4117_n2374), 
	.I(FE_PHN5975_n2374));
   BUFCKLHD FE_PHC4116_n4238 (.O(FE_PHN4116_n4238), 
	.I(FE_PHN5479_n4238));
   BUFCKEHD FE_PHC4115_n4146 (.O(FE_PHN4115_n4146), 
	.I(FE_PHN3413_n4146));
   BUFCKLHD FE_PHC4114_n4340 (.O(FE_PHN4114_n4340), 
	.I(n4340));
   BUFCKEHD FE_PHC4113_n3915 (.O(FE_PHN4113_n3915), 
	.I(n3915));
   BUFCKIHD FE_PHC4112_n2400 (.O(FE_PHN4112_n2400), 
	.I(n2400));
   BUFCKEHD FE_PHC4111_n4387 (.O(FE_PHN4111_n4387), 
	.I(FE_PHN5010_n4387));
   BUFCKJHD FE_PHC4110_n3134 (.O(FE_PHN4110_n3134), 
	.I(FE_PHN5428_n3134));
   BUFCKNHD FE_PHC4109_n4138 (.O(FE_PHN4109_n4138), 
	.I(FE_PHN5595_n4138));
   BUFNHD FE_PHC4108_n3099 (.O(FE_PHN4108_n3099), 
	.I(FE_PHN3328_n3099));
   BUFCKEHD FE_PHC4107_n2994 (.O(FE_PHN4107_n2994), 
	.I(FE_PHN4998_n2994));
   BUFCHD FE_PHC4106_n3010 (.O(FE_PHN4106_n3010), 
	.I(FE_PHN5024_n3010));
   BUFCKMHD FE_PHC4105_ram_221__1_ (.O(FE_PHN4105_ram_221__1_), 
	.I(FE_PHN3488_ram_221__1_));
   BUFCHD FE_PHC4104_n958 (.O(FE_PHN4104_n958), 
	.I(FE_PHN4982_n958));
   BUFCKJHD FE_PHC4103_n876 (.O(FE_PHN4103_n876), 
	.I(FE_PHN3931_n876));
   BUFCKEHD FE_PHC4102_n2961 (.O(FE_PHN4102_n2961), 
	.I(FE_PHN4972_n2961));
   BUFLHD FE_PHC4101_n3102 (.O(FE_PHN4101_n3102), 
	.I(FE_PHN3590_n3102));
   BUFCHD FE_PHC4100_n4006 (.O(FE_PHN4100_n4006), 
	.I(FE_PHN5075_n4006));
   BUFCKEHD FE_PHC4099_n4371 (.O(FE_PHN4099_n4371), 
	.I(FE_PHN4995_n4371));
   BUFNHD FE_PHC4098_n3084 (.O(FE_PHN4098_n3084), 
	.I(FE_PHN3739_n3084));
   BUFCKEHD FE_PHC4097_n2991 (.O(FE_PHN4097_n2991), 
	.I(FE_PHN5197_n2991));
   BUFCKJHD FE_PHC4096_n3124 (.O(FE_PHN4096_n3124), 
	.I(FE_PHN5412_n3124));
   BUFCKEHD FE_PHC4095_n4356 (.O(FE_PHN4095_n4356), 
	.I(FE_PHN5049_n4356));
   BUFCHD FE_PHC4094_n4263 (.O(FE_PHN4094_n4263), 
	.I(FE_PHN5082_n4263));
   BUFCHD FE_PHC4093_n4389 (.O(FE_PHN4093_n4389), 
	.I(FE_PHN4981_n4389));
   BUFCKLHD FE_PHC4092_ram_17__14_ (.O(FE_PHN4092_ram_17__14_), 
	.I(FE_PHN5480_ram_17__14_));
   BUFNHD FE_PHC4091_n4367 (.O(FE_PHN4091_n4367), 
	.I(FE_PHN5512_n4367));
   BUFCKEHD FE_PHC4090_n2955 (.O(FE_PHN4090_n2955), 
	.I(FE_PHN5052_n2955));
   BUFCHD FE_PHC4089_n3948 (.O(FE_PHN4089_n3948), 
	.I(FE_PHN5126_n3948));
   BUFNHD FE_PHC4088_n3127 (.O(FE_PHN4088_n3127), 
	.I(FE_PHN3438_n3127));
   BUFCKEHD FE_PHC4087_ram_98__3_ (.O(FE_PHN4087_ram_98__3_), 
	.I(FE_PHN3347_ram_98__3_));
   BUFCKEHD FE_PHC4086_n4142 (.O(FE_PHN4086_n4142), 
	.I(FE_PHN6443_n4142));
   BUFCKJHD FE_PHC4085_n3048 (.O(FE_PHN4085_n3048), 
	.I(n3048));
   BUFCKEHD FE_PHC4084_n2956 (.O(FE_PHN4084_n2956), 
	.I(FE_PHN5067_n2956));
   BUFCHD FE_PHC4083_n855 (.O(FE_PHN4083_n855), 
	.I(FE_PHN5066_n855));
   BUFCKEHD FE_PHC4082_n914 (.O(FE_PHN4082_n914), 
	.I(FE_PHN6440_n914));
   BUFCKMHD FE_PHC4081_n2973 (.O(FE_PHN4081_n2973), 
	.I(FE_PHN5516_n2973));
   BUFCHD FE_PHC4080_n3105 (.O(FE_PHN4080_n3105), 
	.I(FE_PHN5300_n3105));
   BUFCHD FE_PHC4079_n3092 (.O(FE_PHN4079_n3092), 
	.I(FE_PHN5104_n3092));
   BUFCHD FE_PHC4078_n3104 (.O(FE_PHN4078_n3104), 
	.I(FE_PHN5193_n3104));
   BUFCHD FE_PHC4077_n3107 (.O(FE_PHN4077_n3107), 
	.I(FE_PHN5091_n3107));
   BUFCKLHD FE_PHC4076_n4406 (.O(FE_PHN4076_n4406), 
	.I(FE_PHN5518_n4406));
   BUFCKEHD FE_PHC4075_n2962 (.O(FE_PHN4075_n2962), 
	.I(FE_PHN3810_n2962));
   BUFCKEHD FE_PHC4074_n4359 (.O(FE_PHN4074_n4359), 
	.I(FE_PHN5048_n4359));
   BUFCKLHD FE_PHC4073_n1005 (.O(FE_PHN4073_n1005), 
	.I(FE_PHN3340_n1005));
   BUFCKMHD FE_PHC4072_n3939 (.O(FE_PHN4072_n3939), 
	.I(FE_PHN5557_n3939));
   BUFCKMHD FE_PHC4071_n4003 (.O(FE_PHN4071_n4003), 
	.I(FE_PHN5533_n4003));
   BUFCKEHD FE_PHC4070_n4323 (.O(FE_PHN4070_n4323), 
	.I(FE_PHN4961_n4323));
   BUFCKEHD FE_PHC4069_n3260 (.O(FE_PHN4069_n3260), 
	.I(FE_PHN6484_n3260));
   BUFCKJHD FE_PHC4068_n3108 (.O(FE_PHN4068_n3108), 
	.I(FE_PHN5423_n3108));
   BUFEHD FE_PHC4067_n1045 (.O(FE_PHN4067_n1045), 
	.I(FE_PHN5004_n1045));
   BUFNHD FE_PHC4066_n4339 (.O(FE_PHN4066_n4339), 
	.I(n4339));
   BUFCKEHD FE_PHC4065_n3128 (.O(FE_PHN4065_n3128), 
	.I(FE_PHN5017_n3128));
   BUFCKEHD FE_PHC4064_n4005 (.O(FE_PHN4064_n4005), 
	.I(FE_PHN4996_n4005));
   BUFCKEHD FE_PHC4063_n2979 (.O(FE_PHN4063_n2979), 
	.I(FE_PHN4983_n2979));
   BUFCKEHD FE_PHC4062_n2431 (.O(FE_PHN4062_n2431), 
	.I(FE_PHN5023_n2431));
   BUFCKJHD FE_PHC4061_n3118 (.O(FE_PHN4061_n3118), 
	.I(FE_PHN5387_n3118));
   BUFLHD FE_PHC4060_n4251 (.O(FE_PHN4060_n4251), 
	.I(FE_PHN3357_n4251));
   BUFCKMHD FE_PHC4059_n3001 (.O(FE_PHN4059_n3001), 
	.I(FE_PHN3338_n3001));
   BUFCKLHD FE_PHC4058_n2178 (.O(FE_PHN4058_n2178), 
	.I(n2178));
   BUFCKEHD FE_PHC4057_n2977 (.O(FE_PHN4057_n2977), 
	.I(FE_PHN4999_n2977));
   BUFCKLHD FE_PHC4056_n4388 (.O(FE_PHN4056_n4388), 
	.I(FE_PHN3267_n4388));
   BUFCHD FE_PHC4055_n4405 (.O(FE_PHN4055_n4405), 
	.I(FE_PHN5086_n4405));
   BUFCHD FE_PHC4054_n984 (.O(FE_PHN4054_n984), 
	.I(FE_PHN5000_n984));
   BUFHHD FE_PHC4053_n1093 (.O(FE_PHN4053_n1093), 
	.I(FE_PHN3408_n1093));
   BUFNHD FE_PHC4052_n3116 (.O(FE_PHN4052_n3116), 
	.I(FE_PHN3372_n3116));
   BUFCHD FE_PHC4051_n1048 (.O(FE_PHN4051_n1048), 
	.I(FE_PHN4965_n1048));
   BUFCKEHD FE_PHC4050_n2981 (.O(FE_PHN4050_n2981), 
	.I(FE_PHN4994_n2981));
   BUFCKJHD FE_PHC4049_n3022 (.O(FE_PHN4049_n3022), 
	.I(FE_PHN5376_n3022));
   BUFCKEHD FE_PHC4048_n4372 (.O(FE_PHN4048_n4372), 
	.I(FE_PHN5030_n4372));
   BUFCKEHD FE_PHC4047_n2978 (.O(FE_PHN4047_n2978), 
	.I(FE_PHN4986_n2978));
   BUFCKEHD FE_PHC4046_n960 (.O(FE_PHN4046_n960), 
	.I(FE_PHN4976_n960));
   BUFLHD FE_PHC4045_n3112 (.O(FE_PHN4045_n3112), 
	.I(FE_PHN3629_n3112));
   BUFCHD FE_PHC4044_n3999 (.O(FE_PHN4044_n3999), 
	.I(FE_PHN4967_n3999));
   BUFCHD FE_PHC4043_n3930 (.O(FE_PHN4043_n3930), 
	.I(FE_PHN5039_n3930));
   BUFNHD FE_PHC4042_n3035 (.O(FE_PHN4042_n3035), 
	.I(FE_PHN3337_n3035));
   BUFCKMHD FE_PHC4041_n3100 (.O(FE_PHN4041_n3100), 
	.I(FE_PHN3264_n3100));
   BUFCHD FE_PHC4040_n4385 (.O(FE_PHN4040_n4385), 
	.I(FE_PHN5061_n4385));
   BUFCKMHD FE_PHC4039_n4384 (.O(FE_PHN4039_n4384), 
	.I(FE_PHN5547_n4384));
   BUFNHD FE_PHC4038_n856 (.O(FE_PHN4038_n856), 
	.I(FE_PHN3345_n856));
   BUFCKEHD FE_PHC4037_n1090 (.O(FE_PHN4037_n1090), 
	.I(FE_PHN3368_n1090));
   BUFNHD FE_PHC4036_n3914 (.O(FE_PHN4036_n3914), 
	.I(FE_PHN3601_n3914));
   BUFCKLHD FE_PHC4035_n4230 (.O(FE_PHN4035_n4230), 
	.I(FE_PHN3321_n4230));
   BUFCKEHD FE_PHC4034_n3937 (.O(FE_PHN4034_n3937), 
	.I(FE_PHN5097_n3937));
   BUFCKMHD FE_PHC4033_n918 (.O(FE_PHN4033_n918), 
	.I(FE_PHN3363_n918));
   BUFHHD FE_PHC4032_n4204 (.O(FE_PHN4032_n4204), 
	.I(FE_PHN3675_n4204));
   BUFCKEHD FE_PHC4031_n3947 (.O(FE_PHN4031_n3947), 
	.I(FE_PHN3346_n3947));
   BUFCHD FE_PHC4030_n2976 (.O(FE_PHN4030_n2976), 
	.I(FE_PHN5096_n2976));
   BUFNHD FE_PHC4029_n3032 (.O(FE_PHN4029_n3032), 
	.I(FE_PHN3411_n3032));
   BUFNHD FE_PHC4028_n3922 (.O(FE_PHN4028_n3922), 
	.I(FE_PHN3356_n3922));
   BUFCKEHD FE_PHC4027_n970 (.O(FE_PHN4027_n970), 
	.I(FE_PHN4966_n970));
   BUFCHD FE_PHC4026_ram_145__10_ (.O(FE_PHN4026_ram_145__10_), 
	.I(FE_PHN5074_ram_145__10_));
   BUFCHD FE_PHC4025_n3931 (.O(FE_PHN4025_n3931), 
	.I(FE_PHN4973_n3931));
   BUFCHD FE_PHC4024_n4324 (.O(FE_PHN4024_n4324), 
	.I(FE_PHN5032_n4324));
   BUFHHD FE_PHC4023_n4343 (.O(FE_PHN4023_n4343), 
	.I(FE_PHN3261_n4343));
   BUFCHD FE_PHC4022_n899 (.O(FE_PHN4022_n899), 
	.I(FE_PHN6110_n899));
   BUFCKEHD FE_PHC4021_n4399 (.O(FE_PHN4021_n4399), 
	.I(FE_PHN5014_n4399));
   BUFNHD FE_PHC4020_n3096 (.O(FE_PHN4020_n3096), 
	.I(FE_PHN3461_n3096));
   BUFCHD FE_PHC4019_n2966 (.O(FE_PHN4019_n2966), 
	.I(FE_PHN4984_n2966));
   BUFCKLHD FE_PHC4018_n3094 (.O(FE_PHN4018_n3094), 
	.I(FE_PHN5448_n3094));
   BUFCHD FE_PHC4017_n3926 (.O(FE_PHN4017_n3926), 
	.I(FE_PHN5107_n3926));
   BUFNHD FE_PHC4016_n3954 (.O(FE_PHN4016_n3954), 
	.I(FE_PHN3278_n3954));
   BUFLHD FE_PHC4015_n3993 (.O(FE_PHN4015_n3993), 
	.I(FE_PHN3273_n3993));
   BUFCKGHD FE_PHC4014_n4377 (.O(FE_PHN4014_n4377), 
	.I(FE_PHN5211_n4377));
   BUFCKGHD FE_PHC4013_n3998 (.O(FE_PHN4013_n3998), 
	.I(FE_PHN3274_n3998));
   BUFCKLHD FE_PHC4012_n4195 (.O(FE_PHN4012_n4195), 
	.I(FE_PHN5470_n4195));
   BUFCHD FE_PHC4011_n3125 (.O(FE_PHN4011_n3125), 
	.I(FE_PHN5305_n3125));
   BUFCHD FE_PHC4009_n2297 (.O(FE_PHN4009_n2297), 
	.I(n2297));
   BUFCHD FE_PHC4008_n889 (.O(FE_PHN4008_n889), 
	.I(FE_PHN5427_n889));
   BUFHHD FE_PHC4007_n4416 (.O(FE_PHN4007_n4416), 
	.I(n4416));
   BUFEHD FE_PHC4006_n961 (.O(FE_PHN4006_n961), 
	.I(n961));
   BUFEHD FE_PHC4005_n898 (.O(FE_PHN4005_n898), 
	.I(n898));
   BUFEHD FE_PHC4004_n3034 (.O(FE_PHN4004_n3034), 
	.I(n3034));
   BUFCHD FE_PHC4003_n4032 (.O(FE_PHN4003_n4032), 
	.I(n4032));
   BUFCHD FE_PHC4002_n1143 (.O(FE_PHN4002_n1143), 
	.I(n1143));
   BUFEHD FE_PHC4001_n3004 (.O(FE_PHN4001_n3004), 
	.I(n3004));
   BUFEHD FE_PHC4000_n4370 (.O(FE_PHN4000_n4370), 
	.I(n4370));
   BUFCHD FE_PHC3999_n1042 (.O(FE_PHN3999_n1042), 
	.I(n1042));
   BUFCHD FE_PHC3998_n896 (.O(FE_PHN3998_n896), 
	.I(n896));
   BUFKHD FE_PHC3997_n892 (.O(FE_PHN3997_n892), 
	.I(n892));
   BUFCHD FE_PHC3996_n2944 (.O(FE_PHN3996_n2944), 
	.I(FE_PHN5472_n2944));
   BUFLHD FE_PHC3995_n3135 (.O(FE_PHN3995_n3135), 
	.I(n3135));
   BUFEHD FE_PHC3994_n4407 (.O(FE_PHN3994_n4407), 
	.I(n4407));
   BUFEHD FE_PHC3993_n2954 (.O(FE_PHN3993_n2954), 
	.I(n2954));
   BUFEHD FE_PHC3992_n2388 (.O(FE_PHN3992_n2388), 
	.I(n2388));
   BUFHHD FE_PHC3991_n3130 (.O(FE_PHN3991_n3130), 
	.I(n3130));
   BUFHHD FE_PHC3990_n870 (.O(FE_PHN3990_n870), 
	.I(n870));
   BUFEHD FE_PHC3989_n976 (.O(FE_PHN3989_n976), 
	.I(n976));
   BUFLHD FE_PHC3988_n4202 (.O(FE_PHN3988_n4202), 
	.I(n4202));
   BUFEHD FE_PHC3987_n2963 (.O(FE_PHN3987_n2963), 
	.I(n2963));
   BUFEHD FE_PHC3986_n3977 (.O(FE_PHN3986_n3977), 
	.I(n3977));
   BUFHHD FE_PHC3985_n3257 (.O(FE_PHN3985_n3257), 
	.I(n3257));
   BUFEHD FE_PHC3984_n1000 (.O(FE_PHN3984_n1000), 
	.I(n1000));
   BUFCHD FE_PHC3983_n2722 (.O(FE_PHN3983_n2722), 
	.I(n2722));
   BUFCKMHD FE_PHC3982_n3920 (.O(FE_PHN3982_n3920), 
	.I(n3920));
   BUFCKEHD FE_PHC3981_n4403 (.O(FE_PHN3981_n4403), 
	.I(n4403));
   BUFEHD FE_PHC3980_n2952 (.O(FE_PHN3980_n2952), 
	.I(n2952));
   BUFCKEHD FE_PHC3979_n2933 (.O(FE_PHN3979_n2933), 
	.I(n2933));
   BUFCHD FE_PHC3978_n2959 (.O(FE_PHN3978_n2959), 
	.I(n2959));
   BUFCHD FE_PHC3977_n846 (.O(FE_PHN3977_n846), 
	.I(n846));
   BUFEHD FE_PHC3976_n944 (.O(FE_PHN3976_n944), 
	.I(n944));
   BUFEHD FE_PHC3975_n4289 (.O(FE_PHN3975_n4289), 
	.I(n4289));
   BUFCHD FE_PHC3974_n1911 (.O(FE_PHN3974_n1911), 
	.I(n1911));
   BUFEHD FE_PHC3973_n3114 (.O(FE_PHN3973_n3114), 
	.I(n3114));
   BUFCKNHD FE_PHC3972_n2258 (.O(FE_PHN3972_n2258), 
	.I(FE_PHN4765_n2258));
   BUFEHD FE_PHC3971_n891 (.O(FE_PHN3971_n891), 
	.I(n891));
   BUFEHD FE_PHC3970_n4361 (.O(FE_PHN3970_n4361), 
	.I(n4361));
   BUFHHD FE_PHC3969_n2623 (.O(FE_PHN3969_n2623), 
	.I(n2623));
   BUFIHD FE_PHC3968_n3255 (.O(FE_PHN3968_n3255), 
	.I(n3255));
   BUFEHD FE_PHC3967_n3066 (.O(FE_PHN3967_n3066), 
	.I(n3066));
   BUFCKEHD FE_PHC3966_n3962 (.O(FE_PHN3966_n3962), 
	.I(n3962));
   BUFEHD FE_PHC3965_n4248 (.O(FE_PHN3965_n4248), 
	.I(n4248));
   BUFHHD FE_PHC3964_n4401 (.O(FE_PHN3964_n4401), 
	.I(n4401));
   BUFCHD FE_PHC3963_n3943 (.O(FE_PHN3963_n3943), 
	.I(n3943));
   BUFEHD FE_PHC3962_n2621 (.O(FE_PHN3962_n2621), 
	.I(n2621));
   BUFIHD FE_PHC3961_n4276 (.O(FE_PHN3961_n4276), 
	.I(n4276));
   BUFCHD FE_PHC3960_n885 (.O(FE_PHN3960_n885), 
	.I(n885));
   BUFEHD FE_PHC3959_n3076 (.O(FE_PHN3959_n3076), 
	.I(n3076));
   BUFEHD FE_PHC3958_n3122 (.O(FE_PHN3958_n3122), 
	.I(n3122));
   BUFCHD FE_PHC3957_n969 (.O(FE_PHN3957_n969), 
	.I(n969));
   BUFCHD FE_PHC3956_n966 (.O(FE_PHN3956_n966), 
	.I(FE_PHN5431_n966));
   BUFCKNHD FE_PHC3955_n2605 (.O(FE_PHN3955_n2605), 
	.I(n2605));
   BUFEHD FE_PHC3954_n3080 (.O(FE_PHN3954_n3080), 
	.I(n3080));
   BUFCKEHD FE_PHC3953_n4268 (.O(FE_PHN3953_n4268), 
	.I(n4268));
   BUFEHD FE_PHC3952_n4036 (.O(FE_PHN3952_n4036), 
	.I(n4036));
   BUFEHD FE_PHC3951_n2946 (.O(FE_PHN3951_n2946), 
	.I(n2946));
   BUFNHD FE_PHC3950_n4097 (.O(FE_PHN3950_n4097), 
	.I(n4097));
   BUFJHD FE_PHC3949_n2564 (.O(FE_PHN3949_n2564), 
	.I(n2564));
   BUFCHD FE_PHC3948_n4168 (.O(FE_PHN3948_n4168), 
	.I(FE_PHN5584_n4168));
   BUFCHD FE_PHC3947_n4273 (.O(FE_PHN3947_n4273), 
	.I(n4273));
   BUFCHD FE_PHC3946_n3141 (.O(FE_PHN3946_n3141), 
	.I(n3141));
   BUFMHD FE_PHC3945_n4420 (.O(FE_PHN3945_n4420), 
	.I(n4420));
   BUFEHD FE_PHC3944_n3960 (.O(FE_PHN3944_n3960), 
	.I(n3960));
   BUFEHD FE_PHC3943_n4387 (.O(FE_PHN3943_n4387), 
	.I(n4387));
   BUFCHD FE_PHC3942_n3139 (.O(FE_PHN3942_n3139), 
	.I(n3139));
   BUFCKEHD FE_PHC3941_n3953 (.O(FE_PHN3941_n3953), 
	.I(n3953));
   BUFEHD FE_PHC3940_n968 (.O(FE_PHN3940_n968), 
	.I(n968));
   BUFCKEHD FE_PHC3939_n2385 (.O(FE_PHN3939_n2385), 
	.I(n2385));
   BUFCHD FE_PHC3938_n1110 (.O(FE_PHN3938_n1110), 
	.I(n1110));
   BUFEHD FE_PHC3937_n4225 (.O(FE_PHN3937_n4225), 
	.I(n4225));
   BUFEHD FE_PHC3936_n4333 (.O(FE_PHN3936_n4333), 
	.I(n4333));
   BUFEHD FE_PHC3935_n1034 (.O(FE_PHN3935_n1034), 
	.I(n1034));
   BUFCKEHD FE_PHC3934_n4185 (.O(FE_PHN3934_n4185), 
	.I(n4185));
   BUFCHD FE_PHC3933_n4241 (.O(FE_PHN3933_n4241), 
	.I(n4241));
   BUFEHD FE_PHC3932_n3050 (.O(FE_PHN3932_n3050), 
	.I(n3050));
   BUFEHD FE_PHC3931_n876 (.O(FE_PHN3931_n876), 
	.I(n876));
   BUFCHD FE_PHC3930_n4210 (.O(FE_PHN3930_n4210), 
	.I(FE_PHN4680_n4210));
   BUFHHD FE_PHC3929_n2945 (.O(FE_PHN3929_n2945), 
	.I(n2945));
   BUFCHD FE_PHC3928_n3975 (.O(FE_PHN3928_n3975), 
	.I(n3975));
   BUFJHD FE_PHC3927_n4046 (.O(FE_PHN3927_n4046), 
	.I(n4046));
   BUFJHD FE_PHC3926_n886 (.O(FE_PHN3926_n886), 
	.I(n886));
   BUFEHD FE_PHC3925_n4259 (.O(FE_PHN3925_n4259), 
	.I(n4259));
   BUFCHD FE_PHC3924_ram_20__10_ (.O(FE_PHN3924_ram_20__10_), 
	.I(\ram[20][10] ));
   BUFCHD FE_PHC3923_n4368 (.O(FE_PHN3923_n4368), 
	.I(n4368));
   BUFCHD FE_PHC3922_n988 (.O(FE_PHN3922_n988), 
	.I(n988));
   BUFEHD FE_PHC3921_n2419 (.O(FE_PHN3921_n2419), 
	.I(n2419));
   BUFKHD FE_PHC3920_n2580 (.O(FE_PHN3920_n2580), 
	.I(n2580));
   BUFCHD FE_PHC3919_n936 (.O(FE_PHN3919_n936), 
	.I(n936));
   BUFCHD FE_PHC3918_n4187 (.O(FE_PHN3918_n4187), 
	.I(FE_PHN5563_n4187));
   BUFCHD FE_PHC3917_n2554 (.O(FE_PHN3917_n2554), 
	.I(n2554));
   BUFCKEHD FE_PHC3916_n3219 (.O(FE_PHN3916_n3219), 
	.I(n3219));
   BUFCKEHD FE_PHC3915_n4215 (.O(FE_PHN3915_n4215), 
	.I(FE_PHN4704_n4215));
   BUFEHD FE_PHC3914_n4410 (.O(FE_PHN3914_n4410), 
	.I(n4410));
   BUFNHD FE_PHC3913_n4094 (.O(FE_PHN3913_n4094), 
	.I(n4094));
   BUFEHD FE_PHC3912_n4373 (.O(FE_PHN3912_n4373), 
	.I(n4373));
   BUFEHD FE_PHC3911_n3085 (.O(FE_PHN3911_n3085), 
	.I(n3085));
   BUFEHD FE_PHC3910_n4242 (.O(FE_PHN3910_n4242), 
	.I(n4242));
   BUFEHD FE_PHC3909_n951 (.O(FE_PHN3909_n951), 
	.I(n951));
   BUFEHD FE_PHC3908_n3207 (.O(FE_PHN3908_n3207), 
	.I(n3207));
   BUFHHD FE_PHC3907_n986 (.O(FE_PHN3907_n986), 
	.I(n986));
   BUFCHD FE_PHC3906_n3067 (.O(FE_PHN3906_n3067), 
	.I(FE_PHN5323_n3067));
   BUFCHD FE_PHC3905_n3217 (.O(FE_PHN3905_n3217), 
	.I(n3217));
   BUFHHD FE_PHC3904_n2965 (.O(FE_PHN3904_n2965), 
	.I(n2965));
   BUFCKEHD FE_PHC3903_n851 (.O(FE_PHN3903_n851), 
	.I(n851));
   BUFCKEHD FE_PHC3902_n4217 (.O(FE_PHN3902_n4217), 
	.I(n4217));
   BUFEHD FE_PHC3901_n3011 (.O(FE_PHN3901_n3011), 
	.I(n3011));
   BUFEHD FE_PHC3900_n2735 (.O(FE_PHN3900_n2735), 
	.I(n2735));
   BUFEHD FE_PHC3899_n954 (.O(FE_PHN3899_n954), 
	.I(n954));
   BUFCHD FE_PHC3898_n4183 (.O(FE_PHN3898_n4183), 
	.I(n4183));
   BUFEHD FE_PHC3897_n3036 (.O(FE_PHN3897_n3036), 
	.I(n3036));
   BUFEHD FE_PHC3896_n4338 (.O(FE_PHN3896_n4338), 
	.I(n4338));
   BUFEHD FE_PHC3895_n2993 (.O(FE_PHN3895_n2993), 
	.I(n2993));
   BUFCHD FE_PHC3894_n900 (.O(FE_PHN3894_n900), 
	.I(n900));
   BUFEHD FE_PHC3893_n1918 (.O(FE_PHN3893_n1918), 
	.I(n1918));
   BUFEHD FE_PHC3892_n945 (.O(FE_PHN3892_n945), 
	.I(n945));
   BUFCKEHD FE_PHC3891_n3025 (.O(FE_PHN3891_n3025), 
	.I(n3025));
   BUFIHD FE_PHC3890_n850 (.O(FE_PHN3890_n850), 
	.I(n850));
   BUFCHD FE_PHC3889_n3079 (.O(FE_PHN3889_n3079), 
	.I(FE_PHN5140_n3079));
   BUFEHD FE_PHC3888_n3082 (.O(FE_PHN3888_n3082), 
	.I(n3082));
   BUFCHD FE_PHC3887_n2383 (.O(FE_PHN3887_n2383), 
	.I(FE_PHN5063_n2383));
   BUFCKEHD FE_PHC3886_n3016 (.O(FE_PHN3886_n3016), 
	.I(n3016));
   BUFEHD FE_PHC3885_n1024 (.O(FE_PHN3885_n1024), 
	.I(n1024));
   BUFLHD FE_PHC3884_n895 (.O(FE_PHN3884_n895), 
	.I(n895));
   BUFEHD FE_PHC3883_n2163 (.O(FE_PHN3883_n2163), 
	.I(n2163));
   BUFEHD FE_PHC3882_n1023 (.O(FE_PHN3882_n1023), 
	.I(n1023));
   BUFCHD FE_PHC3881_n3129 (.O(FE_PHN3881_n3129), 
	.I(FE_PHN4348_n3129));
   BUFCHD FE_PHC3880_n2995 (.O(FE_PHN3880_n2995), 
	.I(FE_PHN4544_n2995));
   BUFHHD FE_PHC3879_n3020 (.O(FE_PHN3879_n3020), 
	.I(n3020));
   BUFEHD FE_PHC3878_n2900 (.O(FE_PHN3878_n2900), 
	.I(n2900));
   BUFEHD FE_PHC3877_n999 (.O(FE_PHN3877_n999), 
	.I(n999));
   BUFCHD FE_PHC3876_n920 (.O(FE_PHN3876_n920), 
	.I(n920));
   BUFCHD FE_PHC3875_n1006 (.O(FE_PHN3875_n1006), 
	.I(FE_PHN5306_n1006));
   BUFEHD FE_PHC3874_n2408 (.O(FE_PHN3874_n2408), 
	.I(n2408));
   BUFCHD FE_PHC3873_n3058 (.O(FE_PHN3873_n3058), 
	.I(n3058));
   BUFNHD FE_PHC3872_n873 (.O(FE_PHN3872_n873), 
	.I(n873));
   BUFNHD FE_PHC3871_n3951 (.O(FE_PHN3871_n3951), 
	.I(n3951));
   BUFEHD FE_PHC3870_n904 (.O(FE_PHN3870_n904), 
	.I(n904));
   BUFEHD FE_PHC3869_n1921 (.O(FE_PHN3869_n1921), 
	.I(n1921));
   BUFEHD FE_PHC3868_n3075 (.O(FE_PHN3868_n3075), 
	.I(n3075));
   BUFIHD FE_PHC3867_n2970 (.O(FE_PHN3867_n2970), 
	.I(n2970));
   BUFEHD FE_PHC3866_n3074 (.O(FE_PHN3866_n3074), 
	.I(n3074));
   BUFCHD FE_PHC3865_n902 (.O(FE_PHN3865_n902), 
	.I(FE_PHN5449_n902));
   BUFEHD FE_PHC3864_n1899 (.O(FE_PHN3864_n1899), 
	.I(n1899));
   BUFCHD FE_PHC3863_n844 (.O(FE_PHN3863_n844), 
	.I(FE_PHN5466_n844));
   BUFCHD FE_PHC3862_ram_31__2_ (.O(FE_PHN3862_ram_31__2_), 
	.I(\ram[31][2] ));
   BUFHHD FE_PHC3861_n905 (.O(FE_PHN3861_n905), 
	.I(n905));
   BUFEHD FE_PHC3860_n3946 (.O(FE_PHN3860_n3946), 
	.I(n3946));
   BUFHHD FE_PHC3859_n2967 (.O(FE_PHN3859_n2967), 
	.I(n2967));
   BUFEHD FE_PHC3858_n2896 (.O(FE_PHN3858_n2896), 
	.I(n2896));
   BUFEHD FE_PHC3857_n840 (.O(FE_PHN3857_n840), 
	.I(n840));
   BUFCHD FE_PHC3856_n2753 (.O(FE_PHN3856_n2753), 
	.I(FE_PHN4513_n2753));
   BUFCHD FE_PHC3855_n4229 (.O(FE_PHN3855_n4229), 
	.I(FE_PHN4503_n4229));
   BUFEHD FE_PHC3854_ram_238__0_ (.O(FE_PHN3854_ram_238__0_), 
	.I(\ram[238][0] ));
   BUFCHD FE_PHC3853_n1874 (.O(FE_PHN3853_n1874), 
	.I(n1874));
   BUFJHD FE_PHC3852_n2916 (.O(FE_PHN3852_n2916), 
	.I(n2916));
   BUFCHD FE_PHC3851_n3119 (.O(FE_PHN3851_n3119), 
	.I(n3119));
   BUFHHD FE_PHC3850_n3109 (.O(FE_PHN3850_n3109), 
	.I(n3109));
   BUFEHD FE_PHC3849_n3054 (.O(FE_PHN3849_n3054), 
	.I(n3054));
   BUFCKEHD FE_PHC3848_n4397 (.O(FE_PHN3848_n4397), 
	.I(n4397));
   BUFCHD FE_PHC3847_n934 (.O(FE_PHN3847_n934), 
	.I(n934));
   BUFEHD FE_PHC3846_n913 (.O(FE_PHN3846_n913), 
	.I(n913));
   BUFEHD FE_PHC3845_n952 (.O(FE_PHN3845_n952), 
	.I(n952));
   BUFCHD FE_PHC3844_n4227 (.O(FE_PHN3844_n4227), 
	.I(FE_PHN5558_n4227));
   BUFEHD FE_PHC3843_n2986 (.O(FE_PHN3843_n2986), 
	.I(n2986));
   BUFCHD FE_PHC3842_n1079 (.O(FE_PHN3842_n1079), 
	.I(n1079));
   BUFCHD FE_PHC3841_n3060 (.O(FE_PHN3841_n3060), 
	.I(n3060));
   BUFCHD FE_PHC3840_n1922 (.O(FE_PHN3840_n1922), 
	.I(FE_PHN6491_n1922));
   BUFCKEHD FE_PHC3839_n2384 (.O(FE_PHN3839_n2384), 
	.I(n2384));
   BUFEHD FE_PHC3838_n3090 (.O(FE_PHN3838_n3090), 
	.I(n3090));
   BUFCHD FE_PHC3837_n3029 (.O(FE_PHN3837_n3029), 
	.I(n3029));
   BUFEHD FE_PHC3836_n906 (.O(FE_PHN3836_n906), 
	.I(n906));
   BUFEHD FE_PHC3835_n3262 (.O(FE_PHN3835_n3262), 
	.I(n3262));
   BUFJHD FE_PHC3834_n4209 (.O(FE_PHN3834_n4209), 
	.I(n4209));
   BUFEHD FE_PHC3833_n1880 (.O(FE_PHN3833_n1880), 
	.I(n1880));
   BUFEHD FE_PHC3832_n949 (.O(FE_PHN3832_n949), 
	.I(n949));
   BUFCKEHD FE_PHC3831_n1906 (.O(FE_PHN3831_n1906), 
	.I(n1906));
   BUFCKEHD FE_PHC3830_n3015 (.O(FE_PHN3830_n3015), 
	.I(n3015));
   BUFHHD FE_PHC3829_n1021 (.O(FE_PHN3829_n1021), 
	.I(n1021));
   BUFEHD FE_PHC3828_n4400 (.O(FE_PHN3828_n4400), 
	.I(n4400));
   BUFCHD FE_PHC3827_n959 (.O(FE_PHN3827_n959), 
	.I(n959));
   BUFCKJHD FE_PHC3826_n2943 (.O(FE_PHN3826_n2943), 
	.I(n2943));
   BUFCHD FE_PHC3825_n4283 (.O(FE_PHN3825_n4283), 
	.I(n4283));
   BUFMHD FE_PHC3824_n4265 (.O(FE_PHN3824_n4265), 
	.I(n4265));
   BUFCHD FE_PHC3823_n4134 (.O(FE_PHN3823_n4134), 
	.I(FE_PHN5524_n4134));
   BUFMHD FE_PHC3822_n4366 (.O(FE_PHN3822_n4366), 
	.I(n4366));
   BUFHHD FE_PHC3821_n2574 (.O(FE_PHN3821_n2574), 
	.I(n2574));
   BUFCKEHD FE_PHC3820_n1030 (.O(FE_PHN3820_n1030), 
	.I(n1030));
   BUFCHD FE_PHC3819_n3994 (.O(FE_PHN3819_n3994), 
	.I(n3994));
   BUFEHD FE_PHC3818_n4111 (.O(FE_PHN3818_n4111), 
	.I(n4111));
   BUFEHD FE_PHC3817_n1916 (.O(FE_PHN3817_n1916), 
	.I(n1916));
   BUFHHD FE_PHC3816_n1037 (.O(FE_PHN3816_n1037), 
	.I(n1037));
   BUFHHD FE_PHC3815_n3963 (.O(FE_PHN3815_n3963), 
	.I(n3963));
   BUFEHD FE_PHC3814_n1896 (.O(FE_PHN3814_n1896), 
	.I(n1896));
   BUFEHD FE_PHC3813_n888 (.O(FE_PHN3813_n888), 
	.I(n888));
   BUFLHD FE_PHC3812_n3210 (.O(FE_PHN3812_n3210), 
	.I(n3210));
   BUFCKEHD FE_PHC3811_n841 (.O(FE_PHN3811_n841), 
	.I(n841));
   BUFEHD FE_PHC3810_n2962 (.O(FE_PHN3810_n2962), 
	.I(n2962));
   BUFEHD FE_PHC3809_n2437 (.O(FE_PHN3809_n2437), 
	.I(n2437));
   BUFEHD FE_PHC3808_n4291 (.O(FE_PHN3808_n4291), 
	.I(n4291));
   BUFLHD FE_PHC3807_n3062 (.O(FE_PHN3807_n3062), 
	.I(n3062));
   BUFCHD FE_PHC3806_n845 (.O(FE_PHN3806_n845), 
	.I(n845));
   BUFNHD FE_PHC3805_n2990 (.O(FE_PHN3805_n2990), 
	.I(n2990));
   BUFEHD FE_PHC3804_n4037 (.O(FE_PHN3804_n4037), 
	.I(n4037));
   BUFJHD FE_PHC3803_n962 (.O(FE_PHN3803_n962), 
	.I(n962));
   BUFCHD FE_PHC3802_n1038 (.O(FE_PHN3802_n1038), 
	.I(n1038));
   BUFKHD FE_PHC3801_n3916 (.O(FE_PHN3801_n3916), 
	.I(n3916));
   BUFCKEHD FE_PHC3800_n4231 (.O(FE_PHN3800_n4231), 
	.I(n4231));
   BUFCHD FE_PHC3799_n3942 (.O(FE_PHN3799_n3942), 
	.I(n3942));
   BUFEHD FE_PHC3798_n3968 (.O(FE_PHN3798_n3968), 
	.I(n3968));
   BUFEHD FE_PHC3797_n4362 (.O(FE_PHN3797_n4362), 
	.I(n4362));
   BUFEHD FE_PHC3796_n1077 (.O(FE_PHN3796_n1077), 
	.I(n1077));
   BUFMHD FE_PHC3795_n3940 (.O(FE_PHN3795_n3940), 
	.I(n3940));
   BUFHHD FE_PHC3794_n4277 (.O(FE_PHN3794_n4277), 
	.I(n4277));
   BUFEHD FE_PHC3793_n3046 (.O(FE_PHN3793_n3046), 
	.I(n3046));
   BUFEHD FE_PHC3792_n1919 (.O(FE_PHN3792_n1919), 
	.I(n1919));
   BUFCKEHD FE_PHC3791_n1002 (.O(FE_PHN3791_n1002), 
	.I(n1002));
   BUFEHD FE_PHC3790_n910 (.O(FE_PHN3790_n910), 
	.I(n910));
   BUFEHD FE_PHC3789_n965 (.O(FE_PHN3789_n965), 
	.I(n965));
   BUFMHD FE_PHC3788_n3956 (.O(FE_PHN3788_n3956), 
	.I(n3956));
   BUFEHD FE_PHC3787_n3019 (.O(FE_PHN3787_n3019), 
	.I(n3019));
   BUFCKEHD FE_PHC3786_n4158 (.O(FE_PHN3786_n4158), 
	.I(n4158));
   BUFEHD FE_PHC3785_n2898 (.O(FE_PHN3785_n2898), 
	.I(n2898));
   BUFCHD FE_PHC3784_n853 (.O(FE_PHN3784_n853), 
	.I(n853));
   BUFCHD FE_PHC3783_n943 (.O(FE_PHN3783_n943), 
	.I(n943));
   BUFEHD FE_PHC3782_n2415 (.O(FE_PHN3782_n2415), 
	.I(n2415));
   BUFNHD FE_PHC3781_n4076 (.O(FE_PHN3781_n4076), 
	.I(n4076));
   BUFEHD FE_PHC3780_n3955 (.O(FE_PHN3780_n3955), 
	.I(n3955));
   BUFCHD FE_PHC3779_n3026 (.O(FE_PHN3779_n3026), 
	.I(n3026));
   BUFNHD FE_PHC3778_n2957 (.O(FE_PHN3778_n2957), 
	.I(n2957));
   BUFCKNHD FE_PHC3777_n2732 (.O(FE_PHN3777_n2732), 
	.I(n2732));
   BUFKHD FE_PHC3776_n843 (.O(FE_PHN3776_n843), 
	.I(n843));
   BUFCHD FE_PHC3775_n3965 (.O(FE_PHN3775_n3965), 
	.I(FE_PHN5698_n3965));
   BUFCHD FE_PHC3774_n3932 (.O(FE_PHN3774_n3932), 
	.I(FE_PHN4670_n3932));
   BUFMHD FE_PHC3773_n4207 (.O(FE_PHN3773_n4207), 
	.I(n4207));
   BUFEHD FE_PHC3772_n3110 (.O(FE_PHN3772_n3110), 
	.I(n3110));
   BUFIHD FE_PHC3771_n880 (.O(FE_PHN3771_n880), 
	.I(n880));
   BUFCKEHD FE_PHC3770_n4409 (.O(FE_PHN3770_n4409), 
	.I(n4409));
   BUFCHD FE_PHC3769_n2598 (.O(FE_PHN3769_n2598), 
	.I(n2598));
   BUFEHD FE_PHC3768_n3077 (.O(FE_PHN3768_n3077), 
	.I(n3077));
   BUFEHD FE_PHC3767_n947 (.O(FE_PHN3767_n947), 
	.I(n947));
   BUFCHD FE_PHC3766_n2897 (.O(FE_PHN3766_n2897), 
	.I(n2897));
   BUFEHD FE_PHC3765_n2975 (.O(FE_PHN3765_n2975), 
	.I(n2975));
   BUFEHD FE_PHC3764_n1902 (.O(FE_PHN3764_n1902), 
	.I(n1902));
   BUFEHD FE_PHC3763_n1873 (.O(FE_PHN3763_n1873), 
	.I(n1873));
   BUFEHD FE_PHC3762_n2958 (.O(FE_PHN3762_n2958), 
	.I(n2958));
   BUFJHD FE_PHC3761_n3126 (.O(FE_PHN3761_n3126), 
	.I(n3126));
   BUFEHD FE_PHC3760_n1864 (.O(FE_PHN3760_n1864), 
	.I(n1864));
   BUFCHD FE_PHC3759_n3028 (.O(FE_PHN3759_n3028), 
	.I(FE_PHN4646_n3028));
   BUFEHD FE_PHC3758_n3042 (.O(FE_PHN3758_n3042), 
	.I(n3042));
   BUFCHD FE_PHC3757_n919 (.O(FE_PHN3757_n919), 
	.I(n919));
   BUFEHD FE_PHC3756_n2969 (.O(FE_PHN3756_n2969), 
	.I(n2969));
   BUFHHD FE_PHC3755_n4172 (.O(FE_PHN3755_n4172), 
	.I(n4172));
   BUFEHD FE_PHC3754_n2922 (.O(FE_PHN3754_n2922), 
	.I(n2922));
   BUFCHD FE_PHC3753_n4218 (.O(FE_PHN3753_n4218), 
	.I(n4218));
   BUFEHD FE_PHC3752_n1905 (.O(FE_PHN3752_n1905), 
	.I(n1905));
   BUFCKEHD FE_PHC3751_n3989 (.O(FE_PHN3751_n3989), 
	.I(n3989));
   BUFCKEHD FE_PHC3750_n4035 (.O(FE_PHN3750_n4035), 
	.I(n4035));
   BUFCHD FE_PHC3749_n3005 (.O(FE_PHN3749_n3005), 
	.I(FE_PHN5583_n3005));
   BUFCKEHD FE_PHC3748_n4062 (.O(FE_PHN3748_n4062), 
	.I(n4062));
   BUFJHD FE_PHC3747_n4222 (.O(FE_PHN3747_n4222), 
	.I(n4222));
   BUFCHD FE_PHC3746_n3040 (.O(FE_PHN3746_n3040), 
	.I(FE_PHN4629_n3040));
   BUFCHD FE_PHC3745_n1020 (.O(FE_PHN3745_n1020), 
	.I(FE_PHN5408_n1020));
   BUFEHD FE_PHC3744_n928 (.O(FE_PHN3744_n928), 
	.I(n928));
   BUFCHD FE_PHC3743_n3069 (.O(FE_PHN3743_n3069), 
	.I(n3069));
   BUFCHD FE_PHC3742_n4027 (.O(FE_PHN3742_n4027), 
	.I(n4027));
   BUFJHD FE_PHC3741_n3980 (.O(FE_PHN3741_n3980), 
	.I(n3980));
   BUFEHD FE_PHC3740_n3012 (.O(FE_PHN3740_n3012), 
	.I(n3012));
   BUFEHD FE_PHC3739_n3084 (.O(FE_PHN3739_n3084), 
	.I(n3084));
   BUFEHD FE_PHC3738_n3000 (.O(FE_PHN3738_n3000), 
	.I(n3000));
   BUFEHD FE_PHC3737_n2991 (.O(FE_PHN3737_n2991), 
	.I(n2991));
   BUFHHD FE_PHC3736_n2997 (.O(FE_PHN3736_n2997), 
	.I(n2997));
   BUFCHD FE_PHC3735_n4255 (.O(FE_PHN3735_n4255), 
	.I(n4255));
   BUFEHD FE_PHC3734_n978 (.O(FE_PHN3734_n978), 
	.I(n978));
   BUFEHD FE_PHC3733_n2982 (.O(FE_PHN3733_n2982), 
	.I(n2982));
   BUFEHD FE_PHC3732_n872 (.O(FE_PHN3732_n872), 
	.I(n872));
   BUFMHD FE_PHC3731_n4236 (.O(FE_PHN3731_n4236), 
	.I(n4236));
   BUFEHD FE_PHC3730_n3007 (.O(FE_PHN3730_n3007), 
	.I(n3007));
   BUFEHD FE_PHC3729_n2961 (.O(FE_PHN3729_n2961), 
	.I(n2961));
   BUFMHD FE_PHC3728_n4395 (.O(FE_PHN3728_n4395), 
	.I(n4395));
   BUFCKEHD FE_PHC3727_n1029 (.O(FE_PHN3727_n1029), 
	.I(n1029));
   BUFIHD FE_PHC3726_n903 (.O(FE_PHN3726_n903), 
	.I(n903));
   BUFEHD FE_PHC3725_n1072 (.O(FE_PHN3725_n1072), 
	.I(n1072));
   BUFEHD FE_PHC3724_n3926 (.O(FE_PHN3724_n3926), 
	.I(n3926));
   BUFHHD FE_PHC3723_n972 (.O(FE_PHN3723_n972), 
	.I(n972));
   BUFCHD FE_PHC3722_ram_154__5_ (.O(FE_PHN3722_ram_154__5_), 
	.I(\ram[154][5] ));
   BUFIHD FE_PHC3721_n4049 (.O(FE_PHN3721_n4049), 
	.I(n4049));
   BUFEHD FE_PHC3720_n3966 (.O(FE_PHN3720_n3966), 
	.I(n3966));
   BUFEHD FE_PHC3719_n3083 (.O(FE_PHN3719_n3083), 
	.I(n3083));
   BUFLHD FE_PHC3718_n2928 (.O(FE_PHN3718_n2928), 
	.I(n2928));
   BUFJHD FE_PHC3717_n1920 (.O(FE_PHN3717_n1920), 
	.I(n1920));
   BUFCHD FE_PHC3716_n1904 (.O(FE_PHN3716_n1904), 
	.I(FE_PHN5055_n1904));
   BUFCHD FE_PHC3715_n1106 (.O(FE_PHN3715_n1106), 
	.I(FE_PHN5276_n1106));
   BUFCKNHD FE_PHC3714_n4175 (.O(FE_PHN3714_n4175), 
	.I(n4175));
   BUFCHD FE_PHC3713_n4103 (.O(FE_PHN3713_n4103), 
	.I(FE_PHN5554_n4103));
   BUFIHD FE_PHC3712_n3136 (.O(FE_PHN3712_n3136), 
	.I(n3136));
   BUFEHD FE_PHC3711_n991 (.O(FE_PHN3711_n991), 
	.I(n991));
   BUFCHD FE_PHC3710_n3921 (.O(FE_PHN3710_n3921), 
	.I(n3921));
   BUFEHD FE_PHC3709_n925 (.O(FE_PHN3709_n925), 
	.I(n925));
   BUFEHD FE_PHC3708_n941 (.O(FE_PHN3708_n941), 
	.I(n941));
   BUFEHD FE_PHC3707_n2955 (.O(FE_PHN3707_n2955), 
	.I(n2955));
   BUFHHD FE_PHC3706_n2983 (.O(FE_PHN3706_n2983), 
	.I(n2983));
   BUFIHD FE_PHC3705_n4232 (.O(FE_PHN3705_n4232), 
	.I(n4232));
   BUFCKEHD FE_PHC3704_n3964 (.O(FE_PHN3704_n3964), 
	.I(FE_PHN4653_n3964));
   BUFEHD FE_PHC3703_n3070 (.O(FE_PHN3703_n3070), 
	.I(n3070));
   BUFCKNHD FE_PHC3702_n2733 (.O(FE_PHN3702_n2733), 
	.I(n2733));
   BUFIHD FE_PHC3701_n2405 (.O(FE_PHN3701_n2405), 
	.I(n2405));
   BUFHHD FE_PHC3700_n2599 (.O(FE_PHN3700_n2599), 
	.I(n2599));
   BUFCHD FE_PHC3699_n4261 (.O(FE_PHN3699_n4261), 
	.I(n4261));
   BUFCKNHD FE_PHC3698_n4170 (.O(FE_PHN3698_n4170), 
	.I(n4170));
   BUFCHD FE_PHC3697_n2968 (.O(FE_PHN3697_n2968), 
	.I(n2968));
   BUFEHD FE_PHC3696_n887 (.O(FE_PHN3696_n887), 
	.I(n887));
   BUFCHD FE_PHC3695_n1088 (.O(FE_PHN3695_n1088), 
	.I(n1088));
   BUFCKNHD FE_PHC3694_n3241 (.O(FE_PHN3694_n3241), 
	.I(FE_PHN4755_n3241));
   BUFCKEHD FE_PHC3693_n3984 (.O(FE_PHN3693_n3984), 
	.I(n3984));
   BUFEHD FE_PHC3692_n2430 (.O(FE_PHN3692_n2430), 
	.I(n2430));
   BUFCHD FE_PHC3691_ram_214__13_ (.O(FE_PHN3691_ram_214__13_), 
	.I(\ram[214][13] ));
   BUFEHD FE_PHC3690_ram_153__11_ (.O(FE_PHN3690_ram_153__11_), 
	.I(\ram[153][11] ));
   BUFHHD FE_PHC3689_n4148 (.O(FE_PHN3689_n4148), 
	.I(n4148));
   BUFCHD FE_PHC3688_n3265 (.O(FE_PHN3688_n3265), 
	.I(n3265));
   BUFCHD FE_PHC3687_n4269 (.O(FE_PHN3687_n4269), 
	.I(n4269));
   BUFCHD FE_PHC3686_n1051 (.O(FE_PHN3686_n1051), 
	.I(n1051));
   BUFCKNHD FE_PHC3685_n1068 (.O(FE_PHN3685_n1068), 
	.I(FE_PHN4767_n1068));
   BUFCHD FE_PHC3684_n871 (.O(FE_PHN3684_n871), 
	.I(n871));
   BUFCKEHD FE_PHC3683_n4308 (.O(FE_PHN3683_n4308), 
	.I(n4308));
   BUFCHD FE_PHC3682_n957 (.O(FE_PHN3682_n957), 
	.I(FE_PHN5280_n957));
   BUFCHD FE_PHC3681_n3918 (.O(FE_PHN3681_n3918), 
	.I(FE_PHN5450_n3918));
   BUFCKEHD FE_PHC3680_n4016 (.O(FE_PHN3680_n4016), 
	.I(n4016));
   BUFCHD FE_PHC3679_n3072 (.O(FE_PHN3679_n3072), 
	.I(FE_PHN4493_n3072));
   BUFCKEHD FE_PHC3678_n4181 (.O(FE_PHN3678_n4181), 
	.I(n4181));
   BUFCKEHD FE_PHC3677_n2960 (.O(FE_PHN3677_n2960), 
	.I(n2960));
   BUFCHD FE_PHC3676_n1082 (.O(FE_PHN3676_n1082), 
	.I(FE_PHN4533_n1082));
   BUFCHD FE_PHC3675_n4204 (.O(FE_PHN3675_n4204), 
	.I(n4204));
   BUFCHD FE_PHC3674_n4290 (.O(FE_PHN3674_n4290), 
	.I(n4290));
   BUFEHD FE_PHC3673_n1069 (.O(FE_PHN3673_n1069), 
	.I(n1069));
   BUFCKNHD FE_PHC3672_n1027 (.O(FE_PHN3672_n1027), 
	.I(FE_PHN4773_n1027));
   BUFEHD FE_PHC3671_n3006 (.O(FE_PHN3671_n3006), 
	.I(n3006));
   BUFCHD FE_PHC3670_n950 (.O(FE_PHN3670_n950), 
	.I(n950));
   BUFHHD FE_PHC3669_n3013 (.O(FE_PHN3669_n3013), 
	.I(n3013));
   BUFEHD FE_PHC3668_n852 (.O(FE_PHN3668_n852), 
	.I(n852));
   BUFCKEHD FE_PHC3667_n4365 (.O(FE_PHN3667_n4365), 
	.I(n4365));
   BUFHHD FE_PHC3666_n2998 (.O(FE_PHN3666_n2998), 
	.I(n2998));
   BUFJHD FE_PHC3665_n4178 (.O(FE_PHN3665_n4178), 
	.I(n4178));
   BUFEHD FE_PHC3664_n842 (.O(FE_PHN3664_n842), 
	.I(n842));
   BUFEHD FE_PHC3663_n2953 (.O(FE_PHN3663_n2953), 
	.I(n2953));
   BUFEHD FE_PHC3662_n3978 (.O(FE_PHN3662_n3978), 
	.I(n3978));
   BUFEHD FE_PHC3661_n4007 (.O(FE_PHN3661_n4007), 
	.I(n4007));
   BUFLHD FE_PHC3660_n839 (.O(FE_PHN3660_n839), 
	.I(n839));
   BUFEHD FE_PHC3659_n1040 (.O(FE_PHN3659_n1040), 
	.I(n1040));
   BUFEHD FE_PHC3658_n1087 (.O(FE_PHN3658_n1087), 
	.I(n1087));
   BUFLHD FE_PHC3657_n4240 (.O(FE_PHN3657_n4240), 
	.I(n4240));
   BUFEHD FE_PHC3656_n3088 (.O(FE_PHN3656_n3088), 
	.I(n3088));
   BUFCKEHD FE_PHC3655_n4025 (.O(FE_PHN3655_n4025), 
	.I(n4025));
   BUFLHD FE_PHC3654_n863 (.O(FE_PHN3654_n863), 
	.I(n863));
   BUFJHD FE_PHC3653_n2989 (.O(FE_PHN3653_n2989), 
	.I(n2989));
   BUFEHD FE_PHC3652_n4271 (.O(FE_PHN3652_n4271), 
	.I(n4271));
   BUFHHD FE_PHC3651_n2971 (.O(FE_PHN3651_n2971), 
	.I(n2971));
   BUFEHD FE_PHC3650_n4000 (.O(FE_PHN3650_n4000), 
	.I(n4000));
   BUFEHD FE_PHC3649_n3128 (.O(FE_PHN3649_n3128), 
	.I(n3128));
   BUFCHD FE_PHC3648_n3056 (.O(FE_PHN3648_n3056), 
	.I(n3056));
   BUFCHD FE_PHC3647_n992 (.O(FE_PHN3647_n992), 
	.I(n992));
   BUFCHD FE_PHC3646_n2985 (.O(FE_PHN3646_n2985), 
	.I(n2985));
   BUFLHD FE_PHC3645_n4329 (.O(FE_PHN3645_n4329), 
	.I(n4329));
   BUFCHD FE_PHC3644_n4213 (.O(FE_PHN3644_n4213), 
	.I(FE_PHN5549_n4213));
   BUFCHD FE_PHC3643_n4415 (.O(FE_PHN3643_n4415), 
	.I(FE_PHN5304_n4415));
   BUFJHD FE_PHC3642_n3086 (.O(FE_PHN3642_n3086), 
	.I(n3086));
   BUFEHD FE_PHC3641_ram_144__8_ (.O(FE_PHN3641_ram_144__8_), 
	.I(\ram[144][8] ));
   BUFCHD FE_PHC3640_n3023 (.O(FE_PHN3640_n3023), 
	.I(n3023));
   BUFKHD FE_PHC3639_n2420 (.O(FE_PHN3639_n2420), 
	.I(n2420));
   BUFEHD FE_PHC3638_n4279 (.O(FE_PHN3638_n4279), 
	.I(n4279));
   BUFEHD FE_PHC3637_n3133 (.O(FE_PHN3637_n3133), 
	.I(n3133));
   BUFIHD FE_PHC3636_n847 (.O(FE_PHN3636_n847), 
	.I(n847));
   BUFEHD FE_PHC3635_n2399 (.O(FE_PHN3635_n2399), 
	.I(n2399));
   BUFEHD FE_PHC3634_n4009 (.O(FE_PHN3634_n4009), 
	.I(n4009));
   BUFEHD FE_PHC3633_n922 (.O(FE_PHN3633_n922), 
	.I(n922));
   BUFMHD FE_PHC3632_n4267 (.O(FE_PHN3632_n4267), 
	.I(n4267));
   BUFEHD FE_PHC3631_n3055 (.O(FE_PHN3631_n3055), 
	.I(n3055));
   BUFCHD FE_PHC3630_n4219 (.O(FE_PHN3630_n4219), 
	.I(FE_PHN4604_n4219));
   BUFCHD FE_PHC3629_n3112 (.O(FE_PHN3629_n3112), 
	.I(n3112));
   BUFCHD FE_PHC3628_n4274 (.O(FE_PHN3628_n4274), 
	.I(n4274));
   BUFCHD FE_PHC3627_n4245 (.O(FE_PHN3627_n4245), 
	.I(n4245));
   BUFCKNHD FE_PHC3626_n1206 (.O(FE_PHN3626_n1206), 
	.I(n1206));
   BUFCHD FE_PHC3625_n1025 (.O(FE_PHN3625_n1025), 
	.I(n1025));
   BUFCHD FE_PHC3624_n4239 (.O(FE_PHN3624_n4239), 
	.I(n4239));
   BUFCHD FE_PHC3623_n1018 (.O(FE_PHN3623_n1018), 
	.I(FE_PHN5272_n1018));
   BUFCHD FE_PHC3622_n2754 (.O(FE_PHN3622_n2754), 
	.I(FE_PHN5335_n2754));
   BUFEHD FE_PHC3621_n4367 (.O(FE_PHN3621_n4367), 
	.I(n4367));
   BUFCKEHD FE_PHC3620_n4392 (.O(FE_PHN3620_n4392), 
	.I(n4392));
   BUFEHD FE_PHC3619_n909 (.O(FE_PHN3619_n909), 
	.I(n909));
   BUFEHD FE_PHC3618_n3073 (.O(FE_PHN3618_n3073), 
	.I(n3073));
   BUFCHD FE_PHC3617_n2891 (.O(FE_PHN3617_n2891), 
	.I(n2891));
   BUFKHD FE_PHC3616_n3098 (.O(FE_PHN3616_n3098), 
	.I(n3098));
   BUFEHD FE_PHC3615_n4316 (.O(FE_PHN3615_n4316), 
	.I(n4316));
   BUFEHD FE_PHC3614_n3003 (.O(FE_PHN3614_n3003), 
	.I(n3003));
   BUFCKNHD FE_PHC3613_n2262 (.O(FE_PHN3613_n2262), 
	.I(FE_PHN4769_n2262));
   BUFCHD FE_PHC3612_n3024 (.O(FE_PHN3612_n3024), 
	.I(FE_PHN5409_n3024));
   BUFCHD FE_PHC3611_n4382 (.O(FE_PHN3611_n4382), 
	.I(FE_PHN5561_n4382));
   BUFHHD FE_PHC3610_n4334 (.O(FE_PHN3610_n4334), 
	.I(n4334));
   BUFCKEHD FE_PHC3609_n3117 (.O(FE_PHN3609_n3117), 
	.I(n3117));
   BUFHHD FE_PHC3608_n2996 (.O(FE_PHN3608_n2996), 
	.I(n2996));
   BUFCKEHD FE_PHC3607_n2432 (.O(FE_PHN3607_n2432), 
	.I(n2432));
   BUFCKEHD FE_PHC3606_n4116 (.O(FE_PHN3606_n4116), 
	.I(n4116));
   BUFCHD FE_PHC3605_n2403 (.O(FE_PHN3605_n2403), 
	.I(FE_PHN6457_n2403));
   BUFMHD FE_PHC3604_n4171 (.O(FE_PHN3604_n4171), 
	.I(n4171));
   BUFCHD FE_PHC3603_n1009 (.O(FE_PHN3603_n1009), 
	.I(n1009));
   BUFCKNHD FE_PHC3602_n2727 (.O(FE_PHN3602_n2727), 
	.I(n2727));
   BUFEHD FE_PHC3601_n3914 (.O(FE_PHN3601_n3914), 
	.I(n3914));
   BUFCHD FE_PHC3600_n2935 (.O(FE_PHN3600_n2935), 
	.I(n2935));
   BUFEHD FE_PHC3599_n4238 (.O(FE_PHN3599_n4238), 
	.I(n4238));
   BUFKHD FE_PHC3598_n4299 (.O(FE_PHN3598_n4299), 
	.I(n4299));
   BUFIHD FE_PHC3597_n4404 (.O(FE_PHN3597_n4404), 
	.I(n4404));
   BUFCKEHD FE_PHC3596_n4413 (.O(FE_PHN3596_n4413), 
	.I(n4413));
   BUFLHD FE_PHC3595_n911 (.O(FE_PHN3595_n911), 
	.I(n911));
   BUFCKEHD FE_PHC3594_n4228 (.O(FE_PHN3594_n4228), 
	.I(n4228));
   BUFCKEHD FE_PHC3593_ram_145__7_ (.O(FE_PHN3593_ram_145__7_), 
	.I(\ram[145][7] ));
   BUFCHD FE_PHC3592_n3982 (.O(FE_PHN3592_n3982), 
	.I(n3982));
   BUFNHD FE_PHC3591_n3950 (.O(FE_PHN3591_n3950), 
	.I(n3950));
   BUFCHD FE_PHC3590_n3102 (.O(FE_PHN3590_n3102), 
	.I(n3102));
   BUFCKEHD FE_PHC3589_n4188 (.O(FE_PHN3589_n4188), 
	.I(n4188));
   BUFEHD FE_PHC3588_n3134 (.O(FE_PHN3588_n3134), 
	.I(n3134));
   BUFEHD FE_PHC3587_n3971 (.O(FE_PHN3587_n3971), 
	.I(n3971));
   BUFHHD FE_PHC3586_n3263 (.O(FE_PHN3586_n3263), 
	.I(n3263));
   BUFEHD FE_PHC3585_n964 (.O(FE_PHN3585_n964), 
	.I(n964));
   BUFEHD FE_PHC3584_n2994 (.O(FE_PHN3584_n2994), 
	.I(n2994));
   BUFEHD FE_PHC3583_n3027 (.O(FE_PHN3583_n3027), 
	.I(n3027));
   BUFEHD FE_PHC3582_n4371 (.O(FE_PHN3582_n4371), 
	.I(n4371));
   BUFEHD FE_PHC3581_n4359 (.O(FE_PHN3581_n4359), 
	.I(n4359));
   BUFIHD FE_PHC3580_n2951 (.O(FE_PHN3580_n2951), 
	.I(n2951));
   BUFCHD FE_PHC3579_n901 (.O(FE_PHN3579_n901), 
	.I(n901));
   BUFIHD FE_PHC3578_n3992 (.O(FE_PHN3578_n3992), 
	.I(n3992));
   BUFEHD FE_PHC3577_n2978 (.O(FE_PHN3577_n2978), 
	.I(n2978));
   BUFCKEHD FE_PHC3576_n3091 (.O(FE_PHN3576_n3091), 
	.I(n3091));
   BUFJHD FE_PHC3575_n3044 (.O(FE_PHN3575_n3044), 
	.I(n3044));
   BUFHHD FE_PHC3574_n4294 (.O(FE_PHN3574_n4294), 
	.I(n4294));
   BUFIHD FE_PHC3573_n935 (.O(FE_PHN3573_n935), 
	.I(n935));
   BUFCHD FE_PHC3572_n2992 (.O(FE_PHN3572_n2992), 
	.I(FE_PHN5333_n2992));
   BUFCHD FE_PHC3571_ram_133__9_ (.O(FE_PHN3571_ram_133__9_), 
	.I(\ram[133][9] ));
   BUFCHD FE_PHC3570_n890 (.O(FE_PHN3570_n890), 
	.I(n890));
   BUFCHD FE_PHC3569_n998 (.O(FE_PHN3569_n998), 
	.I(FE_PHN5020_n998));
   BUFCHD FE_PHC3568_n997 (.O(FE_PHN3568_n997), 
	.I(n997));
   BUFEHD FE_PHC3567_n2431 (.O(FE_PHN3567_n2431), 
	.I(n2431));
   BUFEHD FE_PHC3566_n927 (.O(FE_PHN3566_n927), 
	.I(n927));
   BUFCHD FE_PHC3565_n3970 (.O(FE_PHN3565_n3970), 
	.I(FE_PHN4514_n3970));
   BUFCKMHD FE_PHC3564_n3917 (.O(FE_PHN3564_n3917), 
	.I(n3917));
   BUFMHD FE_PHC3563_n1066 (.O(FE_PHN3563_n1066), 
	.I(n1066));
   BUFCKEHD FE_PHC3562_n3095 (.O(FE_PHN3562_n3095), 
	.I(n3095));
   BUFCKEHD FE_PHC3561_n3911 (.O(FE_PHN3561_n3911), 
	.I(n3911));
   BUFCHD FE_PHC3560_n989 (.O(FE_PHN3560_n989), 
	.I(FE_PHN5124_n989));
   BUFEHD FE_PHC3559_n3009 (.O(FE_PHN3559_n3009), 
	.I(n3009));
   BUFCKEHD FE_PHC3558_n3132 (.O(FE_PHN3558_n3132), 
	.I(n3132));
   BUFJHD FE_PHC3557_n874 (.O(FE_PHN3557_n874), 
	.I(n874));
   BUFIHD FE_PHC3556_n2987 (.O(FE_PHN3556_n2987), 
	.I(n2987));
   BUFCHD FE_PHC3555_n849 (.O(FE_PHN3555_n849), 
	.I(n849));
   BUFJHD FE_PHC3554_n2927 (.O(FE_PHN3554_n2927), 
	.I(n2927));
   BUFCHD FE_PHC3553_n3137 (.O(FE_PHN3553_n3137), 
	.I(FE_PHN4507_n3137));
   BUFEHD FE_PHC3552_n2389 (.O(FE_PHN3552_n2389), 
	.I(n2389));
   BUFJHD FE_PHC3551_n1870 (.O(FE_PHN3551_n1870), 
	.I(n1870));
   BUFJHD FE_PHC3550_n4226 (.O(FE_PHN3550_n4226), 
	.I(n4226));
   BUFHHD FE_PHC3549_n3018 (.O(FE_PHN3549_n3018), 
	.I(n3018));
   BUFIHD FE_PHC3548_n4364 (.O(FE_PHN3548_n4364), 
	.I(n4364));
   BUFCKEHD FE_PHC3547_n3140 (.O(FE_PHN3547_n3140), 
	.I(n3140));
   BUFCHD FE_PHC3546_n984 (.O(FE_PHN3546_n984), 
	.I(n984));
   BUFCHD FE_PHC3545_n1048 (.O(FE_PHN3545_n1048), 
	.I(n1048));
   BUFCHD FE_PHC3544_n3010 (.O(FE_PHN3544_n3010), 
	.I(n3010));
   BUFHHD FE_PHC3543_n4169 (.O(FE_PHN3543_n4169), 
	.I(n4169));
   BUFCHD FE_PHC3542_n2932 (.O(FE_PHN3542_n2932), 
	.I(n2932));
   BUFCHD FE_PHC3541_n4179 (.O(FE_PHN3541_n4179), 
	.I(FE_PHN4610_n4179));
   BUFHHD FE_PHC3540_n4212 (.O(FE_PHN3540_n4212), 
	.I(n4212));
   BUFCKEHD FE_PHC3539_n4295 (.O(FE_PHN3539_n4295), 
	.I(n4295));
   BUFHHD FE_PHC3538_n4211 (.O(FE_PHN3538_n4211), 
	.I(n4211));
   BUFCHD FE_PHC3537_n4340 (.O(FE_PHN3537_n4340), 
	.I(FE_PHN5344_n4340));
   BUFMHD FE_PHC3536_n4414 (.O(FE_PHN3536_n4414), 
	.I(n4414));
   BUFCHD FE_PHC3535_n938 (.O(FE_PHN3535_n938), 
	.I(FE_PHN4458_n938));
   BUFCKEHD FE_PHC3534_n3913 (.O(FE_PHN3534_n3913), 
	.I(n3913));
   BUFCKEHD FE_PHC3533_n897 (.O(FE_PHN3533_n897), 
	.I(n897));
   BUFCHD FE_PHC3532_n3052 (.O(FE_PHN3532_n3052), 
	.I(FE_PHN4578_n3052));
   BUFEHD FE_PHC3531_ram_229__12_ (.O(FE_PHN3531_ram_229__12_), 
	.I(\ram[229][12] ));
   BUFCKNHD FE_PHC3530_n2923 (.O(FE_PHN3530_n2923), 
	.I(n2923));
   BUFEHD FE_PHC3529_n857 (.O(FE_PHN3529_n857), 
	.I(n857));
   BUFHHD FE_PHC3528_n878 (.O(FE_PHN3528_n878), 
	.I(n878));
   BUFCHD FE_PHC3527_n975 (.O(FE_PHN3527_n975), 
	.I(FE_PHN4585_n975));
   BUFEHD FE_PHC3526_n3972 (.O(FE_PHN3526_n3972), 
	.I(n3972));
   BUFEHD FE_PHC3525_n1056 (.O(FE_PHN3525_n1056), 
	.I(n1056));
   BUFHHD FE_PHC3524_n3958 (.O(FE_PHN3524_n3958), 
	.I(n3958));
   BUFEHD FE_PHC3523_n4356 (.O(FE_PHN3523_n4356), 
	.I(n4356));
   BUFCHD FE_PHC3522_n894 (.O(FE_PHN3522_n894), 
	.I(FE_PHN5247_n894));
   BUFMHD FE_PHC3521_n4262 (.O(FE_PHN3521_n4262), 
	.I(n4262));
   BUFCHD FE_PHC3520_n3002 (.O(FE_PHN3520_n3002), 
	.I(FE_PHN5242_n3002));
   BUFEHD FE_PHC3519_ram_229__3_ (.O(FE_PHN3519_ram_229__3_), 
	.I(\ram[229][3] ));
   BUFCHD FE_PHC3518_n2980 (.O(FE_PHN3518_n2980), 
	.I(n2980));
   BUFNHD FE_PHC3517_n3952 (.O(FE_PHN3517_n3952), 
	.I(n3952));
   BUFCHD FE_PHC3516_n4034 (.O(FE_PHN3516_n4034), 
	.I(n4034));
   BUFLHD FE_PHC3515_n3258 (.O(FE_PHN3515_n3258), 
	.I(n3258));
   BUFEHD FE_PHC3514_n4369 (.O(FE_PHN3514_n4369), 
	.I(n4369));
   BUFCHD FE_PHC3513_n4220 (.O(FE_PHN3513_n4220), 
	.I(n4220));
   BUFCKEHD FE_PHC3512_n4292 (.O(FE_PHN3512_n4292), 
	.I(n4292));
   BUFEHD FE_PHC3511_n982 (.O(FE_PHN3511_n982), 
	.I(n982));
   BUFCHD FE_PHC3510_n4022 (.O(FE_PHN3510_n4022), 
	.I(n4022));
   BUFEHD FE_PHC3509_n929 (.O(FE_PHN3509_n929), 
	.I(n929));
   BUFMHD FE_PHC3508_n4233 (.O(FE_PHN3508_n4233), 
	.I(n4233));
   BUFCHD FE_PHC3507_n2400 (.O(FE_PHN3507_n2400), 
	.I(FE_PHN5109_n2400));
   BUFCKNHD FE_PHC3506_n971 (.O(FE_PHN3506_n971), 
	.I(FE_PHN4764_n971));
   BUFIHD FE_PHC3505_n4412 (.O(FE_PHN3505_n4412), 
	.I(n4412));
   BUFEHD FE_PHC3504_n914 (.O(FE_PHN3504_n914), 
	.I(n914));
   BUFEHD FE_PHC3503_n4323 (.O(FE_PHN3503_n4323), 
	.I(n4323));
   BUFCHD FE_PHC3502_ram_145__1_ (.O(FE_PHN3502_ram_145__1_), 
	.I(\ram[145][1] ));
   BUFEHD FE_PHC3501_n3923 (.O(FE_PHN3501_n3923), 
	.I(n3923));
   BUFCHD FE_PHC3500_n3948 (.O(FE_PHN3500_n3948), 
	.I(n3948));
   BUFNHD FE_PHC3499_n4087 (.O(FE_PHN3499_n4087), 
	.I(n4087));
   BUFKHD FE_PHC3498_n3945 (.O(FE_PHN3498_n3945), 
	.I(n3945));
   BUFCKNHD FE_PHC3497_n2413 (.O(FE_PHN3497_n2413), 
	.I(FE_PHN4772_n2413));
   BUFCHD FE_PHC3496_n2703 (.O(FE_PHN3496_n2703), 
	.I(FE_PHN5019_n2703));
   BUFJHD FE_PHC3495_n4284 (.O(FE_PHN3495_n4284), 
	.I(n4284));
   BUFEHD FE_PHC3494_n893 (.O(FE_PHN3494_n893), 
	.I(n893));
   BUFEHD FE_PHC3493_n4138 (.O(FE_PHN3493_n4138), 
	.I(n4138));
   BUFHHD FE_PHC3492_n882 (.O(FE_PHN3492_n882), 
	.I(n882));
   BUFHHD FE_PHC3491_n4350 (.O(FE_PHN3491_n4350), 
	.I(n4350));
   BUFCHD FE_PHC3490_n2964 (.O(FE_PHN3490_n2964), 
	.I(FE_PHN4302_n2964));
   BUFCKEHD FE_PHC3489_n3065 (.O(FE_PHN3489_n3065), 
	.I(n3065));
   BUFCHD FE_PHC3488_ram_221__1_ (.O(FE_PHN3488_ram_221__1_), 
	.I(\ram[221][1] ));
   BUFCHD FE_PHC3487_n899 (.O(FE_PHN3487_n899), 
	.I(n899));
   BUFCHD FE_PHC3486_n2374 (.O(FE_PHN3486_n2374), 
	.I(n2374));
   BUFCKEHD FE_PHC3485_n3089 (.O(FE_PHN3485_n3089), 
	.I(n3089));
   BUFCKNHD FE_PHC3484_n2600 (.O(FE_PHN3484_n2600), 
	.I(n2600));
   BUFCKEHD FE_PHC3483_n4331 (.O(FE_PHN3483_n4331), 
	.I(n4331));
   BUFCHD FE_PHC3482_n2906 (.O(FE_PHN3482_n2906), 
	.I(FE_PHN4975_n2906));
   BUFCKEHD FE_PHC3481_n3078 (.O(FE_PHN3481_n3078), 
	.I(n3078));
   BUFCKEHD FE_PHC3480_n4266 (.O(FE_PHN3480_n4266), 
	.I(n4266));
   BUFCKEHD FE_PHC3479_n4418 (.O(FE_PHN3479_n4418), 
	.I(n4418));
   BUFEHD FE_PHC3478_n2981 (.O(FE_PHN3478_n2981), 
	.I(n2981));
   BUFHHD FE_PHC3477_n3910 (.O(FE_PHN3477_n3910), 
	.I(n3910));
   BUFCKEHD FE_PHC3476_n1078 (.O(FE_PHN3476_n1078), 
	.I(n1078));
   BUFEHD FE_PHC3475_n2976 (.O(FE_PHN3475_n2976), 
	.I(n2976));
   BUFEHD FE_PHC3474_n4244 (.O(FE_PHN3474_n4244), 
	.I(n4244));
   BUFEHD FE_PHC3473_n4419 (.O(FE_PHN3473_n4419), 
	.I(n4419));
   BUFEHD FE_PHC3472_n3118 (.O(FE_PHN3472_n3118), 
	.I(n3118));
   BUFIHD FE_PHC3471_n948 (.O(FE_PHN3471_n948), 
	.I(n948));
   BUFEHD FE_PHC3470_n2999 (.O(FE_PHN3470_n2999), 
	.I(n2999));
   BUFHHD FE_PHC3469_n1872 (.O(FE_PHN3469_n1872), 
	.I(n1872));
   BUFCKEHD FE_PHC3468_n3123 (.O(FE_PHN3468_n3123), 
	.I(n3123));
   BUFCKEHD FE_PHC3467_n4110 (.O(FE_PHN3467_n4110), 
	.I(n4110));
   BUFJHD FE_PHC3466_n3976 (.O(FE_PHN3466_n3976), 
	.I(n3976));
   BUFEHD FE_PHC3465_n4142 (.O(FE_PHN3465_n4142), 
	.I(n4142));
   BUFIHD FE_PHC3464_n877 (.O(FE_PHN3464_n877), 
	.I(n877));
   BUFEHD FE_PHC3463_n933 (.O(FE_PHN3463_n933), 
	.I(n933));
   BUFEHD FE_PHC3462_n3930 (.O(FE_PHN3462_n3930), 
	.I(n3930));
   BUFEHD FE_PHC3461_n3096 (.O(FE_PHN3461_n3096), 
	.I(n3096));
   BUFCHD FE_PHC3460_n4285 (.O(FE_PHN3460_n4285), 
	.I(FE_PHN5176_n4285));
   BUFJHD FE_PHC3459_n4278 (.O(FE_PHN3459_n4278), 
	.I(n4278));
   BUFCKEHD FE_PHC3458_n4327 (.O(FE_PHN3458_n4327), 
	.I(n4327));
   BUFJHD FE_PHC3457_n4396 (.O(FE_PHN3457_n4396), 
	.I(n4396));
   BUFCKEHD FE_PHC3456_n4378 (.O(FE_PHN3456_n4378), 
	.I(n4378));
   BUFCKEHD FE_PHC3455_n4394 (.O(FE_PHN3455_n4394), 
	.I(n4394));
   BUFCHD FE_PHC3454_n1017 (.O(FE_PHN3454_n1017), 
	.I(FE_PHN4494_n1017));
   BUFKHD FE_PHC3453_n3131 (.O(FE_PHN3453_n3131), 
	.I(n3131));
   BUFCKEHD FE_PHC3452_n2131 (.O(FE_PHN3452_n2131), 
	.I(n2131));
   BUFEHD FE_PHC3451_ram_17__14_ (.O(FE_PHN3451_ram_17__14_), 
	.I(\ram[17][14] ));
   BUFCHD FE_PHC3450_n3944 (.O(FE_PHN3450_n3944), 
	.I(n3944));
   BUFKHD FE_PHC3449_n3924 (.O(FE_PHN3449_n3924), 
	.I(n3924));
   BUFNHD FE_PHC3448_n2974 (.O(FE_PHN3448_n2974), 
	.I(n2974));
   BUFEHD FE_PHC3447_n4399 (.O(FE_PHN3447_n4399), 
	.I(n4399));
   BUFCKEHD FE_PHC3446_n4023 (.O(FE_PHN3446_n4023), 
	.I(n4023));
   BUFCHD FE_PHC3445_n2972 (.O(FE_PHN3445_n2972), 
	.I(FE_PHN6692_n2972));
   BUFCKNHD FE_PHC3444_n2926 (.O(FE_PHN3444_n2926), 
	.I(FE_PHN4766_n2926));
   BUFCKEHD FE_PHC3443_n4026 (.O(FE_PHN3443_n4026), 
	.I(n4026));
   BUFCHD FE_PHC3442_n3979 (.O(FE_PHN3442_n3979), 
	.I(n3979));
   BUFHHD FE_PHC3441_n861 (.O(FE_PHN3441_n861), 
	.I(n861));
   BUFCHD FE_PHC3440_n994 (.O(FE_PHN3440_n994), 
	.I(n994));
   BUFEHD FE_PHC3439_n946 (.O(FE_PHN3439_n946), 
	.I(n946));
   BUFCHD FE_PHC3438_n3127 (.O(FE_PHN3438_n3127), 
	.I(n3127));
   BUFCKEHD FE_PHC3437_n1886 (.O(FE_PHN3437_n1886), 
	.I(n1886));
   BUFCKEHD FE_PHC3436_n958 (.O(FE_PHN3436_n958), 
	.I(n958));
   BUFCHD FE_PHC3435_n2178 (.O(FE_PHN3435_n2178), 
	.I(FE_PHN5297_n2178));
   BUFCKEHD FE_PHC3434_n3103 (.O(FE_PHN3434_n3103), 
	.I(n3103));
   BUFNHD FE_PHC3433_n3008 (.O(FE_PHN3433_n3008), 
	.I(n3008));
   BUFHHD FE_PHC3432_n917 (.O(FE_PHN3432_n917), 
	.I(n917));
   BUFCHD FE_PHC3431_n1022 (.O(FE_PHN3431_n1022), 
	.I(FE_PHN5069_n1022));
   BUFEHD FE_PHC3430_n2956 (.O(FE_PHN3430_n2956), 
	.I(n2956));
   BUFCKMHD FE_PHC3429_n3936 (.O(FE_PHN3429_n3936), 
	.I(n3936));
   BUFCHD FE_PHC3428_n4260 (.O(FE_PHN3428_n4260), 
	.I(n4260));
   BUFCHD FE_PHC3427_n4360 (.O(FE_PHN3427_n4360), 
	.I(FE_PHN5292_n4360));
   BUFLHD FE_PHC3426_n2886 (.O(FE_PHN3426_n2886), 
	.I(n2886));
   BUFCKEHD FE_PHC3425_n4375 (.O(FE_PHN3425_n4375), 
	.I(n4375));
   BUFLHD FE_PHC3424_n2918 (.O(FE_PHN3424_n2918), 
	.I(n2918));
   BUFKHD FE_PHC3423_n2984 (.O(FE_PHN3423_n2984), 
	.I(n2984));
   BUFCKEHD FE_PHC3422_n3111 (.O(FE_PHN3422_n3111), 
	.I(n3111));
   BUFHHD FE_PHC3421_n3093 (.O(FE_PHN3421_n3093), 
	.I(n3093));
   BUFCKEHD FE_PHC3420_n1016 (.O(FE_PHN3420_n1016), 
	.I(n1016));
   BUFCHD FE_PHC3419_n3049 (.O(FE_PHN3419_n3049), 
	.I(FE_PHN5084_n3049));
   BUFCHD FE_PHC3418_n3048 (.O(FE_PHN3418_n3048), 
	.I(FE_PHN5212_n3048));
   BUFCKEHD FE_PHC3417_n4363 (.O(FE_PHN3417_n4363), 
	.I(n4363));
   BUFCKEHD FE_PHC3416_n3120 (.O(FE_PHN3416_n3120), 
	.I(n3120));
   BUFCHD FE_PHC3415_n4174 (.O(FE_PHN3415_n4174), 
	.I(FE_PHN4489_n4174));
   BUFHHD FE_PHC3414_n4199 (.O(FE_PHN3414_n4199), 
	.I(n4199));
   BUFCHD FE_PHC3413_n4146 (.O(FE_PHN3413_n4146), 
	.I(n4146));
   BUFEHD FE_PHC3412_n4005 (.O(FE_PHN3412_n4005), 
	.I(n4005));
   BUFEHD FE_PHC3411_n3032 (.O(FE_PHN3411_n3032), 
	.I(n3032));
   BUFEHD FE_PHC3410_n3223 (.O(FE_PHN3410_n3223), 
	.I(n3223));
   BUFKHD FE_PHC3409_n993 (.O(FE_PHN3409_n993), 
	.I(n993));
   BUFCKEHD FE_PHC3408_n1093 (.O(FE_PHN3408_n1093), 
	.I(n1093));
   BUFHHD FE_PHC3407_n3071 (.O(FE_PHN3407_n3071), 
	.I(n3071));
   BUFCKEHD FE_PHC3406_n4031 (.O(FE_PHN3406_n4031), 
	.I(n4031));
   BUFCKEHD FE_PHC3405_n1045 (.O(FE_PHN3405_n1045), 
	.I(n1045));
   BUFCHD FE_PHC3404_n2904 (.O(FE_PHN3404_n2904), 
	.I(FE_PHN6453_n2904));
   BUFCHD FE_PHC3403_n3915 (.O(FE_PHN3403_n3915), 
	.I(FE_PHN5129_n3915));
   BUFJHD FE_PHC3402_n4029 (.O(FE_PHN3402_n4029), 
	.I(n4029));
   BUFCKEHD FE_PHC3401_n930 (.O(FE_PHN3401_n930), 
	.I(n930));
   BUFEHD FE_PHC3400_n2433 (.O(FE_PHN3400_n2433), 
	.I(n2433));
   BUFCKEHD FE_PHC3399_n4206 (.O(FE_PHN3399_n4206), 
	.I(n4206));
   BUFEHD FE_PHC3398_n3022 (.O(FE_PHN3398_n3022), 
	.I(n3022));
   BUFHHD FE_PHC3397_n4017 (.O(FE_PHN3397_n4017), 
	.I(n4017));
   BUFCKEHD FE_PHC3396_n4196 (.O(FE_PHN3396_n4196), 
	.I(n4196));
   BUFCHD FE_PHC3395_n866 (.O(FE_PHN3395_n866), 
	.I(FE_PHN5355_n866));
   BUFCKEHD FE_PHC3394_n4417 (.O(FE_PHN3394_n4417), 
	.I(n4417));
   BUFCKEHD FE_PHC3393_n1008 (.O(FE_PHN3393_n1008), 
	.I(n1008));
   BUFHHD FE_PHC3392_n4030 (.O(FE_PHN3392_n4030), 
	.I(n4030));
   BUFCHD FE_PHC3391_n974 (.O(FE_PHN3391_n974), 
	.I(FE_PHN4355_n974));
   BUFCKEHD FE_PHC3390_n3212 (.O(FE_PHN3390_n3212), 
	.I(n3212));
   BUFCHD FE_PHC3389_ram_237__7_ (.O(FE_PHN3389_ram_237__7_), 
	.I(\ram[237][7] ));
   BUFEHD FE_PHC3388_n3260 (.O(FE_PHN3388_n3260), 
	.I(n3260));
   BUFLHD FE_PHC3387_n2920 (.O(FE_PHN3387_n2920), 
	.I(n2920));
   BUFCKEHD FE_PHC3386_n3108 (.O(FE_PHN3386_n3108), 
	.I(n3108));
   BUFCHD FE_PHC3385_n4421 (.O(FE_PHN3385_n4421), 
	.I(n4421));
   BUFEHD FE_PHC3384_n4372 (.O(FE_PHN3384_n4372), 
	.I(n4372));
   BUFCHD FE_PHC3383_n4201 (.O(FE_PHN3383_n4201), 
	.I(FE_PHN4495_n4201));
   BUFLHD FE_PHC3382_n4164 (.O(FE_PHN3382_n4164), 
	.I(n4164));
   BUFNHD FE_PHC3381_n3038 (.O(FE_PHN3381_n3038), 
	.I(n3038));
   BUFCKEHD FE_PHC3380_n4300 (.O(FE_PHN3380_n4300), 
	.I(n4300));
   BUFJHD FE_PHC3379_n2950 (.O(FE_PHN3379_n2950), 
	.I(n2950));
   BUFCKEHD FE_PHC3378_n4166 (.O(FE_PHN3378_n4166), 
	.I(n4166));
   BUFCKEHD FE_PHC3377_n4408 (.O(FE_PHN3377_n4408), 
	.I(n4408));
   BUFCKEHD FE_PHC3376_n848 (.O(FE_PHN3376_n848), 
	.I(n848));
   BUFCHD FE_PHC3375_n1014 (.O(FE_PHN3375_n1014), 
	.I(FE_PHN4624_n1014));
   BUFCHD FE_PHC3374_ram_158__11_ (.O(FE_PHN3374_ram_158__11_), 
	.I(\ram[158][11] ));
   BUFCHD FE_PHC3373_ram_153__7_ (.O(FE_PHN3373_ram_153__7_), 
	.I(\ram[153][7] ));
   BUFEHD FE_PHC3372_n3116 (.O(FE_PHN3372_n3116), 
	.I(n3116));
   BUFCKNHD FE_PHC3371_n2127 (.O(FE_PHN3371_n2127), 
	.I(FE_PHN4768_n2127));
   BUFJHD FE_PHC3370_n4281 (.O(FE_PHN3370_n4281), 
	.I(n4281));
   BUFCKLHD FE_PHC3369_n4235 (.O(FE_PHN3369_n4235), 
	.I(n4235));
   BUFCHD FE_PHC3368_n1090 (.O(FE_PHN3368_n1090), 
	.I(n1090));
   BUFEHD FE_PHC3367_n2977 (.O(FE_PHN3367_n2977), 
	.I(n2977));
   BUFNHD FE_PHC3366_n838 (.O(FE_PHN3366_n838), 
	.I(n838));
   BUFEHD FE_PHC3365_n960 (.O(FE_PHN3365_n960), 
	.I(n960));
   BUFCKEHD FE_PHC3364_n4270 (.O(FE_PHN3364_n4270), 
	.I(n4270));
   BUFCHD FE_PHC3363_n918 (.O(FE_PHN3363_n918), 
	.I(n918));
   BUFCHD FE_PHC3362_n3031 (.O(FE_PHN3362_n3031), 
	.I(n3031));
   BUFCKEHD FE_PHC3361_n4028 (.O(FE_PHN3361_n4028), 
	.I(n4028));
   BUFCKEHD FE_PHC3360_n4254 (.O(FE_PHN3360_n4254), 
	.I(n4254));
   BUFCKEHD FE_PHC3359_n1032 (.O(FE_PHN3359_n1032), 
	.I(n1032));
   BUFEHD FE_PHC3358_ram_145__0_ (.O(FE_PHN3358_ram_145__0_), 
	.I(\ram[145][0] ));
   BUFEHD FE_PHC3357_n4251 (.O(FE_PHN3357_n4251), 
	.I(n4251));
   BUFCHD FE_PHC3356_n3922 (.O(FE_PHN3356_n3922), 
	.I(n3922));
   BUFEHD FE_PHC3355_n4405 (.O(FE_PHN3355_n4405), 
	.I(n4405));
   BUFJHD FE_PHC3354_n4355 (.O(FE_PHN3354_n4355), 
	.I(n4355));
   BUFCHD FE_PHC3353_n4214 (.O(FE_PHN3353_n4214), 
	.I(FE_PHN5128_n4214));
   BUFCHD FE_PHC3352_n3959 (.O(FE_PHN3352_n3959), 
	.I(FE_PHN5425_n3959));
   BUFCHD FE_PHC3351_n3104 (.O(FE_PHN3351_n3104), 
	.I(FE_PHN4078_n3104));
   BUFCKEHD FE_PHC3350_n3053 (.O(FE_PHN3350_n3053), 
	.I(n3053));
   BUFHHD FE_PHC3349_n4307 (.O(FE_PHN3349_n4307), 
	.I(n4307));
   BUFCKEHD FE_PHC3348_n2930 (.O(FE_PHN3348_n2930), 
	.I(n2930));
   BUFCHD FE_PHC3347_ram_98__3_ (.O(FE_PHN3347_ram_98__3_), 
	.I(\ram[98][3] ));
   BUFCHD FE_PHC3346_n3947 (.O(FE_PHN3346_n3947), 
	.I(n3947));
   BUFEHD FE_PHC3345_n856 (.O(FE_PHN3345_n856), 
	.I(n856));
   BUFCKEHD FE_PHC3344_n3138 (.O(FE_PHN3344_n3138), 
	.I(n3138));
   BUFEHD FE_PHC3343_n2979 (.O(FE_PHN3343_n2979), 
	.I(n2979));
   BUFCKEHD FE_PHC3342_n3983 (.O(FE_PHN3342_n3983), 
	.I(n3983));
   BUFCHD FE_PHC3341_n3927 (.O(FE_PHN3341_n3927), 
	.I(FE_PHN5009_n3927));
   BUFCKEHD FE_PHC3340_n1005 (.O(FE_PHN3340_n1005), 
	.I(n1005));
   BUFCKEHD FE_PHC3339_n3124 (.O(FE_PHN3339_n3124), 
	.I(n3124));
   BUFCKEHD FE_PHC3338_n3001 (.O(FE_PHN3338_n3001), 
	.I(n3001));
   BUFEHD FE_PHC3337_n3035 (.O(FE_PHN3337_n3035), 
	.I(n3035));
   BUFCKEHD FE_PHC3336_n3115 (.O(FE_PHN3336_n3115), 
	.I(n3115));
   BUFCHD FE_PHC3335_n869 (.O(FE_PHN3335_n869), 
	.I(FE_PHN5429_n869));
   BUFCHD FE_PHC3334_n3064 (.O(FE_PHN3334_n3064), 
	.I(FE_PHN5317_n3064));
   BUFLHD FE_PHC3333_n2888 (.O(FE_PHN3333_n2888), 
	.I(n2888));
   BUFLHD FE_PHC3332_n4311 (.O(FE_PHN3332_n4311), 
	.I(n4311));
   BUFCHD FE_PHC3331_n4398 (.O(FE_PHN3331_n4398), 
	.I(FE_PHN4273_n4398));
   BUFCKNHD FE_PHC3330_n1062 (.O(FE_PHN3330_n1062), 
	.I(FE_PHN4771_n1062));
   BUFCKEHD FE_PHC3329_n3081 (.O(FE_PHN3329_n3081), 
	.I(n3081));
   BUFEHD FE_PHC3328_n3099 (.O(FE_PHN3328_n3099), 
	.I(n3099));
   BUFHHD FE_PHC3327_n4001 (.O(FE_PHN3327_n4001), 
	.I(n4001));
   BUFCKEHD FE_PHC3326_n4406 (.O(FE_PHN3326_n4406), 
	.I(n4406));
   BUFKHD FE_PHC3325_n4393 (.O(FE_PHN3325_n4393), 
	.I(n4393));
   BUFEHD FE_PHC3324_n3094 (.O(FE_PHN3324_n3094), 
	.I(n3094));
   BUFEHD FE_PHC3323_n970 (.O(FE_PHN3323_n970), 
	.I(n970));
   BUFCHD FE_PHC3322_n4342 (.O(FE_PHN3322_n4342), 
	.I(FE_PHN5227_n4342));
   BUFCHD FE_PHC3321_n4230 (.O(FE_PHN3321_n4230), 
	.I(n4230));
   BUFEHD FE_PHC3320_n2973 (.O(FE_PHN3320_n2973), 
	.I(n2973));
   BUFHHD FE_PHC3319_n4358 (.O(FE_PHN3319_n4358), 
	.I(n4358));
   BUFCKEHD FE_PHC3318_n884 (.O(FE_PHN3318_n884), 
	.I(n884));
   BUFHHD FE_PHC3317_n4194 (.O(FE_PHN3317_n4194), 
	.I(n4194));
   BUFCKEHD FE_PHC3316_n4411 (.O(FE_PHN3316_n4411), 
	.I(n4411));
   BUFCKEHD FE_PHC3315_n2988 (.O(FE_PHN3315_n2988), 
	.I(n2988));
   BUFHHD FE_PHC3314_n3988 (.O(FE_PHN3314_n3988), 
	.I(n3988));
   BUFEHD FE_PHC3313_n3937 (.O(FE_PHN3313_n3937), 
	.I(n3937));
   BUFCKEHD FE_PHC3312_n3092 (.O(FE_PHN3312_n3092), 
	.I(n3092));
   BUFJHD FE_PHC3311_n858 (.O(FE_PHN3311_n858), 
	.I(n858));
   BUFCHD FE_PHC3310_n3043 (.O(FE_PHN3310_n3043), 
	.I(FE_PHN5103_n3043));
   BUFCKEHD FE_PHC3309_n881 (.O(FE_PHN3309_n881), 
	.I(n881));
   BUFCKEHD FE_PHC3308_n865 (.O(FE_PHN3308_n865), 
	.I(n865));
   BUFCKEHD FE_PHC3307_n3961 (.O(FE_PHN3307_n3961), 
	.I(n3961));
   BUFCKEHD FE_PHC3306_n4286 (.O(FE_PHN3306_n4286), 
	.I(n4286));
   BUFCHD FE_PHC3305_n879 (.O(FE_PHN3305_n879), 
	.I(FE_PHN5122_n879));
   BUFEHD FE_PHC3304_n4377 (.O(FE_PHN3304_n4377), 
	.I(n4377));
   BUFCKEHD FE_PHC3303_n3939 (.O(FE_PHN3303_n3939), 
	.I(n3939));
   BUFCKEHD FE_PHC3302_n4263 (.O(FE_PHN3302_n4263), 
	.I(n4263));
   BUFCKEHD FE_PHC3301_n3014 (.O(FE_PHN3301_n3014), 
	.I(n3014));
   BUFCKEHD FE_PHC3300_n3105 (.O(FE_PHN3300_n3105), 
	.I(n3105));
   BUFCHD FE_PHC3299_n4180 (.O(FE_PHN3299_n4180), 
	.I(FE_PHN4429_n4180));
   BUFCKEHD FE_PHC3298_n2421 (.O(FE_PHN3298_n2421), 
	.I(n2421));
   BUFMHD FE_PHC3297_n4402 (.O(FE_PHN3297_n4402), 
	.I(n4402));
   BUFEHD FE_PHC3296_n4380 (.O(FE_PHN3296_n4380), 
	.I(n4380));
   BUFLHD FE_PHC3295_n854 (.O(FE_PHN3295_n854), 
	.I(n854));
   BUFCKEHD FE_PHC3294_n4003 (.O(FE_PHN3294_n4003), 
	.I(n4003));
   BUFCKEHD FE_PHC3293_n3919 (.O(FE_PHN3293_n3919), 
	.I(n3919));
   BUFHHD FE_PHC3292_n4386 (.O(FE_PHN3292_n4386), 
	.I(n4386));
   BUFCHD FE_PHC3291_n3934 (.O(FE_PHN3291_n3934), 
	.I(FE_PHN6676_n3934));
   BUFCKEHD FE_PHC3290_n3063 (.O(FE_PHN3290_n3063), 
	.I(n3063));
   BUFCKEHD FE_PHC3289_n3969 (.O(FE_PHN3289_n3969), 
	.I(n3969));
   BUFCKEHD FE_PHC3288_n4167 (.O(FE_PHN3288_n4167), 
	.I(n4167));
   BUFCKEHD FE_PHC3287_n4374 (.O(FE_PHN3287_n4374), 
	.I(n4374));
   BUFCKEHD FE_PHC3286_ram_145__10_ (.O(FE_PHN3286_ram_145__10_), 
	.I(\ram[145][10] ));
   BUFCKNHD FE_PHC3285_n1046 (.O(FE_PHN3285_n1046), 
	.I(n1046));
   BUFCKEHD FE_PHC3284_n4014 (.O(FE_PHN3284_n4014), 
	.I(n4014));
   BUFCKNHD FE_PHC3283_n2396 (.O(FE_PHN3283_n2396), 
	.I(FE_PHN4761_n2396));
   BUFHHD FE_PHC3282_n3087 (.O(FE_PHN3282_n3087), 
	.I(n3087));
   BUFCKEHD FE_PHC3281_n1074 (.O(FE_PHN3281_n1074), 
	.I(n1074));
   BUFHHD FE_PHC3280_n4379 (.O(FE_PHN3280_n4379), 
	.I(n4379));
   BUFCHD FE_PHC3279_n864 (.O(FE_PHN3279_n864), 
	.I(FE_PHN5213_n864));
   BUFCHD FE_PHC3278_n3954 (.O(FE_PHN3278_n3954), 
	.I(n3954));
   BUFCKEHD FE_PHC3277_n4195 (.O(FE_PHN3277_n4195), 
	.I(n4195));
   BUFCKEHD FE_PHC3276_n855 (.O(FE_PHN3276_n855), 
	.I(n855));
   BUFCKEHD FE_PHC3275_n3107 (.O(FE_PHN3275_n3107), 
	.I(n3107));
   BUFCHD FE_PHC3274_n3998 (.O(FE_PHN3274_n3998), 
	.I(n3998));
   BUFCHD FE_PHC3273_n3993 (.O(FE_PHN3273_n3993), 
	.I(n3993));
   BUFCHD FE_PHC3272_n2966 (.O(FE_PHN3272_n2966), 
	.I(n2966));
   BUFCKEHD FE_PHC3271_n3974 (.O(FE_PHN3271_n3974), 
	.I(n3974));
   BUFCKNHD FE_PHC3270_n4123 (.O(FE_PHN3270_n4123), 
	.I(FE_PHN4770_n4123));
   BUFCHD FE_PHC3269_n1013 (.O(FE_PHN3269_n1013), 
	.I(FE_PHN4549_n1013));
   BUFIHD FE_PHC3268_n4243 (.O(FE_PHN3268_n4243), 
	.I(n4243));
   BUFCKEHD FE_PHC3267_n4388 (.O(FE_PHN3267_n4388), 
	.I(n4388));
   BUFCKNHD FE_PHC3266_n2158 (.O(FE_PHN3266_n2158), 
	.I(FE_PHN4763_n2158));
   BUFCKNHD FE_PHC3265_n2910 (.O(FE_PHN3265_n2910), 
	.I(n2910));
   BUFCKEHD FE_PHC3264_n3100 (.O(FE_PHN3264_n3100), 
	.I(n3100));
   BUFHHD FE_PHC3263_n4033 (.O(FE_PHN3263_n4033), 
	.I(n4033));
   BUFCKNHD FE_PHC3262_n2141 (.O(FE_PHN3262_n2141), 
	.I(FE_PHN4760_n2141));
   BUFCKEHD FE_PHC3261_n4343 (.O(FE_PHN3261_n4343), 
	.I(n4343));
   BUFHHD FE_PHC3260_n4332 (.O(FE_PHN3260_n4332), 
	.I(n4332));
   BUFCKEHD FE_PHC3259_n3996 (.O(FE_PHN3259_n3996), 
	.I(n3996));
   BUFCKEHD FE_PHC3258_n4391 (.O(FE_PHN3258_n4391), 
	.I(n4391));
   BUFJHD FE_PHC3257_n2936 (.O(FE_PHN3257_n2936), 
	.I(n2936));
   BUFCHD FE_PHC3256_n4339 (.O(FE_PHN3256_n4339), 
	.I(FE_PHN5492_n4339));
   BUFCKEHD FE_PHC3255_n4389 (.O(FE_PHN3255_n4389), 
	.I(n4389));
   BUFCKEHD FE_PHC3254_n4384 (.O(FE_PHN3254_n4384), 
	.I(n4384));
   BUFCKEHD FE_PHC3253_n2934 (.O(FE_PHN3253_n2934), 
	.I(n2934));
   BUFEHD FE_PHC3252_n4383 (.O(FE_PHN3252_n4383), 
	.I(n4383));
   BUFCKEHD FE_PHC3251_n4010 (.O(FE_PHN3251_n4010), 
	.I(n4010));
   BUFCKEHD FE_PHC3250_n1064 (.O(FE_PHN3250_n1064), 
	.I(n1064));
   BUFCHD FE_PHC3249_n4203 (.O(FE_PHN3249_n4203), 
	.I(FE_PHN4562_n4203));
   BUFHHD FE_PHC3248_n4021 (.O(FE_PHN3248_n4021), 
	.I(n4021));
   BUFCHD FE_PHC3247_n3125 (.O(FE_PHN3247_n3125), 
	.I(n3125));
   BUFCKNHD FE_PHC3246_n2391 (.O(FE_PHN3246_n2391), 
	.I(n2391));
   BUFCKEHD FE_PHC3245_n3030 (.O(FE_PHN3245_n3030), 
	.I(n3030));
   BUFCKEHD FE_PHC3244_n3929 (.O(FE_PHN3244_n3929), 
	.I(n3929));
   BUFCKEHD FE_PHC3243_n3985 (.O(FE_PHN3243_n3985), 
	.I(n3985));
   BUFCKEHD FE_PHC3242_n1026 (.O(FE_PHN3242_n1026), 
	.I(n1026));
   BUFCKEHD FE_PHC3241_n4006 (.O(FE_PHN3241_n4006), 
	.I(n4006));
   BUFCKEHD FE_PHC3240_n3999 (.O(FE_PHN3240_n3999), 
	.I(n3999));
   BUFKHD FE_PHC3239_n4252 (.O(FE_PHN3239_n4252), 
	.I(n4252));
   BUFCKEHD FE_PHC3238_n3987 (.O(FE_PHN3238_n3987), 
	.I(n3987));
   BUFCKEHD FE_PHC3237_n4008 (.O(FE_PHN3237_n4008), 
	.I(n4008));
   BUFEHD FE_PHC3236_n4385 (.O(FE_PHN3236_n4385), 
	.I(n4385));
   BUFCKNHD FE_PHC3235_n4015 (.O(FE_PHN3235_n4015), 
	.I(n4015));
   BUFCKEHD FE_PHC3234_n3931 (.O(FE_PHN3234_n3931), 
	.I(n3931));
   BUFCKEHD FE_PHC3233_n4324 (.O(FE_PHN3233_n4324), 
	.I(n4324));
   DELCKHD FE_PHC3230_n1489 (.O(FE_PHN3230_n1489), 
	.I(n1489));
   DELCKHD FE_PHC3229_n3451 (.O(FE_PHN3229_n3451), 
	.I(n3451));
   DELDKHD FE_PHC3228_n1773 (.O(FE_PHN3228_n1773), 
	.I(n1773));
   DELDKHD FE_PHC3227_n649 (.O(FE_PHN3227_n649), 
	.I(n649));
   DELDKHD FE_PHC3226_n2005 (.O(FE_PHN3226_n2005), 
	.I(n2005));
   DELDKHD FE_PHC3225_n809 (.O(FE_PHN3225_n809), 
	.I(n809));
   DELDKHD FE_PHC3224_n713 (.O(FE_PHN3224_n713), 
	.I(n713));
   DELCKHD FE_PHC3223_n1197 (.O(FE_PHN3223_n1197), 
	.I(n1197));
   DELCKHD FE_PHC3222_n1099 (.O(FE_PHN3222_n1099), 
	.I(n1099));
   DELCKHD FE_PHC3221_n2104 (.O(FE_PHN3221_n2104), 
	.I(n2104));
   DELCKHD FE_PHC3220_n1536 (.O(FE_PHN3220_n1536), 
	.I(n1536));
   DELCKHD FE_PHC3219_n3461 (.O(FE_PHN3219_n3461), 
	.I(n3461));
   DELCKHD FE_PHC3218_n625 (.O(FE_PHN3218_n625), 
	.I(n625));
   DELDKHD FE_PHC3217_n3427 (.O(FE_PHN3217_n3427), 
	.I(n3427));
   DELDKHD FE_PHC3216_n1425 (.O(FE_PHN3216_n1425), 
	.I(n1425));
   DELDKHD FE_PHC3215_n1132 (.O(FE_PHN3215_n1132), 
	.I(n1132));
   DELDKHD FE_PHC3214_n1815 (.O(FE_PHN3214_n1815), 
	.I(n1815));
   DELCKHD FE_PHC3213_n3152 (.O(FE_PHN3213_n3152), 
	.I(n3152));
   DELCKHD FE_PHC3212_n3520 (.O(FE_PHN3212_n3520), 
	.I(n3520));
   DELCKHD FE_PHC3211_n1422 (.O(FE_PHN3211_n1422), 
	.I(n1422));
   DELCKHD FE_PHC3210_n4162 (.O(FE_PHN3210_n4162), 
	.I(n4162));
   DELCKHD FE_PHC3209_n768 (.O(FE_PHN3209_n768), 
	.I(n768));
   DELCKHD FE_PHC3208_n1688 (.O(FE_PHN3208_n1688), 
	.I(n1688));
   DELCKHD FE_PHC3207_n3284 (.O(FE_PHN3207_n3284), 
	.I(n3284));
   DELCKHD FE_PHC3206_n3848 (.O(FE_PHN3206_n3848), 
	.I(n3848));
   DELCKHD FE_PHC3205_n3592 (.O(FE_PHN3205_n3592), 
	.I(n3592));
   DELCKHD FE_PHC3204_n590 (.O(FE_PHN3204_n590), 
	.I(n590));
   DELCKHD FE_PHC3203_n3469 (.O(FE_PHN3203_n3469), 
	.I(n3469));
   DELDKHD FE_PHC3202_n4541 (.O(FE_PHN3202_n4541), 
	.I(n4541));
   DELDKHD FE_PHC3201_n1962 (.O(FE_PHN3201_n1962), 
	.I(n1962));
   DELDKHD FE_PHC3200_n2360 (.O(FE_PHN3200_n2360), 
	.I(n2360));
   DELDKHD FE_PHC3199_n2355 (.O(FE_PHN3199_n2355), 
	.I(n2355));
   DELDKHD FE_PHC3198_n1324 (.O(FE_PHN3198_n1324), 
	.I(n1324));
   DELDKHD FE_PHC3197_n3688 (.O(FE_PHN3197_n3688), 
	.I(n3688));
   DELDKHD FE_PHC3196_n1401 (.O(FE_PHN3196_n1401), 
	.I(n1401));
   DELCKHD FE_PHC3195_n706 (.O(FE_PHN3195_n706), 
	.I(n706));
   DELCKHD FE_PHC3194_n1328 (.O(FE_PHN3194_n1328), 
	.I(n1328));
   DELCKHD FE_PHC3193_n2012 (.O(FE_PHN3193_n2012), 
	.I(n2012));
   DELCKHD FE_PHC3192_n3846 (.O(FE_PHN3192_n3846), 
	.I(n3846));
   DELCKHD FE_PHC3191_n1511 (.O(FE_PHN3191_n1511), 
	.I(n1511));
   DELCKHD FE_PHC3190_n1978 (.O(FE_PHN3190_n1978), 
	.I(n1978));
   DELCKHD FE_PHC3189_n749 (.O(FE_PHN3189_n749), 
	.I(n749));
   DELCKHD FE_PHC3188_n1780 (.O(FE_PHN3188_n1780), 
	.I(n1780));
   DELCKHD FE_PHC3187_n1993 (.O(FE_PHN3187_n1993), 
	.I(n1993));
   DELCKHD FE_PHC3186_n3481 (.O(FE_PHN3186_n3481), 
	.I(n3481));
   DELCKHD FE_PHC3185_n1799 (.O(FE_PHN3185_n1799), 
	.I(n1799));
   DELCKHD FE_PHC3184_n1601 (.O(FE_PHN3184_n1601), 
	.I(n1601));
   DELCKHD FE_PHC3183_n3541 (.O(FE_PHN3183_n3541), 
	.I(n3541));
   DELCKHD FE_PHC3182_n1382 (.O(FE_PHN3182_n1382), 
	.I(n1382));
   DELCKHD FE_PHC3181_n2870 (.O(FE_PHN3181_n2870), 
	.I(n2870));
   DELCKHD FE_PHC3180_n592 (.O(FE_PHN3180_n592), 
	.I(n592));
   DELCKHD FE_PHC3179_n717 (.O(FE_PHN3179_n717), 
	.I(n717));
   DELCKHD FE_PHC3178_n1825 (.O(FE_PHN3178_n1825), 
	.I(n1825));
   DELCKHD FE_PHC3177_n4353 (.O(FE_PHN3177_n4353), 
	.I(n4353));
   DELDKHD FE_PHC3176_n832 (.O(FE_PHN3176_n832), 
	.I(n832));
   DELDKHD FE_PHC3175_n2505 (.O(FE_PHN3175_n2505), 
	.I(n2505));
   DELDKHD FE_PHC3174_n3843 (.O(FE_PHN3174_n3843), 
	.I(n3843));
   DELDKHD FE_PHC3173_n3519 (.O(FE_PHN3173_n3519), 
	.I(n3519));
   DELDKHD FE_PHC3172_n3388 (.O(FE_PHN3172_n3388), 
	.I(n3388));
   DELDKHD FE_PHC3171_n3769 (.O(FE_PHN3171_n3769), 
	.I(n3769));
   DELDKHD FE_PHC3170_n1279 (.O(FE_PHN3170_n1279), 
	.I(n1279));
   DELDKHD FE_PHC3169_n3483 (.O(FE_PHN3169_n3483), 
	.I(n3483));
   DELDKHD FE_PHC3168_n3471 (.O(FE_PHN3168_n3471), 
	.I(n3471));
   DELDKHD FE_PHC3167_n3280 (.O(FE_PHN3167_n3280), 
	.I(n3280));
   DELDKHD FE_PHC3166_n2511 (.O(FE_PHN3166_n2511), 
	.I(n2511));
   DELDKHD FE_PHC3165_n2196 (.O(FE_PHN3165_n2196), 
	.I(n2196));
   DELDKHD FE_PHC3164_n594 (.O(FE_PHN3164_n594), 
	.I(n594));
   DELDKHD FE_PHC3163_n2549 (.O(FE_PHN3163_n2549), 
	.I(n2549));
   DELDKHD FE_PHC3162_n4540 (.O(FE_PHN3162_n4540), 
	.I(n4540));
   DELDKHD FE_PHC3161_n2227 (.O(FE_PHN3161_n2227), 
	.I(n2227));
   DELDKHD FE_PHC3160_n1277 (.O(FE_PHN3160_n1277), 
	.I(n1277));
   DELDKHD FE_PHC3159_n1449 (.O(FE_PHN3159_n1449), 
	.I(n1449));
   DELCKHD FE_PHC3158_n801 (.O(FE_PHN3158_n801), 
	.I(n801));
   DELCKHD FE_PHC3157_n4096 (.O(FE_PHN3157_n4096), 
	.I(n4096));
   DELCKHD FE_PHC3156_n1405 (.O(FE_PHN3156_n1405), 
	.I(n1405));
   DELCKHD FE_PHC3155_n3891 (.O(FE_PHN3155_n3891), 
	.I(n3891));
   DELCKHD FE_PHC3154_n1772 (.O(FE_PHN3154_n1772), 
	.I(n1772));
   DELCKHD FE_PHC3153_n1699 (.O(FE_PHN3153_n1699), 
	.I(n1699));
   DELCKHD FE_PHC3152_n812 (.O(FE_PHN3152_n812), 
	.I(n812));
   DELCKHD FE_PHC3151_n1236 (.O(FE_PHN3151_n1236), 
	.I(n1236));
   DELCKHD FE_PHC3150_n651 (.O(FE_PHN3150_n651), 
	.I(n651));
   DELCKHD FE_PHC3149_n770 (.O(FE_PHN3149_n770), 
	.I(n770));
   DELCKHD FE_PHC3148_n1254 (.O(FE_PHN3148_n1254), 
	.I(n1254));
   DELCKHD FE_PHC3147_n2949 (.O(FE_PHN3147_n2949), 
	.I(n2949));
   DELCKHD FE_PHC3146_n3640 (.O(FE_PHN3146_n3640), 
	.I(n3640));
   DELCKHD FE_PHC3145_n1118 (.O(FE_PHN3145_n1118), 
	.I(n1118));
   DELCKHD FE_PHC3144_n1676 (.O(FE_PHN3144_n1676), 
	.I(n1676));
   DELCKHD FE_PHC3143_n1937 (.O(FE_PHN3143_n1937), 
	.I(n1937));
   DELCKHD FE_PHC3142_n1901 (.O(FE_PHN3142_n1901), 
	.I(n1901));
   DELCKHD FE_PHC3141_n1804 (.O(FE_PHN3141_n1804), 
	.I(n1804));
   DELCKHD FE_PHC3140_n1529 (.O(FE_PHN3140_n1529), 
	.I(n1529));
   DELCKHD FE_PHC3139_n3243 (.O(FE_PHN3139_n3243), 
	.I(n3243));
   DELCKHD FE_PHC3138_n1269 (.O(FE_PHN3138_n1269), 
	.I(n1269));
   DELCKHD FE_PHC3137_n758 (.O(FE_PHN3137_n758), 
	.I(n758));
   DELCKHD FE_PHC3136_n2358 (.O(FE_PHN3136_n2358), 
	.I(n2358));
   DELCKHD FE_PHC3135_n688 (.O(FE_PHN3135_n688), 
	.I(n688));
   DELCKHD FE_PHC3134_n3797 (.O(FE_PHN3134_n3797), 
	.I(n3797));
   DELCKHD FE_PHC3133_n715 (.O(FE_PHN3133_n715), 
	.I(n715));
   DELCKHD FE_PHC3132_n1354 (.O(FE_PHN3132_n1354), 
	.I(n1354));
   DELCKHD FE_PHC3131_n2446 (.O(FE_PHN3131_n2446), 
	.I(n2446));
   DELCKHD FE_PHC3130_n2223 (.O(FE_PHN3130_n2223), 
	.I(n2223));
   DELCKHD FE_PHC3129_n1203 (.O(FE_PHN3129_n1203), 
	.I(n1203));
   DELCKHD FE_PHC3128_n2700 (.O(FE_PHN3128_n2700), 
	.I(n2700));
   DELCKHD FE_PHC3127_n1043 (.O(FE_PHN3127_n1043), 
	.I(n1043));
   DELCKHD FE_PHC3126_n1737 (.O(FE_PHN3126_n1737), 
	.I(n1737));
   DELDKHD FE_PHC3125_n1593 (.O(FE_PHN3125_n1593), 
	.I(n1593));
   DELDKHD FE_PHC3124_n4557 (.O(FE_PHN3124_n4557), 
	.I(n4557));
   DELDKHD FE_PHC3123_n3777 (.O(FE_PHN3123_n3777), 
	.I(n3777));
   DELDKHD FE_PHC3122_n3220 (.O(FE_PHN3122_n3220), 
	.I(n3220));
   DELDKHD FE_PHC3121_n4173 (.O(FE_PHN3121_n4173), 
	.I(n4173));
   DELDKHD FE_PHC3120_n2613 (.O(FE_PHN3120_n2613), 
	.I(n2613));
   DELDKHD FE_PHC3119_n3784 (.O(FE_PHN3119_n3784), 
	.I(n3784));
   DELDKHD FE_PHC3118_n2868 (.O(FE_PHN3118_n2868), 
	.I(n2868));
   DELDKHD FE_PHC3117_n1714 (.O(FE_PHN3117_n1714), 
	.I(n1714));
   DELDKHD FE_PHC3116_n3143 (.O(FE_PHN3116_n3143), 
	.I(n3143));
   DELDKHD FE_PHC3115_n3697 (.O(FE_PHN3115_n3697), 
	.I(n3697));
   DELDKHD FE_PHC3114_n781 (.O(FE_PHN3114_n781), 
	.I(n781));
   DELDKHD FE_PHC3113_n1452 (.O(FE_PHN3113_n1452), 
	.I(n1452));
   DELDKHD FE_PHC3112_n2773 (.O(FE_PHN3112_n2773), 
	.I(n2773));
   DELDKHD FE_PHC3111_n1212 (.O(FE_PHN3111_n1212), 
	.I(n1212));
   DELDKHD FE_PHC3110_n2788 (.O(FE_PHN3110_n2788), 
	.I(n2788));
   DELDKHD FE_PHC3109_n1355 (.O(FE_PHN3109_n1355), 
	.I(n1355));
   DELDKHD FE_PHC3108_n3535 (.O(FE_PHN3108_n3535), 
	.I(n3535));
   DELDKHD FE_PHC3107_n3191 (.O(FE_PHN3107_n3191), 
	.I(n3191));
   DELDKHD FE_PHC3106_n1358 (.O(FE_PHN3106_n1358), 
	.I(n1358));
   DELDKHD FE_PHC3105_n1741 (.O(FE_PHN3105_n1741), 
	.I(n1741));
   DELDKHD FE_PHC3104_n2802 (.O(FE_PHN3104_n2802), 
	.I(n2802));
   DELDKHD FE_PHC3103_n1829 (.O(FE_PHN3103_n1829), 
	.I(n1829));
   DELDKHD FE_PHC3102_n2052 (.O(FE_PHN3102_n2052), 
	.I(n2052));
   DELDKHD FE_PHC3101_n2692 (.O(FE_PHN3101_n2692), 
	.I(n2692));
   DELDKHD FE_PHC3100_n2112 (.O(FE_PHN3100_n2112), 
	.I(n2112));
   DELDKHD FE_PHC3099_n2636 (.O(FE_PHN3099_n2636), 
	.I(n2636));
   DELDKHD FE_PHC3098_n1104 (.O(FE_PHN3098_n1104), 
	.I(n1104));
   DELDKHD FE_PHC3097_n1850 (.O(FE_PHN3097_n1850), 
	.I(n1850));
   DELDKHD FE_PHC3096_n1470 (.O(FE_PHN3096_n1470), 
	.I(n1470));
   DELDKHD FE_PHC3095_n3467 (.O(FE_PHN3095_n3467), 
	.I(n3467));
   DELDKHD FE_PHC3094_n3453 (.O(FE_PHN3094_n3453), 
	.I(n3453));
   DELCKHD FE_PHC3093_n1150 (.O(FE_PHN3093_n1150), 
	.I(n1150));
   DELCKHD FE_PHC3092_n3854 (.O(FE_PHN3092_n3854), 
	.I(n3854));
   DELCKHD FE_PHC3091_n2499 (.O(FE_PHN3091_n2499), 
	.I(n2499));
   DELCKHD FE_PHC3090_n3328 (.O(FE_PHN3090_n3328), 
	.I(n3328));
   DELCKHD FE_PHC3089_n3332 (.O(FE_PHN3089_n3332), 
	.I(n3332));
   DELCKHD FE_PHC3088_n907 (.O(FE_PHN3088_n907), 
	.I(n907));
   DELCKHD FE_PHC3087_n1935 (.O(FE_PHN3087_n1935), 
	.I(n1935));
   DELCKHD FE_PHC3086_n4043 (.O(FE_PHN3086_n4043), 
	.I(n4043));
   DELCKHD FE_PHC3085_n1731 (.O(FE_PHN3085_n1731), 
	.I(n1731));
   DELCKHD FE_PHC3084_n641 (.O(FE_PHN3084_n641), 
	.I(n641));
   DELCKHD FE_PHC3083_n1166 (.O(FE_PHN3083_n1166), 
	.I(n1166));
   DELCKHD FE_PHC3082_n3459 (.O(FE_PHN3082_n3459), 
	.I(n3459));
   DELCKHD FE_PHC3081_n2815 (.O(FE_PHN3081_n2815), 
	.I(n2815));
   DELCKHD FE_PHC3080_n1163 (.O(FE_PHN3080_n1163), 
	.I(n1163));
   DELCKHD FE_PHC3079_n4143 (.O(FE_PHN3079_n4143), 
	.I(n4143));
   DELCKHD FE_PHC3078_n1426 (.O(FE_PHN3078_n1426), 
	.I(n1426));
   DELCKHD FE_PHC3077_n1652 (.O(FE_PHN3077_n1652), 
	.I(n1652));
   DELCKHD FE_PHC3076_n1461 (.O(FE_PHN3076_n1461), 
	.I(n1461));
   DELCKHD FE_PHC3075_n1681 (.O(FE_PHN3075_n1681), 
	.I(n1681));
   DELCKHD FE_PHC3074_ram_143__10_ (.O(FE_PHN3074_ram_143__10_), 
	.I(\ram[143][10] ));
   DELCKHD FE_PHC3073_ram_52__15_ (.O(FE_PHN3073_ram_52__15_), 
	.I(\ram[52][15] ));
   DELCKHD FE_PHC3072_n3319 (.O(FE_PHN3072_n3319), 
	.I(n3319));
   DELCKHD FE_PHC3071_n2041 (.O(FE_PHN3071_n2041), 
	.I(n2041));
   DELCKHD FE_PHC3070_n1229 (.O(FE_PHN3070_n1229), 
	.I(n1229));
   DELCKHD FE_PHC3069_n2214 (.O(FE_PHN3069_n2214), 
	.I(n2214));
   DELCKHD FE_PHC3068_n4642 (.O(FE_PHN3068_n4642), 
	.I(n4642));
   DELCKHD FE_PHC3067_n1484 (.O(FE_PHN3067_n1484), 
	.I(n1484));
   DELCKHD FE_PHC3066_n811 (.O(FE_PHN3066_n811), 
	.I(n811));
   DELCKHD FE_PHC3065_n1101 (.O(FE_PHN3065_n1101), 
	.I(n1101));
   DELCKHD FE_PHC3064_n1161 (.O(FE_PHN3064_n1161), 
	.I(n1161));
   DELCKHD FE_PHC3063_n1349 (.O(FE_PHN3063_n1349), 
	.I(n1349));
   DELCKHD FE_PHC3062_n2304 (.O(FE_PHN3062_n2304), 
	.I(n2304));
   DELCKHD FE_PHC3061_n620 (.O(FE_PHN3061_n620), 
	.I(n620));
   DELCKHD FE_PHC3060_n1134 (.O(FE_PHN3060_n1134), 
	.I(n1134));
   DELCKHD FE_PHC3059_n1615 (.O(FE_PHN3059_n1615), 
	.I(n1615));
   DELCKHD FE_PHC3058_n1413 (.O(FE_PHN3058_n1413), 
	.I(n1413));
   DELCKHD FE_PHC3057_n3908 (.O(FE_PHN3057_n3908), 
	.I(n3908));
   DELCKHD FE_PHC3056_n3487 (.O(FE_PHN3056_n3487), 
	.I(n3487));
   DELCKHD FE_PHC3055_n1784 (.O(FE_PHN3055_n1784), 
	.I(n1784));
   DELCKHD FE_PHC3054_n1491 (.O(FE_PHN3054_n1491), 
	.I(n1491));
   DELCKHD FE_PHC3053_n2464 (.O(FE_PHN3053_n2464), 
	.I(n2464));
   DELCKHD FE_PHC3052_n596 (.O(FE_PHN3052_n596), 
	.I(n596));
   DELDKHD FE_PHC3051_n3634 (.O(FE_PHN3051_n3634), 
	.I(n3634));
   DELDKHD FE_PHC3050_n1111 (.O(FE_PHN3050_n1111), 
	.I(n1111));
   DELDKHD FE_PHC3049_n1376 (.O(FE_PHN3049_n1376), 
	.I(n1376));
   DELDKHD FE_PHC3048_n1543 (.O(FE_PHN3048_n1543), 
	.I(n1543));
   DELDKHD FE_PHC3047_n1600 (.O(FE_PHN3047_n1600), 
	.I(n1600));
   DELDKHD FE_PHC3046_n2053 (.O(FE_PHN3046_n2053), 
	.I(n2053));
   DELDKHD FE_PHC3045_n1574 (.O(FE_PHN3045_n1574), 
	.I(n1574));
   DELDKHD FE_PHC3044_n4662 (.O(FE_PHN3044_n4662), 
	.I(n4662));
   DELDKHD FE_PHC3043_n631 (.O(FE_PHN3043_n631), 
	.I(n631));
   DELDKHD FE_PHC3042_n1618 (.O(FE_PHN3042_n1618), 
	.I(n1618));
   DELDKHD FE_PHC3041_n1419 (.O(FE_PHN3041_n1419), 
	.I(n1419));
   DELDKHD FE_PHC3040_n3778 (.O(FE_PHN3040_n3778), 
	.I(n3778));
   DELDKHD FE_PHC3039_n1787 (.O(FE_PHN3039_n1787), 
	.I(n1787));
   DELDKHD FE_PHC3038_n1726 (.O(FE_PHN3038_n1726), 
	.I(n1726));
   DELDKHD FE_PHC3037_n585 (.O(FE_PHN3037_n585), 
	.I(n585));
   DELDKHD FE_PHC3036_n721 (.O(FE_PHN3036_n721), 
	.I(n721));
   DELDKHD FE_PHC3035_n2746 (.O(FE_PHN3035_n2746), 
	.I(n2746));
   DELDKHD FE_PHC3034_n828 (.O(FE_PHN3034_n828), 
	.I(n828));
   DELDKHD FE_PHC3033_n1757 (.O(FE_PHN3033_n1757), 
	.I(n1757));
   DELDKHD FE_PHC3032_n1259 (.O(FE_PHN3032_n1259), 
	.I(n1259));
   DELDKHD FE_PHC3031_n4510 (.O(FE_PHN3031_n4510), 
	.I(n4510));
   DELDKHD FE_PHC3030_n3462 (.O(FE_PHN3030_n3462), 
	.I(n3462));
   DELDKHD FE_PHC3029_n1613 (.O(FE_PHN3029_n1613), 
	.I(n1613));
   DELDKHD FE_PHC3028_n1301 (.O(FE_PHN3028_n1301), 
	.I(n1301));
   DELDKHD FE_PHC3027_n729 (.O(FE_PHN3027_n729), 
	.I(n729));
   DELDKHD FE_PHC3026_n2055 (.O(FE_PHN3026_n2055), 
	.I(n2055));
   DELDKHD FE_PHC3025_n3261 (.O(FE_PHN3025_n3261), 
	.I(n3261));
   DELDKHD FE_PHC3024_n2885 (.O(FE_PHN3024_n2885), 
	.I(n2885));
   DELDKHD FE_PHC3023_n1859 (.O(FE_PHN3023_n1859), 
	.I(n1859));
   DELDKHD FE_PHC3022_n1941 (.O(FE_PHN3022_n1941), 
	.I(n1941));
   DELDKHD FE_PHC3021_n4670 (.O(FE_PHN3021_n4670), 
	.I(n4670));
   DELDKHD FE_PHC3020_n2098 (.O(FE_PHN3020_n2098), 
	.I(n2098));
   DELDKHD FE_PHC3019_n1856 (.O(FE_PHN3019_n1856), 
	.I(n1856));
   DELDKHD FE_PHC3018_n2665 (.O(FE_PHN3018_n2665), 
	.I(n2665));
   DELDKHD FE_PHC3017_n1579 (.O(FE_PHN3017_n1579), 
	.I(n1579));
   DELDKHD FE_PHC3016_n2240 (.O(FE_PHN3016_n2240), 
	.I(n2240));
   DELDKHD FE_PHC3015_n2845 (.O(FE_PHN3015_n2845), 
	.I(n2845));
   DELDKHD FE_PHC3014_n1417 (.O(FE_PHN3014_n1417), 
	.I(n1417));
   DELDKHD FE_PHC3013_ram_244__10_ (.O(FE_PHN3013_ram_244__10_), 
	.I(\ram[244][10] ));
   DELDKHD FE_PHC3012_n2031 (.O(FE_PHN3012_n2031), 
	.I(n2031));
   DELDKHD FE_PHC3011_n616 (.O(FE_PHN3011_n616), 
	.I(n616));
   DELDKHD FE_PHC3010_n1361 (.O(FE_PHN3010_n1361), 
	.I(n1361));
   DELDKHD FE_PHC3009_n1540 (.O(FE_PHN3009_n1540), 
	.I(n1540));
   DELDKHD FE_PHC3008_n3443 (.O(FE_PHN3008_n3443), 
	.I(n3443));
   DELDKHD FE_PHC3007_n1289 (.O(FE_PHN3007_n1289), 
	.I(n1289));
   DELDKHD FE_PHC3006_n2051 (.O(FE_PHN3006_n2051), 
	.I(n2051));
   DELDKHD FE_PHC3005_n1451 (.O(FE_PHN3005_n1451), 
	.I(n1451));
   DELDKHD FE_PHC3004_n4542 (.O(FE_PHN3004_n4542), 
	.I(n4542));
   DELDKHD FE_PHC3003_n3466 (.O(FE_PHN3003_n3466), 
	.I(n3466));
   DELDKHD FE_PHC3002_n1969 (.O(FE_PHN3002_n1969), 
	.I(n1969));
   DELDKHD FE_PHC3001_n3639 (.O(FE_PHN3001_n3639), 
	.I(n3639));
   DELDKHD FE_PHC3000_n4304 (.O(FE_PHN3000_n4304), 
	.I(n4304));
   DELDKHD FE_PHC2999_n2804 (.O(FE_PHN2999_n2804), 
	.I(n2804));
   DELDKHD FE_PHC2998_n785 (.O(FE_PHN2998_n785), 
	.I(n785));
   DELDKHD FE_PHC2997_n1448 (.O(FE_PHN2997_n1448), 
	.I(n1448));
   DELDKHD FE_PHC2996_n3816 (.O(FE_PHN2996_n3816), 
	.I(n3816));
   DELCKHD FE_PHC2995_ram_250__1_ (.O(FE_PHN2995_ram_250__1_), 
	.I(\ram[250][1] ));
   DELCKHD FE_PHC2994_n1984 (.O(FE_PHN2994_n1984), 
	.I(n1984));
   DELCKHD FE_PHC2993_n1553 (.O(FE_PHN2993_n1553), 
	.I(n1553));
   DELCKHD FE_PHC2992_n4208 (.O(FE_PHN2992_n4208), 
	.I(n4208));
   DELCKHD FE_PHC2991_n1705 (.O(FE_PHN2991_n1705), 
	.I(n1705));
   DELCKHD FE_PHC2990_n4109 (.O(FE_PHN2990_n4109), 
	.I(n4109));
   DELCKHD FE_PHC2989_n2083 (.O(FE_PHN2989_n2083), 
	.I(n2083));
   DELCKHD FE_PHC2988_n2217 (.O(FE_PHN2988_n2217), 
	.I(n2217));
   DELCKHD FE_PHC2987_n1350 (.O(FE_PHN2987_n1350), 
	.I(n1350));
   DELCKHD FE_PHC2986_n1468 (.O(FE_PHN2986_n1468), 
	.I(n1468));
   DELCKHD FE_PHC2985_n2036 (.O(FE_PHN2985_n2036), 
	.I(n2036));
   DELCKHD FE_PHC2984_n583 (.O(FE_PHN2984_n583), 
	.I(n583));
   DELCKHD FE_PHC2983_n588 (.O(FE_PHN2983_n588), 
	.I(n588));
   DELCKHD FE_PHC2982_n1609 (.O(FE_PHN2982_n1609), 
	.I(n1609));
   DELCKHD FE_PHC2981_n1642 (.O(FE_PHN2981_n1642), 
	.I(n1642));
   DELCKHD FE_PHC2980_n2111 (.O(FE_PHN2980_n2111), 
	.I(n2111));
   DELCKHD FE_PHC2979_ram_46__2_ (.O(FE_PHN2979_ram_46__2_), 
	.I(\ram[46][2] ));
   DELCKHD FE_PHC2978_n4104 (.O(FE_PHN2978_n4104), 
	.I(n4104));
   DELCKHD FE_PHC2977_n3440 (.O(FE_PHN2977_n3440), 
	.I(n3440));
   DELCKHD FE_PHC2976_n2471 (.O(FE_PHN2976_n2471), 
	.I(n2471));
   DELCKHD FE_PHC2975_n699 (.O(FE_PHN2975_n699), 
	.I(n699));
   DELCKHD FE_PHC2974_n2506 (.O(FE_PHN2974_n2506), 
	.I(n2506));
   DELCKHD FE_PHC2973_n2030 (.O(FE_PHN2973_n2030), 
	.I(n2030));
   DELCKHD FE_PHC2972_n1897 (.O(FE_PHN2972_n1897), 
	.I(n1897));
   DELCKHD FE_PHC2971_n1103 (.O(FE_PHN2971_n1103), 
	.I(n1103));
   DELCKHD FE_PHC2970_n3714 (.O(FE_PHN2970_n3714), 
	.I(n3714));
   DELCKHD FE_PHC2969_n2105 (.O(FE_PHN2969_n2105), 
	.I(n2105));
   DELCKHD FE_PHC2968_n2445 (.O(FE_PHN2968_n2445), 
	.I(n2445));
   DELCKHD FE_PHC2967_n3503 (.O(FE_PHN2967_n3503), 
	.I(n3503));
   DELCKHD FE_PHC2966_n1164 (.O(FE_PHN2966_n1164), 
	.I(n1164));
   DELCKHD FE_PHC2965_n1336 (.O(FE_PHN2965_n1336), 
	.I(n1336));
   DELCKHD FE_PHC2964_n1914 (.O(FE_PHN2964_n1914), 
	.I(n1914));
   DELCKHD FE_PHC2963_n1963 (.O(FE_PHN2963_n1963), 
	.I(n1963));
   DELCKHD FE_PHC2962_n746 (.O(FE_PHN2962_n746), 
	.I(n746));
   DELCKHD FE_PHC2961_n3321 (.O(FE_PHN2961_n3321), 
	.I(n3321));
   DELCKHD FE_PHC2960_n2869 (.O(FE_PHN2960_n2869), 
	.I(n2869));
   DELCKHD FE_PHC2959_n3387 (.O(FE_PHN2959_n3387), 
	.I(n3387));
   DELCKHD FE_PHC2958_n1381 (.O(FE_PHN2958_n1381), 
	.I(n1381));
   DELCKHD FE_PHC2957_n1727 (.O(FE_PHN2957_n1727), 
	.I(n1727));
   DELCKHD FE_PHC2956_n1147 (.O(FE_PHN2956_n1147), 
	.I(n1147));
   DELCKHD FE_PHC2955_n2674 (.O(FE_PHN2955_n2674), 
	.I(n2674));
   DELCKHD FE_PHC2954_n2793 (.O(FE_PHN2954_n2793), 
	.I(n2793));
   DELCKHD FE_PHC2953_n1454 (.O(FE_PHN2953_n1454), 
	.I(n1454));
   DELCKHD FE_PHC2952_n2630 (.O(FE_PHN2952_n2630), 
	.I(n2630));
   DELCKHD FE_PHC2951_n655 (.O(FE_PHN2951_n655), 
	.I(n655));
   DELCKHD FE_PHC2950_n1325 (.O(FE_PHN2950_n1325), 
	.I(n1325));
   DELCKHD FE_PHC2949_n1750 (.O(FE_PHN2949_n1750), 
	.I(n1750));
   DELCKHD FE_PHC2948_n1725 (.O(FE_PHN2948_n1725), 
	.I(n1725));
   DELCKHD FE_PHC2947_n3392 (.O(FE_PHN2947_n3392), 
	.I(n3392));
   DELCKHD FE_PHC2946_n4497 (.O(FE_PHN2946_n4497), 
	.I(n4497));
   DELCKHD FE_PHC2945_n1271 (.O(FE_PHN2945_n1271), 
	.I(n1271));
   DELCKHD FE_PHC2944_n2060 (.O(FE_PHN2944_n2060), 
	.I(n2060));
   DELCKHD FE_PHC2943_ram_254__9_ (.O(FE_PHN2943_ram_254__9_), 
	.I(\ram[254][9] ));
   DELCKHD FE_PHC2942_n4667 (.O(FE_PHN2942_n4667), 
	.I(n4667));
   DELCKHD FE_PHC2941_n4141 (.O(FE_PHN2941_n4141), 
	.I(n4141));
   DELCKHD FE_PHC2940_n3635 (.O(FE_PHN2940_n3635), 
	.I(n3635));
   DELCKHD FE_PHC2939_n3540 (.O(FE_PHN2939_n3540), 
	.I(n3540));
   DELCKHD FE_PHC2938_n1281 (.O(FE_PHN2938_n1281), 
	.I(n1281));
   DELCKHD FE_PHC2937_n3447 (.O(FE_PHN2937_n3447), 
	.I(n3447));
   DELCKHD FE_PHC2936_n4093 (.O(FE_PHN2936_n4093), 
	.I(n4093));
   DELCKHD FE_PHC2935_n1213 (.O(FE_PHN2935_n1213), 
	.I(n1213));
   DELCKHD FE_PHC2934_n4538 (.O(FE_PHN2934_n4538), 
	.I(n4538));
   DELCKHD FE_PHC2933_n3786 (.O(FE_PHN2933_n3786), 
	.I(n3786));
   DELCKHD FE_PHC2932_n803 (.O(FE_PHN2932_n803), 
	.I(n803));
   DELCKHD FE_PHC2931_n613 (.O(FE_PHN2931_n613), 
	.I(n613));
   DELCKHD FE_PHC2930_n2306 (.O(FE_PHN2930_n2306), 
	.I(n2306));
   DELCKHD FE_PHC2929_n2546 (.O(FE_PHN2929_n2546), 
	.I(n2546));
   DELCKHD FE_PHC2928_n1455 (.O(FE_PHN2928_n1455), 
	.I(n1455));
   DELCKHD FE_PHC2927_n3826 (.O(FE_PHN2927_n3826), 
	.I(n3826));
   DELCKHD FE_PHC2926_n761 (.O(FE_PHN2926_n761), 
	.I(n761));
   DELCKHD FE_PHC2925_n1487 (.O(FE_PHN2925_n1487), 
	.I(n1487));
   DELCKHD FE_PHC2924_n1407 (.O(FE_PHN2924_n1407), 
	.I(n1407));
   DELCKHD FE_PHC2923_n2480 (.O(FE_PHN2923_n2480), 
	.I(n2480));
   DELCKHD FE_PHC2922_n2086 (.O(FE_PHN2922_n2086), 
	.I(n2086));
   DELCKHD FE_PHC2921_n3275 (.O(FE_PHN2921_n3275), 
	.I(n3275));
   DELDKHD FE_PHC2920_n2103 (.O(FE_PHN2920_n2103), 
	.I(n2103));
   DELDKHD FE_PHC2919_n3641 (.O(FE_PHN2919_n3641), 
	.I(n3641));
   DELDKHD FE_PHC2918_n1807 (.O(FE_PHN2918_n1807), 
	.I(n1807));
   DELDKHD FE_PHC2917_n3616 (.O(FE_PHN2917_n3616), 
	.I(n3616));
   DELDKHD FE_PHC2916_n3674 (.O(FE_PHN2916_n3674), 
	.I(n3674));
   DELDKHD FE_PHC2915_n3372 (.O(FE_PHN2915_n3372), 
	.I(n3372));
   DELDKHD FE_PHC2914_n691 (.O(FE_PHN2914_n691), 
	.I(n691));
   DELDKHD FE_PHC2913_n3370 (.O(FE_PHN2913_n3370), 
	.I(n3370));
   DELDKHD FE_PHC2912_n3598 (.O(FE_PHN2912_n3598), 
	.I(n3598));
   DELDKHD FE_PHC2911_n1752 (.O(FE_PHN2911_n1752), 
	.I(n1752));
   DELDKHD FE_PHC2910_n1779 (.O(FE_PHN2910_n1779), 
	.I(n1779));
   DELDKHD FE_PHC2909_n2048 (.O(FE_PHN2909_n2048), 
	.I(n2048));
   DELDKHD FE_PHC2908_n1977 (.O(FE_PHN2908_n1977), 
	.I(n1977));
   DELDKHD FE_PHC2907_n2320 (.O(FE_PHN2907_n2320), 
	.I(n2320));
   DELDKHD FE_PHC2906_n1917 (.O(FE_PHN2906_n1917), 
	.I(n1917));
   DELDKHD FE_PHC2905_n1266 (.O(FE_PHN2905_n1266), 
	.I(n1266));
   DELDKHD FE_PHC2904_n4462 (.O(FE_PHN2904_n4462), 
	.I(n4462));
   DELDKHD FE_PHC2903_n1533 (.O(FE_PHN2903_n1533), 
	.I(n1533));
   DELDKHD FE_PHC2902_n1225 (.O(FE_PHN2902_n1225), 
	.I(n1225));
   DELDKHD FE_PHC2901_n4606 (.O(FE_PHN2901_n4606), 
	.I(n4606));
   DELDKHD FE_PHC2900_n1205 (.O(FE_PHN2900_n1205), 
	.I(n1205));
   DELDKHD FE_PHC2899_n1488 (.O(FE_PHN2899_n1488), 
	.I(n1488));
   DELDKHD FE_PHC2898_n1748 (.O(FE_PHN2898_n1748), 
	.I(n1748));
   DELDKHD FE_PHC2897_n2247 (.O(FE_PHN2897_n2247), 
	.I(n2247));
   DELDKHD FE_PHC2896_n2565 (.O(FE_PHN2896_n2565), 
	.I(n2565));
   DELDKHD FE_PHC2895_n837 (.O(FE_PHN2895_n837), 
	.I(n837));
   DELDKHD FE_PHC2894_n3343 (.O(FE_PHN2894_n3343), 
	.I(n3343));
   DELDKHD FE_PHC2893_n2065 (.O(FE_PHN2893_n2065), 
	.I(n2065));
   DELDKHD FE_PHC2892_n1430 (.O(FE_PHN2892_n1430), 
	.I(n1430));
   DELDKHD FE_PHC2891_n702 (.O(FE_PHN2891_n702), 
	.I(n702));
   DELDKHD FE_PHC2890_n1806 (.O(FE_PHN2890_n1806), 
	.I(n1806));
   DELDKHD FE_PHC2889_n1133 (.O(FE_PHN2889_n1133), 
	.I(n1133));
   DELDKHD FE_PHC2888_n1309 (.O(FE_PHN2888_n1309), 
	.I(n1309));
   DELDKHD FE_PHC2887_n1545 (.O(FE_PHN2887_n1545), 
	.I(n1545));
   DELDKHD FE_PHC2886_n2001 (.O(FE_PHN2886_n2001), 
	.I(n2001));
   DELDKHD FE_PHC2885_n657 (.O(FE_PHN2885_n657), 
	.I(n657));
   DELDKHD FE_PHC2884_n4575 (.O(FE_PHN2884_n4575), 
	.I(n4575));
   DELDKHD FE_PHC2883_n2310 (.O(FE_PHN2883_n2310), 
	.I(n2310));
   DELDKHD FE_PHC2882_n1395 (.O(FE_PHN2882_n1395), 
	.I(n1395));
   DELDKHD FE_PHC2881_n1472 (.O(FE_PHN2881_n1472), 
	.I(n1472));
   DELDKHD FE_PHC2880_n643 (.O(FE_PHN2880_n643), 
	.I(n643));
   DELDKHD FE_PHC2879_n1107 (.O(FE_PHN2879_n1107), 
	.I(n1107));
   DELDKHD FE_PHC2878_n650 (.O(FE_PHN2878_n650), 
	.I(n650));
   DELDKHD FE_PHC2877_n2561 (.O(FE_PHN2877_n2561), 
	.I(n2561));
   DELDKHD FE_PHC2876_n2043 (.O(FE_PHN2876_n2043), 
	.I(n2043));
   DELDKHD FE_PHC2875_n2317 (.O(FE_PHN2875_n2317), 
	.I(n2317));
   DELDKHD FE_PHC2874_n2522 (.O(FE_PHN2874_n2522), 
	.I(n2522));
   DELDKHD FE_PHC2873_n4341 (.O(FE_PHN2873_n4341), 
	.I(n4341));
   DELDKHD FE_PHC2872_n1420 (.O(FE_PHN2872_n1420), 
	.I(n1420));
   DELDKHD FE_PHC2871_n633 (.O(FE_PHN2871_n633), 
	.I(n633));
   DELDKHD FE_PHC2870_n2370 (.O(FE_PHN2870_n2370), 
	.I(n2370));
   DELDKHD FE_PHC2869_n3426 (.O(FE_PHN2869_n3426), 
	.I(n3426));
   DELDKHD FE_PHC2868_n2078 (.O(FE_PHN2868_n2078), 
	.I(n2078));
   DELDKHD FE_PHC2867_n4216 (.O(FE_PHN2867_n4216), 
	.I(n4216));
   DELDKHD FE_PHC2866_n3626 (.O(FE_PHN2866_n3626), 
	.I(n3626));
   DELDKHD FE_PHC2865_n2093 (.O(FE_PHN2865_n2093), 
	.I(n2093));
   DELDKHD FE_PHC2864_n1280 (.O(FE_PHN2864_n1280), 
	.I(n1280));
   DELDKHD FE_PHC2863_n1117 (.O(FE_PHN2863_n1117), 
	.I(n1117));
   DELDKHD FE_PHC2862_n4460 (.O(FE_PHN2862_n4460), 
	.I(n4460));
   DELDKHD FE_PHC2861_n1083 (.O(FE_PHN2861_n1083), 
	.I(n1083));
   DELDKHD FE_PHC2860_n684 (.O(FE_PHN2860_n684), 
	.I(n684));
   DELDKHD FE_PHC2859_n1222 (.O(FE_PHN2859_n1222), 
	.I(n1222));
   DELDKHD FE_PHC2858_n1228 (.O(FE_PHN2858_n1228), 
	.I(n1228));
   DELDKHD FE_PHC2857_n2453 (.O(FE_PHN2857_n2453), 
	.I(n2453));
   DELDKHD FE_PHC2856_n3433 (.O(FE_PHN2856_n3433), 
	.I(n3433));
   DELDKHD FE_PHC2855_n3458 (.O(FE_PHN2855_n3458), 
	.I(n3458));
   DELDKHD FE_PHC2854_n1602 (.O(FE_PHN2854_n1602), 
	.I(n1602));
   DELDKHD FE_PHC2853_n3179 (.O(FE_PHN2853_n3179), 
	.I(n3179));
   DELDKHD FE_PHC2852_n1596 (.O(FE_PHN2852_n1596), 
	.I(n1596));
   DELDKHD FE_PHC2851_ram_78__8_ (.O(FE_PHN2851_ram_78__8_), 
	.I(\ram[78][8] ));
   DELDKHD FE_PHC2850_n2575 (.O(FE_PHN2850_n2575), 
	.I(n2575));
   DELDKHD FE_PHC2849_ram_104__13_ (.O(FE_PHN2849_ram_104__13_), 
	.I(\ram[104][13] ));
   DELDKHD FE_PHC2848_n658 (.O(FE_PHN2848_n658), 
	.I(n658));
   DELDKHD FE_PHC2847_n1848 (.O(FE_PHN2847_n1848), 
	.I(n1848));
   DELDKHD FE_PHC2846_n795 (.O(FE_PHN2846_n795), 
	.I(n795));
   DELDKHD FE_PHC2845_n754 (.O(FE_PHN2845_n754), 
	.I(n754));
   DELDKHD FE_PHC2844_n2756 (.O(FE_PHN2844_n2756), 
	.I(n2756));
   DELDKHD FE_PHC2843_n1457 (.O(FE_PHN2843_n1457), 
	.I(n1457));
   DELDKHD FE_PHC2842_n4098 (.O(FE_PHN2842_n4098), 
	.I(n4098));
   DELDKHD FE_PHC2841_n2215 (.O(FE_PHN2841_n2215), 
	.I(n2215));
   DELDKHD FE_PHC2840_n3830 (.O(FE_PHN2840_n3830), 
	.I(n3830));
   DELDKHD FE_PHC2839_n4430 (.O(FE_PHN2839_n4430), 
	.I(n4430));
   DELDKHD FE_PHC2838_n1759 (.O(FE_PHN2838_n1759), 
	.I(n1759));
   DELDKHD FE_PHC2837_n653 (.O(FE_PHN2837_n653), 
	.I(n653));
   DELDKHD FE_PHC2836_n645 (.O(FE_PHN2836_n645), 
	.I(n645));
   DELDKHD FE_PHC2835_n773 (.O(FE_PHN2835_n773), 
	.I(n773));
   DELDKHD FE_PHC2834_n3631 (.O(FE_PHN2834_n3631), 
	.I(n3631));
   DELDKHD FE_PHC2833_n1531 (.O(FE_PHN2833_n1531), 
	.I(n1531));
   DELDKHD FE_PHC2832_n3142 (.O(FE_PHN2832_n3142), 
	.I(n3142));
   DELDKHD FE_PHC2831_n2517 (.O(FE_PHN2831_n2517), 
	.I(n2517));
   DELDKHD FE_PHC2830_n1363 (.O(FE_PHN2830_n1363), 
	.I(n1363));
   DELDKHD FE_PHC2829_n623 (.O(FE_PHN2829_n623), 
	.I(n623));
   DELCKHD FE_PHC2828_ram_120__14_ (.O(FE_PHN2828_ram_120__14_), 
	.I(\ram[120][14] ));
   DELCKHD FE_PHC2827_n3475 (.O(FE_PHN2827_n3475), 
	.I(n3475));
   DELCKHD FE_PHC2826_n2675 (.O(FE_PHN2826_n2675), 
	.I(n2675));
   DELCKHD FE_PHC2825_n1290 (.O(FE_PHN2825_n1290), 
	.I(n1290));
   DELCKHD FE_PHC2824_n652 (.O(FE_PHN2824_n652), 
	.I(n652));
   DELCKHD FE_PHC2823_n2817 (.O(FE_PHN2823_n2817), 
	.I(n2817));
   DELCKHD FE_PHC2822_n3285 (.O(FE_PHN2822_n3285), 
	.I(n3285));
   DELCKHD FE_PHC2821_n719 (.O(FE_PHN2821_n719), 
	.I(n719));
   DELCKHD FE_PHC2820_n4464 (.O(FE_PHN2820_n4464), 
	.I(n4464));
   DELCKHD FE_PHC2819_n3518 (.O(FE_PHN2819_n3518), 
	.I(n3518));
   DELCKHD FE_PHC2818_n3669 (.O(FE_PHN2818_n3669), 
	.I(n3669));
   DELCKHD FE_PHC2817_n2766 (.O(FE_PHN2817_n2766), 
	.I(n2766));
   DELCKHD FE_PHC2816_n3896 (.O(FE_PHN2816_n3896), 
	.I(n3896));
   DELCKHD FE_PHC2815_n755 (.O(FE_PHN2815_n755), 
	.I(n755));
   DELCKHD FE_PHC2814_n1162 (.O(FE_PHN2814_n1162), 
	.I(n1162));
   DELCKHD FE_PHC2813_n1687 (.O(FE_PHN2813_n1687), 
	.I(n1687));
   DELCKHD FE_PHC2812_n1747 (.O(FE_PHN2812_n1747), 
	.I(n1747));
   DELCKHD FE_PHC2811_n629 (.O(FE_PHN2811_n629), 
	.I(n629));
   DELCKHD FE_PHC2810_n3320 (.O(FE_PHN2810_n3320), 
	.I(n3320));
   DELCKHD FE_PHC2809_n3455 (.O(FE_PHN2809_n3455), 
	.I(n3455));
   DELCKHD FE_PHC2808_n1476 (.O(FE_PHN2808_n1476), 
	.I(n1476));
   DELCKHD FE_PHC2807_n2116 (.O(FE_PHN2807_n2116), 
	.I(n2116));
   DELCKHD FE_PHC2806_n1961 (.O(FE_PHN2806_n1961), 
	.I(n1961));
   DELCKHD FE_PHC2805_n2109 (.O(FE_PHN2805_n2109), 
	.I(n2109));
   DELCKHD FE_PHC2804_n1293 (.O(FE_PHN2804_n1293), 
	.I(n1293));
   DELCKHD FE_PHC2803_n711 (.O(FE_PHN2803_n711), 
	.I(n711));
   DELCKHD FE_PHC2802_ram_45__11_ (.O(FE_PHN2802_ram_45__11_), 
	.I(\ram[45][11] ));
   DELCKHD FE_PHC2801_n2016 (.O(FE_PHN2801_n2016), 
	.I(n2016));
   DELCKHD FE_PHC2800_n4176 (.O(FE_PHN2800_n4176), 
	.I(n4176));
   DELCKHD FE_PHC2799_n1823 (.O(FE_PHN2799_n1823), 
	.I(n1823));
   DELCKHD FE_PHC2798_n2209 (.O(FE_PHN2798_n2209), 
	.I(n2209));
   DELCKHD FE_PHC2797_n710 (.O(FE_PHN2797_n710), 
	.I(n710));
   DELCKHD FE_PHC2796_n1569 (.O(FE_PHN2796_n1569), 
	.I(n1569));
   DELCKHD FE_PHC2795_n3860 (.O(FE_PHN2795_n3860), 
	.I(n3860));
   DELCKHD FE_PHC2794_n2050 (.O(FE_PHN2794_n2050), 
	.I(n2050));
   DELCKHD FE_PHC2793_n4305 (.O(FE_PHN2793_n4305), 
	.I(n4305));
   DELCKHD FE_PHC2792_n4547 (.O(FE_PHN2792_n4547), 
	.I(n4547));
   DELCKHD FE_PHC2791_n2479 (.O(FE_PHN2791_n2479), 
	.I(n2479));
   DELCKHD FE_PHC2790_n2210 (.O(FE_PHN2790_n2210), 
	.I(n2210));
   DELCKHD FE_PHC2789_n2769 (.O(FE_PHN2789_n2769), 
	.I(n2769));
   DELCKHD FE_PHC2788_n830 (.O(FE_PHN2788_n830), 
	.I(n830));
   DELCKHD FE_PHC2787_n3250 (.O(FE_PHN2787_n3250), 
	.I(n3250));
   DELCKHD FE_PHC2786_n1264 (.O(FE_PHN2786_n1264), 
	.I(n1264));
   DELCKHD FE_PHC2785_n1399 (.O(FE_PHN2785_n1399), 
	.I(n1399));
   DELCKHD FE_PHC2784_n1344 (.O(FE_PHN2784_n1344), 
	.I(n1344));
   DELCKHD FE_PHC2783_n3331 (.O(FE_PHN2783_n3331), 
	.I(n3331));
   DELCKHD FE_PHC2782_n1866 (.O(FE_PHN2782_n1866), 
	.I(n1866));
   DELCKHD FE_PHC2781_n1296 (.O(FE_PHN2781_n1296), 
	.I(n1296));
   DELCKHD FE_PHC2780_n1341 (.O(FE_PHN2780_n1341), 
	.I(n1341));
   DELCKHD FE_PHC2779_n4634 (.O(FE_PHN2779_n4634), 
	.I(n4634));
   DELCKHD FE_PHC2778_n3448 (.O(FE_PHN2778_n3448), 
	.I(n3448));
   DELCKHD FE_PHC2777_n2235 (.O(FE_PHN2777_n2235), 
	.I(n2235));
   DELCKHD FE_PHC2776_n1492 (.O(FE_PHN2776_n1492), 
	.I(n1492));
   DELCKHD FE_PHC2775_n3377 (.O(FE_PHN2775_n3377), 
	.I(n3377));
   DELCKHD FE_PHC2774_n2282 (.O(FE_PHN2774_n2282), 
	.I(n2282));
   DELCKHD FE_PHC2773_n1447 (.O(FE_PHN2773_n1447), 
	.I(n1447));
   DELCKHD FE_PHC2772_n3624 (.O(FE_PHN2772_n3624), 
	.I(n3624));
   DELCKHD FE_PHC2771_n1365 (.O(FE_PHN2771_n1365), 
	.I(n1365));
   DELCKHD FE_PHC2770_n3205 (.O(FE_PHN2770_n3205), 
	.I(n3205));
   DELCKHD FE_PHC2769_n4631 (.O(FE_PHN2769_n4631), 
	.I(n4631));
   DELCKHD FE_PHC2768_n1481 (.O(FE_PHN2768_n1481), 
	.I(n1481));
   DELCKHD FE_PHC2767_n1337 (.O(FE_PHN2767_n1337), 
	.I(n1337));
   DELCKHD FE_PHC2766_n2362 (.O(FE_PHN2766_n2362), 
	.I(n2362));
   DELCKHD FE_PHC2765_n1268 (.O(FE_PHN2765_n1268), 
	.I(n1268));
   DELCKHD FE_PHC2764_n2438 (.O(FE_PHN2764_n2438), 
	.I(n2438));
   DELCKHD FE_PHC2763_n1331 (.O(FE_PHN2763_n1331), 
	.I(n1331));
   DELCKHD FE_PHC2762_n3272 (.O(FE_PHN2762_n3272), 
	.I(n3272));
   DELCKHD FE_PHC2761_n3478 (.O(FE_PHN2761_n3478), 
	.I(n3478));
   DELCKHD FE_PHC2760_n2003 (.O(FE_PHN2760_n2003), 
	.I(n2003));
   DELCKHD FE_PHC2759_n3445 (.O(FE_PHN2759_n3445), 
	.I(n3445));
   DELCKHD FE_PHC2758_n2102 (.O(FE_PHN2758_n2102), 
	.I(n2102));
   DELCKHD FE_PHC2757_n1463 (.O(FE_PHN2757_n1463), 
	.I(n1463));
   DELCKHD FE_PHC2756_n1501 (.O(FE_PHN2756_n1501), 
	.I(n1501));
   DELCKHD FE_PHC2755_n1719 (.O(FE_PHN2755_n1719), 
	.I(n1719));
   DELCKHD FE_PHC2754_n2004 (.O(FE_PHN2754_n2004), 
	.I(n2004));
   DELCKHD FE_PHC2753_n2542 (.O(FE_PHN2753_n2542), 
	.I(n2542));
   DELCKHD FE_PHC2752_n1580 (.O(FE_PHN2752_n1580), 
	.I(n1580));
   DELCKHD FE_PHC2751_n2659 (.O(FE_PHN2751_n2659), 
	.I(n2659));
   DELCKHD FE_PHC2750_n819 (.O(FE_PHN2750_n819), 
	.I(n819));
   DELCKHD FE_PHC2749_n3668 (.O(FE_PHN2749_n3668), 
	.I(n3668));
   DELCKHD FE_PHC2748_n2723 (.O(FE_PHN2748_n2723), 
	.I(n2723));
   DELCKHD FE_PHC2747_n3665 (.O(FE_PHN2747_n3665), 
	.I(n3665));
   DELCKHD FE_PHC2746_n1940 (.O(FE_PHN2746_n1940), 
	.I(n1940));
   DELCKHD FE_PHC2745_n2037 (.O(FE_PHN2745_n2037), 
	.I(n2037));
   DELCKHD FE_PHC2744_n778 (.O(FE_PHN2744_n778), 
	.I(n778));
   DELCKHD FE_PHC2743_n2470 (.O(FE_PHN2743_n2470), 
	.I(n2470));
   DELCKHD FE_PHC2742_n3430 (.O(FE_PHN2742_n3430), 
	.I(n3430));
   DELCKHD FE_PHC2741_n2875 (.O(FE_PHN2741_n2875), 
	.I(n2875));
   DELCKHD FE_PHC2740_n2256 (.O(FE_PHN2740_n2256), 
	.I(n2256));
   DELCKHD FE_PHC2739_n1342 (.O(FE_PHN2739_n1342), 
	.I(n1342));
   DELCKHD FE_PHC2738_n2545 (.O(FE_PHN2738_n2545), 
	.I(n2545));
   DELCKHD FE_PHC2737_n2113 (.O(FE_PHN2737_n2113), 
	.I(n2113));
   DELCKHD FE_PHC2736_n2500 (.O(FE_PHN2736_n2500), 
	.I(n2500));
   DELCKHD FE_PHC2735_n1532 (.O(FE_PHN2735_n1532), 
	.I(n1532));
   DELCKHD FE_PHC2734_n3409 (.O(FE_PHN2734_n3409), 
	.I(n3409));
   DELCKHD FE_PHC2733_n1578 (.O(FE_PHN2733_n1578), 
	.I(n1578));
   DELDKHD FE_PHC2732_n1109 (.O(FE_PHN2732_n1109), 
	.I(n1109));
   DELDKHD FE_PHC2731_n2002 (.O(FE_PHN2731_n2002), 
	.I(n2002));
   DELDKHD FE_PHC2730_n814 (.O(FE_PHN2730_n814), 
	.I(n814));
   DELDKHD FE_PHC2729_n1127 (.O(FE_PHN2729_n1127), 
	.I(n1127));
   DELDKHD FE_PHC2728_n4330 (.O(FE_PHN2728_n4330), 
	.I(n4330));
   DELDKHD FE_PHC2727_n2326 (.O(FE_PHN2727_n2326), 
	.I(n2326));
   DELDKHD FE_PHC2726_n2066 (.O(FE_PHN2726_n2066), 
	.I(n2066));
   DELDKHD FE_PHC2725_n1789 (.O(FE_PHN2725_n1789), 
	.I(n1789));
   DELDKHD FE_PHC2724_n681 (.O(FE_PHN2724_n681), 
	.I(n681));
   DELDKHD FE_PHC2723_n2079 (.O(FE_PHN2723_n2079), 
	.I(n2079));
   DELDKHD FE_PHC2722_n799 (.O(FE_PHN2722_n799), 
	.I(n799));
   DELDKHD FE_PHC2721_n2757 (.O(FE_PHN2721_n2757), 
	.I(n2757));
   DELDKHD FE_PHC2720_n664 (.O(FE_PHN2720_n664), 
	.I(n664));
   DELDKHD FE_PHC2719_n937 (.O(FE_PHN2719_n937), 
	.I(n937));
   DELDKHD FE_PHC2718_n1200 (.O(FE_PHN2718_n1200), 
	.I(n1200));
   DELDKHD FE_PHC2717_n1097 (.O(FE_PHN2717_n1097), 
	.I(n1097));
   DELDKHD FE_PHC2716_n2368 (.O(FE_PHN2716_n2368), 
	.I(n2368));
   DELDKHD FE_PHC2715_n2351 (.O(FE_PHN2715_n2351), 
	.I(n2351));
   DELDKHD FE_PHC2714_n2367 (.O(FE_PHN2714_n2367), 
	.I(n2367));
   DELDKHD FE_PHC2713_n3738 (.O(FE_PHN2713_n3738), 
	.I(n3738));
   DELDKHD FE_PHC2712_n1739 (.O(FE_PHN2712_n1739), 
	.I(n1739));
   DELDKHD FE_PHC2711_n1467 (.O(FE_PHN2711_n1467), 
	.I(n1467));
   DELDKHD FE_PHC2710_n4480 (.O(FE_PHN2710_n4480), 
	.I(n4480));
   DELDKHD FE_PHC2709_n593 (.O(FE_PHN2709_n593), 
	.I(n593));
   DELDKHD FE_PHC2708_n2068 (.O(FE_PHN2708_n2068), 
	.I(n2068));
   DELDKHD FE_PHC2707_n1931 (.O(FE_PHN2707_n1931), 
	.I(n1931));
   DELDKHD FE_PHC2706_n2760 (.O(FE_PHN2706_n2760), 
	.I(n2760));
   DELDKHD FE_PHC2705_n1215 (.O(FE_PHN2705_n1215), 
	.I(n1215));
   DELDKHD FE_PHC2704_n2359 (.O(FE_PHN2704_n2359), 
	.I(n2359));
   DELDKHD FE_PHC2703_n3175 (.O(FE_PHN2703_n3175), 
	.I(n3175));
   DELDKHD FE_PHC2702_n2581 (.O(FE_PHN2702_n2581), 
	.I(n2581));
   DELDKHD FE_PHC2701_n2758 (.O(FE_PHN2701_n2758), 
	.I(n2758));
   DELDKHD FE_PHC2700_n3363 (.O(FE_PHN2700_n3363), 
	.I(n3363));
   DELDKHD FE_PHC2699_n2023 (.O(FE_PHN2699_n2023), 
	.I(n2023));
   DELDKHD FE_PHC2698_n1912 (.O(FE_PHN2698_n1912), 
	.I(n1912));
   DELDKHD FE_PHC2697_n2872 (.O(FE_PHN2697_n2872), 
	.I(n2872));
   DELDKHD FE_PHC2696_n2261 (.O(FE_PHN2696_n2261), 
	.I(n2261));
   DELDKHD FE_PHC2695_n4428 (.O(FE_PHN2695_n4428), 
	.I(n4428));
   DELDKHD FE_PHC2694_n2101 (.O(FE_PHN2694_n2101), 
	.I(n2101));
   DELDKHD FE_PHC2693_n1576 (.O(FE_PHN2693_n1576), 
	.I(n1576));
   DELDKHD FE_PHC2692_n2790 (.O(FE_PHN2692_n2790), 
	.I(n2790));
   DELDKHD FE_PHC2691_n1518 (.O(FE_PHN2691_n1518), 
	.I(n1518));
   DELDKHD FE_PHC2690_n2798 (.O(FE_PHN2690_n2798), 
	.I(n2798));
   DELDKHD FE_PHC2689_n2462 (.O(FE_PHN2689_n2462), 
	.I(n2462));
   DELDKHD FE_PHC2688_n1546 (.O(FE_PHN2688_n1546), 
	.I(n1546));
   DELDKHD FE_PHC2687_n3429 (.O(FE_PHN2687_n3429), 
	.I(n3429));
   DELDKHD FE_PHC2686_n2059 (.O(FE_PHN2686_n2059), 
	.I(n2059));
   DELDKHD FE_PHC2685_n1584 (.O(FE_PHN2685_n1584), 
	.I(n1584));
   DELDKHD FE_PHC2684_n1404 (.O(FE_PHN2684_n1404), 
	.I(n1404));
   DELDKHD FE_PHC2683_n2447 (.O(FE_PHN2683_n2447), 
	.I(n2447));
   DELDKHD FE_PHC2682_n1959 (.O(FE_PHN2682_n1959), 
	.I(n1959));
   DELDKHD FE_PHC2681_n1359 (.O(FE_PHN2681_n1359), 
	.I(n1359));
   DELDKHD FE_PHC2680_n3893 (.O(FE_PHN2680_n3893), 
	.I(n3893));
   DELDKHD FE_PHC2679_n584 (.O(FE_PHN2679_n584), 
	.I(n584));
   DELDKHD FE_PHC2678_n2248 (.O(FE_PHN2678_n2248), 
	.I(n2248));
   DELDKHD FE_PHC2677_n1774 (.O(FE_PHN2677_n1774), 
	.I(n1774));
   DELDKHD FE_PHC2676_n2038 (.O(FE_PHN2676_n2038), 
	.I(n2038));
   DELDKHD FE_PHC2675_n2759 (.O(FE_PHN2675_n2759), 
	.I(n2759));
   DELDKHD FE_PHC2674_n4047 (.O(FE_PHN2674_n4047), 
	.I(n4047));
   DELDKHD FE_PHC2673_n1868 (.O(FE_PHN2673_n1868), 
	.I(n1868));
   DELDKHD FE_PHC2672_n831 (.O(FE_PHN2672_n831), 
	.I(n831));
   DELDKHD FE_PHC2671_n1274 (.O(FE_PHN2671_n1274), 
	.I(n1274));
   DELDKHD FE_PHC2670_n2478 (.O(FE_PHN2670_n2478), 
	.I(n2478));
   DELDKHD FE_PHC2669_n1155 (.O(FE_PHN2669_n1155), 
	.I(n1155));
   DELDKHD FE_PHC2668_n2069 (.O(FE_PHN2668_n2069), 
	.I(n2069));
   DELDKHD FE_PHC2667_n1791 (.O(FE_PHN2667_n1791), 
	.I(n1791));
   DELDKHD FE_PHC2666_n1519 (.O(FE_PHN2666_n1519), 
	.I(n1519));
   DELDKHD FE_PHC2665_n2054 (.O(FE_PHN2665_n2054), 
	.I(n2054));
   DELDKHD FE_PHC2664_n1927 (.O(FE_PHN2664_n1927), 
	.I(n1927));
   DELDKHD FE_PHC2663_n3892 (.O(FE_PHN2663_n3892), 
	.I(n3892));
   DELDKHD FE_PHC2662_n3765 (.O(FE_PHN2662_n3765), 
	.I(n3765));
   DELDKHD FE_PHC2661_n1398 (.O(FE_PHN2661_n1398), 
	.I(n1398));
   DELDKHD FE_PHC2660_n2039 (.O(FE_PHN2660_n2039), 
	.I(n2039));
   DELDKHD FE_PHC2659_n2366 (.O(FE_PHN2659_n2366), 
	.I(n2366));
   DELDKHD FE_PHC2658_ram_33__9_ (.O(FE_PHN2658_ram_33__9_), 
	.I(\ram[33][9] ));
   DELDKHD FE_PHC2657_n3525 (.O(FE_PHN2657_n3525), 
	.I(n3525));
   DELDKHD FE_PHC2656_n2670 (.O(FE_PHN2656_n2670), 
	.I(n2670));
   DELDKHD FE_PHC2655_n2309 (.O(FE_PHN2655_n2309), 
	.I(n2309));
   DELDKHD FE_PHC2654_n731 (.O(FE_PHN2654_n731), 
	.I(n731));
   DELDKHD FE_PHC2653_n1924 (.O(FE_PHN2653_n1924), 
	.I(n1924));
   DELDKHD FE_PHC2652_n2241 (.O(FE_PHN2652_n2241), 
	.I(n2241));
   DELDKHD FE_PHC2651_n3394 (.O(FE_PHN2651_n3394), 
	.I(n3394));
   DELDKHD FE_PHC2650_n2242 (.O(FE_PHN2650_n2242), 
	.I(n2242));
   DELDKHD FE_PHC2649_n1555 (.O(FE_PHN2649_n1555), 
	.I(n1555));
   DELDKHD FE_PHC2648_n1672 (.O(FE_PHN2648_n1672), 
	.I(n1672));
   DELDKHD FE_PHC2647_n2629 (.O(FE_PHN2647_n2629), 
	.I(n2629));
   DELDKHD FE_PHC2646_n3792 (.O(FE_PHN2646_n3792), 
	.I(n3792));
   DELDKHD FE_PHC2645_n1148 (.O(FE_PHN2645_n1148), 
	.I(n1148));
   DELDKHD FE_PHC2644_n2560 (.O(FE_PHN2644_n2560), 
	.I(n2560));
   DELDKHD FE_PHC2643_n1744 (.O(FE_PHN2643_n1744), 
	.I(n1744));
   DELDKHD FE_PHC2642_n3376 (.O(FE_PHN2642_n3376), 
	.I(n3376));
   DELDKHD FE_PHC2641_n2642 (.O(FE_PHN2641_n2642), 
	.I(n2642));
   DELDKHD FE_PHC2640_n1278 (.O(FE_PHN2640_n1278), 
	.I(n1278));
   DELDKHD FE_PHC2639_n634 (.O(FE_PHN2639_n634), 
	.I(n634));
   DELDKHD FE_PHC2638_n4605 (.O(FE_PHN2638_n4605), 
	.I(n4605));
   DELDKHD FE_PHC2637_n1456 (.O(FE_PHN2637_n1456), 
	.I(n1456));
   DELDKHD FE_PHC2636_n1483 (.O(FE_PHN2636_n1483), 
	.I(n1483));
   DELDKHD FE_PHC2635_n1786 (.O(FE_PHN2635_n1786), 
	.I(n1786));
   DELDKHD FE_PHC2634_n916 (.O(FE_PHN2634_n916), 
	.I(n916));
   DELDKHD FE_PHC2633_n756 (.O(FE_PHN2633_n756), 
	.I(n756));
   DELDKHD FE_PHC2632_n2501 (.O(FE_PHN2632_n2501), 
	.I(n2501));
   DELDKHD FE_PHC2631_n3617 (.O(FE_PHN2631_n3617), 
	.I(n3617));
   DELDKHD FE_PHC2630_n3657 (.O(FE_PHN2630_n3657), 
	.I(n3657));
   DELDKHD FE_PHC2629_n2057 (.O(FE_PHN2629_n2057), 
	.I(n2057));
   DELDKHD FE_PHC2628_n1216 (.O(FE_PHN2628_n1216), 
	.I(n1216));
   DELDKHD FE_PHC2627_n3401 (.O(FE_PHN2627_n3401), 
	.I(n3401));
   DELDKHD FE_PHC2626_n1619 (.O(FE_PHN2626_n1619), 
	.I(n1619));
   DELDKHD FE_PHC2625_n2871 (.O(FE_PHN2625_n2871), 
	.I(n2871));
   DELDKHD FE_PHC2624_n1428 (.O(FE_PHN2624_n1428), 
	.I(n1428));
   DELDKHD FE_PHC2623_n4423 (.O(FE_PHN2623_n4423), 
	.I(n4423));
   DELDKHD FE_PHC2622_n4090 (.O(FE_PHN2622_n4090), 
	.I(n4090));
   DELDKHD FE_PHC2621_n2716 (.O(FE_PHN2621_n2716), 
	.I(n2716));
   DELDKHD FE_PHC2620_n1374 (.O(FE_PHN2620_n1374), 
	.I(n1374));
   DELDKHD FE_PHC2619_n2035 (.O(FE_PHN2619_n2035), 
	.I(n2035));
   DELDKHD FE_PHC2618_n2220 (.O(FE_PHN2618_n2220), 
	.I(n2220));
   DELDKHD FE_PHC2617_n1654 (.O(FE_PHN2617_n1654), 
	.I(n1654));
   DELDKHD FE_PHC2616_n3782 (.O(FE_PHN2616_n3782), 
	.I(n3782));
   DELDKHD FE_PHC2615_n742 (.O(FE_PHN2615_n742), 
	.I(n742));
   DELDKHD FE_PHC2614_n4205 (.O(FE_PHN2614_n4205), 
	.I(n4205));
   DELDKHD FE_PHC2613_n1875 (.O(FE_PHN2613_n1875), 
	.I(n1875));
   DELDKHD FE_PHC2612_n2281 (.O(FE_PHN2612_n2281), 
	.I(n2281));
   DELDKHD FE_PHC2611_n1436 (.O(FE_PHN2611_n1436), 
	.I(n1436));
   DELDKHD FE_PHC2610_n1263 (.O(FE_PHN2610_n1263), 
	.I(n1263));
   DELDKHD FE_PHC2609_n1767 (.O(FE_PHN2609_n1767), 
	.I(n1767));
   DELDKHD FE_PHC2608_n1421 (.O(FE_PHN2608_n1421), 
	.I(n1421));
   DELDKHD FE_PHC2607_n2115 (.O(FE_PHN2607_n2115), 
	.I(n2115));
   DELDKHD FE_PHC2606_n2708 (.O(FE_PHN2606_n2708), 
	.I(n2708));
   DELDKHD FE_PHC2605_n2008 (.O(FE_PHN2605_n2008), 
	.I(n2008));
   DELDKHD FE_PHC2604_n1153 (.O(FE_PHN2604_n1153), 
	.I(n1153));
   DELDKHD FE_PHC2603_n2882 (.O(FE_PHN2603_n2882), 
	.I(n2882));
   DELDKHD FE_PHC2602_n3567 (.O(FE_PHN2602_n3567), 
	.I(n3567));
   DELDKHD FE_PHC2601_n3856 (.O(FE_PHN2601_n3856), 
	.I(n3856));
   DELDKHD FE_PHC2600_n1938 (.O(FE_PHN2600_n1938), 
	.I(n1938));
   DELDKHD FE_PHC2599_n2117 (.O(FE_PHN2599_n2117), 
	.I(n2117));
   DELCKHD FE_PHC2598_ram_45__0_ (.O(FE_PHN2598_ram_45__0_), 
	.I(\ram[45][0] ));
   DELCKHD FE_PHC2597_ram_93__3_ (.O(FE_PHN2597_ram_93__3_), 
	.I(\ram[93][3] ));
   DELCKHD FE_PHC2596_n622 (.O(FE_PHN2596_n622), 
	.I(n622));
   DELCKHD FE_PHC2595_n1808 (.O(FE_PHN2595_n1808), 
	.I(n1808));
   DELCKHD FE_PHC2594_n1458 (.O(FE_PHN2594_n1458), 
	.I(n1458));
   DELCKHD FE_PHC2593_n1991 (.O(FE_PHN2593_n1991), 
	.I(n1991));
   DELCKHD FE_PHC2592_n766 (.O(FE_PHN2592_n766), 
	.I(n766));
   DELCKHD FE_PHC2591_n1950 (.O(FE_PHN2591_n1950), 
	.I(n1950));
   DELCKHD FE_PHC2590_n2224 (.O(FE_PHN2590_n2224), 
	.I(n2224));
   DELCKHD FE_PHC2589_n1135 (.O(FE_PHN2589_n1135), 
	.I(n1135));
   DELCKHD FE_PHC2588_n598 (.O(FE_PHN2588_n598), 
	.I(n598));
   DELCKHD FE_PHC2587_n3338 (.O(FE_PHN2587_n3338), 
	.I(n3338));
   DELCKHD FE_PHC2586_n1460 (.O(FE_PHN2586_n1460), 
	.I(n1460));
   DELCKHD FE_PHC2585_n3252 (.O(FE_PHN2585_n3252), 
	.I(n3252));
   DELCKHD FE_PHC2584_n3182 (.O(FE_PHN2584_n3182), 
	.I(n3182));
   DELCKHD FE_PHC2583_n1964 (.O(FE_PHN2583_n1964), 
	.I(n1964));
   DELCKHD FE_PHC2582_n3692 (.O(FE_PHN2582_n3692), 
	.I(n3692));
   DELCKHD FE_PHC2581_n3454 (.O(FE_PHN2581_n3454), 
	.I(n3454));
   DELCKHD FE_PHC2580_n3622 (.O(FE_PHN2580_n3622), 
	.I(n3622));
   DELCKHD FE_PHC2579_n3647 (.O(FE_PHN2579_n3647), 
	.I(n3647));
   DELCKHD FE_PHC2578_n2067 (.O(FE_PHN2578_n2067), 
	.I(n2067));
   DELCKHD FE_PHC2577_n1996 (.O(FE_PHN2577_n1996), 
	.I(n1996));
   DELCKHD FE_PHC2576_n3878 (.O(FE_PHN2576_n3878), 
	.I(n3878));
   DELCKHD FE_PHC2575_n2369 (.O(FE_PHN2575_n2369), 
	.I(n2369));
   DELCKHD FE_PHC2574_n1538 (.O(FE_PHN2574_n1538), 
	.I(n1538));
   DELCKHD FE_PHC2573_n782 (.O(FE_PHN2573_n782), 
	.I(n782));
   DELCKHD FE_PHC2572_n2544 (.O(FE_PHN2572_n2544), 
	.I(n2544));
   DELCKHD FE_PHC2571_n2535 (.O(FE_PHN2571_n2535), 
	.I(n2535));
   DELCKHD FE_PHC2570_n4050 (.O(FE_PHN2570_n4050), 
	.I(n4050));
   DELCKHD FE_PHC2569_n3689 (.O(FE_PHN2569_n3689), 
	.I(n3689));
   DELCKHD FE_PHC2568_n3235 (.O(FE_PHN2568_n3235), 
	.I(n3235));
   DELCKHD FE_PHC2567_n3302 (.O(FE_PHN2567_n3302), 
	.I(n3302));
   DELCKHD FE_PHC2566_n1287 (.O(FE_PHN2566_n1287), 
	.I(n1287));
   DELCKHD FE_PHC2565_n2504 (.O(FE_PHN2565_n2504), 
	.I(n2504));
   DELCKHD FE_PHC2564_n687 (.O(FE_PHN2564_n687), 
	.I(n687));
   DELCKHD FE_PHC2563_n1177 (.O(FE_PHN2563_n1177), 
	.I(n1177));
   DELCKHD FE_PHC2562_n3157 (.O(FE_PHN2562_n3157), 
	.I(n3157));
   DELCKHD FE_PHC2561_n3704 (.O(FE_PHN2561_n3704), 
	.I(n3704));
   DELCKHD FE_PHC2560_n4079 (.O(FE_PHN2560_n4079), 
	.I(n4079));
   DELCKHD FE_PHC2559_n1568 (.O(FE_PHN2559_n1568), 
	.I(n1568));
   DELCKHD FE_PHC2558_n4560 (.O(FE_PHN2558_n4560), 
	.I(n4560));
   DELCKHD FE_PHC2557_n1674 (.O(FE_PHN2557_n1674), 
	.I(n1674));
   DELCKHD FE_PHC2556_n3457 (.O(FE_PHN2556_n3457), 
	.I(n3457));
   DELCKHD FE_PHC2555_n2040 (.O(FE_PHN2555_n2040), 
	.I(n2040));
   DELCKHD FE_PHC2554_n1551 (.O(FE_PHN2554_n1551), 
	.I(n1551));
   DELCKHD FE_PHC2553_n1044 (.O(FE_PHN2553_n1044), 
	.I(n1044));
   DELCKHD FE_PHC2552_n1934 (.O(FE_PHN2552_n1934), 
	.I(n1934));
   DELCKHD FE_PHC2551_n1723 (.O(FE_PHN2551_n1723), 
	.I(n1723));
   DELCKHD FE_PHC2550_n3422 (.O(FE_PHN2550_n3422), 
	.I(n3422));
   DELCKHD FE_PHC2549_n1462 (.O(FE_PHN2549_n1462), 
	.I(n1462));
   DELCKHD FE_PHC2548_n3898 (.O(FE_PHN2548_n3898), 
	.I(n3898));
   DELCKHD FE_PHC2547_n1347 (.O(FE_PHN2547_n1347), 
	.I(n1347));
   DELCKHD FE_PHC2546_n1465 (.O(FE_PHN2546_n1465), 
	.I(n1465));
   DELCKHD FE_PHC2545_n4569 (.O(FE_PHN2545_n4569), 
	.I(n4569));
   DELCKHD FE_PHC2544_n4561 (.O(FE_PHN2544_n4561), 
	.I(n4561));
   DELCKHD FE_PHC2543_n3791 (.O(FE_PHN2543_n3791), 
	.I(n3791));
   DELCKHD FE_PHC2542_n2669 (.O(FE_PHN2542_n2669), 
	.I(n2669));
   DELCKHD FE_PHC2541_n3153 (.O(FE_PHN2541_n3153), 
	.I(n3153));
   DELCKHD FE_PHC2540_n2024 (.O(FE_PHN2540_n2024), 
	.I(n2024));
   DELCKHD FE_PHC2539_n2502 (.O(FE_PHN2539_n2502), 
	.I(n2502));
   DELCKHD FE_PHC2538_n3185 (.O(FE_PHN2538_n3185), 
	.I(n3185));
   DELCKHD FE_PHC2537_n3151 (.O(FE_PHN2537_n3151), 
	.I(n3151));
   DELCKHD FE_PHC2536_n3437 (.O(FE_PHN2536_n3437), 
	.I(n3437));
   DELCKHD FE_PHC2535_n3308 (.O(FE_PHN2535_n3308), 
	.I(n3308));
   DELCKHD FE_PHC2534_n2314 (.O(FE_PHN2534_n2314), 
	.I(n2314));
   DELCKHD FE_PHC2533_n2663 (.O(FE_PHN2533_n2663), 
	.I(n2663));
   DELCKHD FE_PHC2532_n4344 (.O(FE_PHN2532_n4344), 
	.I(n4344));
   DELCKHD FE_PHC2531_n939 (.O(FE_PHN2531_n939), 
	.I(n939));
   DELCKHD FE_PHC2530_n3524 (.O(FE_PHN2530_n3524), 
	.I(n3524));
   DELCKHD FE_PHC2529_n3795 (.O(FE_PHN2529_n3795), 
	.I(n3795));
   DELCKHD FE_PHC2528_n1156 (.O(FE_PHN2528_n1156), 
	.I(n1156));
   DELCKHD FE_PHC2527_n1474 (.O(FE_PHN2527_n1474), 
	.I(n1474));
   DELCKHD FE_PHC2526_n1242 (.O(FE_PHN2526_n1242), 
	.I(n1242));
   DELCKHD FE_PHC2525_n1343 (.O(FE_PHN2525_n1343), 
	.I(n1343));
   DELCKHD FE_PHC2524_n2487 (.O(FE_PHN2524_n2487), 
	.I(n2487));
   DELCKHD FE_PHC2523_n3522 (.O(FE_PHN2523_n3522), 
	.I(n3522));
   DELCKHD FE_PHC2522_n1513 (.O(FE_PHN2522_n1513), 
	.I(n1513));
   DELCKHD FE_PHC2521_n1438 (.O(FE_PHN2521_n1438), 
	.I(n1438));
   DELCKHD FE_PHC2520_n3504 (.O(FE_PHN2520_n3504), 
	.I(n3504));
   DELCKHD FE_PHC2519_n1283 (.O(FE_PHN2519_n1283), 
	.I(n1283));
   DELCKHD FE_PHC2518_n2184 (.O(FE_PHN2518_n2184), 
	.I(n2184));
   DELCKHD FE_PHC2517_n1389 (.O(FE_PHN2517_n1389), 
	.I(n1389));
   DELCKHD FE_PHC2516_n1662 (.O(FE_PHN2516_n1662), 
	.I(n1662));
   DELCKHD FE_PHC2515_n2280 (.O(FE_PHN2515_n2280), 
	.I(n2280));
   DELCKHD FE_PHC2514_n3259 (.O(FE_PHN2514_n3259), 
	.I(n3259));
   DELCKHD FE_PHC2513_n3654 (.O(FE_PHN2513_n3654), 
	.I(n3654));
   DELCKHD FE_PHC2512_n3756 (.O(FE_PHN2512_n3756), 
	.I(n3756));
   DELCKHD FE_PHC2511_n627 (.O(FE_PHN2511_n627), 
	.I(n627));
   DELCKHD FE_PHC2510_n2495 (.O(FE_PHN2510_n2495), 
	.I(n2495));
   DELCKHD FE_PHC2509_n1198 (.O(FE_PHN2509_n1198), 
	.I(n1198));
   DELCKHD FE_PHC2508_n1383 (.O(FE_PHN2508_n1383), 
	.I(n1383));
   DELCKHD FE_PHC2507_n1929 (.O(FE_PHN2507_n1929), 
	.I(n1929));
   DELCKHD FE_PHC2506_n2573 (.O(FE_PHN2506_n2573), 
	.I(n2573));
   DELCKHD FE_PHC2505_n1400 (.O(FE_PHN2505_n1400), 
	.I(n1400));
   DELCKHD FE_PHC2504_n1403 (.O(FE_PHN2504_n1403), 
	.I(n1403));
   DELCKHD FE_PHC2503_n3693 (.O(FE_PHN2503_n3693), 
	.I(n3693));
   DELCKHD FE_PHC2502_n3603 (.O(FE_PHN2502_n3603), 
	.I(n3603));
   DELCKHD FE_PHC2501_n1149 (.O(FE_PHN2501_n1149), 
	.I(n1149));
   DELCKHD FE_PHC2500_n1958 (.O(FE_PHN2500_n1958), 
	.I(n1958));
   DELCKHD FE_PHC2499_n1894 (.O(FE_PHN2499_n1894), 
	.I(n1894));
   DELCKHD FE_PHC2498_n2726 (.O(FE_PHN2498_n2726), 
	.I(n2726));
   DELCKHD FE_PHC2497_n2443 (.O(FE_PHN2497_n2443), 
	.I(n2443));
   DELCKHD FE_PHC2496_n1070 (.O(FE_PHN2496_n1070), 
	.I(n1070));
   DELCKHD FE_PHC2495_n2335 (.O(FE_PHN2495_n2335), 
	.I(n2335));
   DELCKHD FE_PHC2494_ram_45__14_ (.O(FE_PHN2494_ram_45__14_), 
	.I(\ram[45][14] ));
   DELCKHD FE_PHC2493_n1416 (.O(FE_PHN2493_n1416), 
	.I(n1416));
   DELCKHD FE_PHC2492_n2448 (.O(FE_PHN2492_n2448), 
	.I(n2448));
   DELCKHD FE_PHC2491_n1322 (.O(FE_PHN2491_n1322), 
	.I(n1322));
   DELCKHD FE_PHC2490_n2074 (.O(FE_PHN2490_n2074), 
	.I(n2074));
   DELCKHD FE_PHC2489_n1573 (.O(FE_PHN2489_n1573), 
	.I(n1573));
   DELCKHD FE_PHC2488_n3638 (.O(FE_PHN2488_n3638), 
	.I(n3638));
   DELCKHD FE_PHC2487_n3408 (.O(FE_PHN2487_n3408), 
	.I(n3408));
   DELCKHD FE_PHC2486_n1589 (.O(FE_PHN2486_n1589), 
	.I(n1589));
   DELCKHD FE_PHC2485_n2285 (.O(FE_PHN2485_n2285), 
	.I(n2285));
   DELCKHD FE_PHC2484_n3844 (.O(FE_PHN2484_n3844), 
	.I(n3844));
   DELCKHD FE_PHC2483_n3903 (.O(FE_PHN2483_n3903), 
	.I(n3903));
   DELCKHD FE_PHC2482_n1776 (.O(FE_PHN2482_n1776), 
	.I(n1776));
   DELCKHD FE_PHC2481_n1167 (.O(FE_PHN2481_n1167), 
	.I(n1167));
   DELCKHD FE_PHC2480_n2534 (.O(FE_PHN2480_n2534), 
	.I(n2534));
   DELCKHD FE_PHC2479_n3895 (.O(FE_PHN2479_n3895), 
	.I(n3895));
   DELCKHD FE_PHC2478_n642 (.O(FE_PHN2478_n642), 
	.I(n642));
   DELCKHD FE_PHC2477_n3523 (.O(FE_PHN2477_n3523), 
	.I(n3523));
   DELCKHD FE_PHC2476_n2631 (.O(FE_PHN2476_n2631), 
	.I(n2631));
   DELCKHD FE_PHC2475_n2483 (.O(FE_PHN2475_n2483), 
	.I(n2483));
   DELCKHD FE_PHC2474_n2863 (.O(FE_PHN2474_n2863), 
	.I(n2863));
   DELCKHD FE_PHC2473_n1219 (.O(FE_PHN2473_n1219), 
	.I(n1219));
   DELCKHD FE_PHC2472_n2693 (.O(FE_PHN2472_n2693), 
	.I(n2693));
   DELCKHD FE_PHC2471_n1992 (.O(FE_PHN2471_n1992), 
	.I(n1992));
   DELCKHD FE_PHC2470_n1171 (.O(FE_PHN2470_n1171), 
	.I(n1171));
   DELCKHD FE_PHC2469_n1464 (.O(FE_PHN2469_n1464), 
	.I(n1464));
   DELCKHD FE_PHC2468_n2510 (.O(FE_PHN2468_n2510), 
	.I(n2510));
   DELCKHD FE_PHC2467_n3722 (.O(FE_PHN2467_n3722), 
	.I(n3722));
   DELCKHD FE_PHC2466_n3432 (.O(FE_PHN2466_n3432), 
	.I(n3432));
   DELCKHD FE_PHC2465_n724 (.O(FE_PHN2465_n724), 
	.I(n724));
   DELCKHD FE_PHC2464_n4437 (.O(FE_PHN2464_n4437), 
	.I(n4437));
   DELCKHD FE_PHC2463_n3310 (.O(FE_PHN2463_n3310), 
	.I(n3310));
   DELCKHD FE_PHC2462_n1983 (.O(FE_PHN2462_n1983), 
	.I(n1983));
   DELCKHD FE_PHC2461_n1434 (.O(FE_PHN2461_n1434), 
	.I(n1434));
   DELCKHD FE_PHC2460_n2771 (.O(FE_PHN2460_n2771), 
	.I(n2771));
   DELCKHD FE_PHC2459_n2044 (.O(FE_PHN2459_n2044), 
	.I(n2044));
   DELCKHD FE_PHC2458_n2706 (.O(FE_PHN2458_n2706), 
	.I(n2706));
   DELCKHD FE_PHC2457_n3402 (.O(FE_PHN2457_n3402), 
	.I(n3402));
   DELCKHD FE_PHC2456_n1936 (.O(FE_PHN2456_n1936), 
	.I(n1936));
   DELDKHD FE_PHC2455_n3242 (.O(FE_PHN2455_n3242), 
	.I(n3242));
   DELDKHD FE_PHC2454_ram_81__1_ (.O(FE_PHN2454_ram_81__1_), 
	.I(\ram[81][1] ));
   DELDKHD FE_PHC2453_n692 (.O(FE_PHN2453_n692), 
	.I(n692));
   DELDKHD FE_PHC2452_n4128 (.O(FE_PHN2452_n4128), 
	.I(n4128));
   DELDKHD FE_PHC2451_n1345 (.O(FE_PHN2451_n1345), 
	.I(n1345));
   DELDKHD FE_PHC2450_n3818 (.O(FE_PHN2450_n3818), 
	.I(n3818));
   DELDKHD FE_PHC2449_n1469 (.O(FE_PHN2449_n1469), 
	.I(n1469));
   DELDKHD FE_PHC2448_n2820 (.O(FE_PHN2448_n2820), 
	.I(n2820));
   DELDKHD FE_PHC2447_n3507 (.O(FE_PHN2447_n3507), 
	.I(n3507));
   DELDKHD FE_PHC2446_n3144 (.O(FE_PHN2446_n3144), 
	.I(n3144));
   DELDKHD FE_PHC2445_n794 (.O(FE_PHN2445_n794), 
	.I(n794));
   DELDKHD FE_PHC2444_n3500 (.O(FE_PHN2444_n3500), 
	.I(n3500));
   DELDKHD FE_PHC2443_n3378 (.O(FE_PHN2443_n3378), 
	.I(n3378));
   DELDKHD FE_PHC2442_n2047 (.O(FE_PHN2442_n2047), 
	.I(n2047));
   DELDKHD FE_PHC2441_n1050 (.O(FE_PHN2441_n1050), 
	.I(n1050));
   DELDKHD FE_PHC2440_n3149 (.O(FE_PHN2440_n3149), 
	.I(n3149));
   DELDKHD FE_PHC2439_n2186 (.O(FE_PHN2439_n2186), 
	.I(n2186));
   DELDKHD FE_PHC2438_n3614 (.O(FE_PHN2438_n3614), 
	.I(n3614));
   DELDKHD FE_PHC2437_n1352 (.O(FE_PHN2437_n1352), 
	.I(n1352));
   DELDKHD FE_PHC2436_n1614 (.O(FE_PHN2436_n1614), 
	.I(n1614));
   DELDKHD FE_PHC2435_n4675 (.O(FE_PHN2435_n4675), 
	.I(n4675));
   DELDKHD FE_PHC2434_n1975 (.O(FE_PHN2434_n1975), 
	.I(n1975));
   DELDKHD FE_PHC2433_n2264 (.O(FE_PHN2433_n2264), 
	.I(n2264));
   DELDKHD FE_PHC2432_n4615 (.O(FE_PHN2432_n4615), 
	.I(n4615));
   DELDKHD FE_PHC2431_n1195 (.O(FE_PHN2431_n1195), 
	.I(n1195));
   DELDKHD FE_PHC2430_n700 (.O(FE_PHN2430_n700), 
	.I(n700));
   DELDKHD FE_PHC2429_n924 (.O(FE_PHN2429_n924), 
	.I(n924));
   DELDKHD FE_PHC2428_n2559 (.O(FE_PHN2428_n2559), 
	.I(n2559));
   DELDKHD FE_PHC2427_n1988 (.O(FE_PHN2427_n1988), 
	.I(n1988));
   DELDKHD FE_PHC2426_n2063 (.O(FE_PHN2426_n2063), 
	.I(n2063));
   DELDKHD FE_PHC2425_n2336 (.O(FE_PHN2425_n2336), 
	.I(n2336));
   DELDKHD FE_PHC2424_n3577 (.O(FE_PHN2424_n3577), 
	.I(n3577));
   DELDKHD FE_PHC2423_n1898 (.O(FE_PHN2423_n1898), 
	.I(n1898));
   DELDKHD FE_PHC2422_n1994 (.O(FE_PHN2422_n1994), 
	.I(n1994));
   DELDKHD FE_PHC2421_n3894 (.O(FE_PHN2421_n3894), 
	.I(n3894));
   DELDKHD FE_PHC2420_n1235 (.O(FE_PHN2420_n1235), 
	.I(n1235));
   DELDKHD FE_PHC2419_n639 (.O(FE_PHN2419_n639), 
	.I(n639));
   DELDKHD FE_PHC2418_n1267 (.O(FE_PHN2418_n1267), 
	.I(n1267));
   DELDKHD FE_PHC2417_n1486 (.O(FE_PHN2417_n1486), 
	.I(n1486));
   DELDKHD FE_PHC2416_n1734 (.O(FE_PHN2416_n1734), 
	.I(n1734));
   DELDKHD FE_PHC2415_n4539 (.O(FE_PHN2415_n4539), 
	.I(n4539));
   DELDKHD FE_PHC2414_n2795 (.O(FE_PHN2414_n2795), 
	.I(n2795));
   DELDKHD FE_PHC2413_n1883 (.O(FE_PHN2413_n1883), 
	.I(n1883));
   DELDKHD FE_PHC2412_n2555 (.O(FE_PHN2412_n2555), 
	.I(n2555));
   DELDKHD FE_PHC2411_n4614 (.O(FE_PHN2411_n4614), 
	.I(n4614));
   DELDKHD FE_PHC2410_n3649 (.O(FE_PHN2410_n3649), 
	.I(n3649));
   DELDKHD FE_PHC2409_n2022 (.O(FE_PHN2409_n2022), 
	.I(n2022));
   DELDKHD FE_PHC2408_n2562 (.O(FE_PHN2408_n2562), 
	.I(n2562));
   DELDKHD FE_PHC2407_n4645 (.O(FE_PHN2407_n4645), 
	.I(n4645));
   DELDKHD FE_PHC2406_n1115 (.O(FE_PHN2406_n1115), 
	.I(n1115));
   DELDKHD FE_PHC2405_n1284 (.O(FE_PHN2405_n1284), 
	.I(n1284));
   DELDKHD FE_PHC2404_n3683 (.O(FE_PHN2404_n3683), 
	.I(n3683));
   DELDKHD FE_PHC2403_n1693 (.O(FE_PHN2403_n1693), 
	.I(n1693));
   DELDKHD FE_PHC2402_n3630 (.O(FE_PHN2402_n3630), 
	.I(n3630));
   DELDKHD FE_PHC2401_n2543 (.O(FE_PHN2401_n2543), 
	.I(n2543));
   DELDKHD FE_PHC2400_n738 (.O(FE_PHN2400_n738), 
	.I(n738));
   DELDKHD FE_PHC2399_n1972 (.O(FE_PHN2399_n1972), 
	.I(n1972));
   DELDKHD FE_PHC2398_n3190 (.O(FE_PHN2398_n3190), 
	.I(n3190));
   DELDKHD FE_PHC2397_n3855 (.O(FE_PHN2397_n3855), 
	.I(n3855));
   DELDKHD FE_PHC2396_n638 (.O(FE_PHN2396_n638), 
	.I(n638));
   DELDKHD FE_PHC2395_n1778 (.O(FE_PHN2395_n1778), 
	.I(n1778));
   DELDKHD FE_PHC2394_n2344 (.O(FE_PHN2394_n2344), 
	.I(n2344));
   DELDKHD FE_PHC2393_n1665 (.O(FE_PHN2393_n1665), 
	.I(n1665));
   DELDKHD FE_PHC2392_n3417 (.O(FE_PHN2392_n3417), 
	.I(n3417));
   DELDKHD FE_PHC2391_n1157 (.O(FE_PHN2391_n1157), 
	.I(n1157));
   DELDKHD FE_PHC2390_n3341 (.O(FE_PHN2390_n3341), 
	.I(n3341));
   DELDKHD FE_PHC2389_n1997 (.O(FE_PHN2389_n1997), 
	.I(n1997));
   DELDKHD FE_PHC2388_n1257 (.O(FE_PHN2388_n1257), 
	.I(n1257));
   DELDKHD FE_PHC2387_n3656 (.O(FE_PHN2387_n3656), 
	.I(n3656));
   DELDKHD FE_PHC2386_n595 (.O(FE_PHN2386_n595), 
	.I(n595));
   DELDKHD FE_PHC2385_n834 (.O(FE_PHN2385_n834), 
	.I(n834));
   DELDKHD FE_PHC2384_n1356 (.O(FE_PHN2384_n1356), 
	.I(n1356));
   DELDKHD FE_PHC2383_n635 (.O(FE_PHN2383_n635), 
	.I(n635));
   DELDKHD FE_PHC2382_n777 (.O(FE_PHN2382_n777), 
	.I(n777));
   DELDKHD FE_PHC2381_n1857 (.O(FE_PHN2381_n1857), 
	.I(n1857));
   DELDKHD FE_PHC2380_n1671 (.O(FE_PHN2380_n1671), 
	.I(n1671));
   DELDKHD FE_PHC2379_n1437 (.O(FE_PHN2379_n1437), 
	.I(n1437));
   DELDKHD FE_PHC2378_n1876 (.O(FE_PHN2378_n1876), 
	.I(n1876));
   DELDKHD FE_PHC2377_n1987 (.O(FE_PHN2377_n1987), 
	.I(n1987));
   DELDKHD FE_PHC2376_n732 (.O(FE_PHN2376_n732), 
	.I(n732));
   DELDKHD FE_PHC2375_n3434 (.O(FE_PHN2375_n3434), 
	.I(n3434));
   DELDKHD FE_PHC2374_n2829 (.O(FE_PHN2374_n2829), 
	.I(n2829));
   DELDKHD FE_PHC2373_n2087 (.O(FE_PHN2373_n2087), 
	.I(n2087));
   DELDKHD FE_PHC2372_n1453 (.O(FE_PHN2372_n1453), 
	.I(n1453));
   DELDKHD FE_PHC2371_ram_241__0_ (.O(FE_PHN2371_ram_241__0_), 
	.I(\ram[241][0] ));
   DELDKHD FE_PHC2370_n4077 (.O(FE_PHN2370_n4077), 
	.I(n4077));
   DELDKHD FE_PHC2369_n1970 (.O(FE_PHN2369_n1970), 
	.I(n1970));
   DELDKHD FE_PHC2368_n2145 (.O(FE_PHN2368_n2145), 
	.I(n2145));
   DELDKHD FE_PHC2367_n2929 (.O(FE_PHN2367_n2929), 
	.I(n2929));
   DELDKHD FE_PHC2366_n4309 (.O(FE_PHN2366_n4309), 
	.I(n4309));
   DELDKHD FE_PHC2365_n4159 (.O(FE_PHN2365_n4159), 
	.I(n4159));
   DELDKHD FE_PHC2364_ram_9__1_ (.O(FE_PHN2364_ram_9__1_), 
	.I(\ram[9][1] ));
   DELDKHD FE_PHC2363_n3435 (.O(FE_PHN2363_n3435), 
	.I(n3435));
   DELDKHD FE_PHC2362_n3723 (.O(FE_PHN2362_n3723), 
	.I(n3723));
   DELDKHD FE_PHC2361_n1306 (.O(FE_PHN2361_n1306), 
	.I(n1306));
   DELDKHD FE_PHC2360_n2842 (.O(FE_PHN2360_n2842), 
	.I(n2842));
   DELDKHD FE_PHC2359_n1762 (.O(FE_PHN2359_n1762), 
	.I(n1762));
   DELDKHD FE_PHC2358_n2883 (.O(FE_PHN2358_n2883), 
	.I(n2883));
   DELDKHD FE_PHC2357_n1183 (.O(FE_PHN2357_n1183), 
	.I(n1183));
   DELDKHD FE_PHC2356_n3148 (.O(FE_PHN2356_n3148), 
	.I(n3148));
   DELDKHD FE_PHC2355_n4629 (.O(FE_PHN2355_n4629), 
	.I(n4629));
   DELDKHD FE_PHC2354_n2029 (.O(FE_PHN2354_n2029), 
	.I(n2029));
   DELDKHD FE_PHC2353_n789 (.O(FE_PHN2353_n789), 
	.I(n789));
   DELDKHD FE_PHC2352_n3374 (.O(FE_PHN2352_n3374), 
	.I(n3374));
   DELDKHD FE_PHC2351_n4549 (.O(FE_PHN2351_n4549), 
	.I(n4549));
   DELDKHD FE_PHC2350_n1587 (.O(FE_PHN2350_n1587), 
	.I(n1587));
   DELDKHD FE_PHC2349_n4596 (.O(FE_PHN2349_n4596), 
	.I(n4596));
   DELDKHD FE_PHC2348_n1974 (.O(FE_PHN2348_n1974), 
	.I(n1974));
   DELDKHD FE_PHC2347_n3351 (.O(FE_PHN2347_n3351), 
	.I(n3351));
   DELDKHD FE_PHC2346_n673 (.O(FE_PHN2346_n673), 
	.I(n673));
   DELDKHD FE_PHC2345_n1326 (.O(FE_PHN2345_n1326), 
	.I(n1326));
   DELDKHD FE_PHC2344_n1366 (.O(FE_PHN2344_n1366), 
	.I(n1366));
   DELDKHD FE_PHC2343_n3707 (.O(FE_PHN2343_n3707), 
	.I(n3707));
   DELDKHD FE_PHC2342_n1318 (.O(FE_PHN2342_n1318), 
	.I(n1318));
   DELDKHD FE_PHC2341_n4469 (.O(FE_PHN2341_n4469), 
	.I(n4469));
   DELDKHD FE_PHC2340_n1530 (.O(FE_PHN2340_n1530), 
	.I(n1530));
   DELDKHD FE_PHC2339_n2049 (.O(FE_PHN2339_n2049), 
	.I(n2049));
   DELDKHD FE_PHC2338_n2090 (.O(FE_PHN2338_n2090), 
	.I(n2090));
   DELDKHD FE_PHC2337_n3750 (.O(FE_PHN2337_n3750), 
	.I(n3750));
   DELDKHD FE_PHC2336_n1256 (.O(FE_PHN2336_n1256), 
	.I(n1256));
   DELDKHD FE_PHC2335_n1946 (.O(FE_PHN2335_n1946), 
	.I(n1946));
   DELDKHD FE_PHC2334_n4073 (.O(FE_PHN2334_n4073), 
	.I(n4073));
   DELDKHD FE_PHC2333_n2021 (.O(FE_PHN2333_n2021), 
	.I(n2021));
   DELDKHD FE_PHC2332_n2569 (.O(FE_PHN2332_n2569), 
	.I(n2569));
   DELDKHD FE_PHC2331_n4482 (.O(FE_PHN2331_n4482), 
	.I(n4482));
   DELDKHD FE_PHC2330_n1427 (.O(FE_PHN2330_n1427), 
	.I(n1427));
   DELDKHD FE_PHC2329_n3456 (.O(FE_PHN2329_n3456), 
	.I(n3456));
   DELDKHD FE_PHC2328_n3849 (.O(FE_PHN2328_n3849), 
	.I(n3849));
   DELDKHD FE_PHC2327_n1311 (.O(FE_PHN2327_n1311), 
	.I(n1311));
   DELCKHD FE_PHC2326_ram_67__9_ (.O(FE_PHN2326_ram_67__9_), 
	.I(\ram[67][9] ));
   DELCKHD FE_PHC2325_n646 (.O(FE_PHN2325_n646), 
	.I(n646));
   DELCKHD FE_PHC2324_n4544 (.O(FE_PHN2324_n4544), 
	.I(n4544));
   DELCKHD FE_PHC2323_n3298 (.O(FE_PHN2323_n3298), 
	.I(n3298));
   DELCKHD FE_PHC2322_n3776 (.O(FE_PHN2322_n3776), 
	.I(n3776));
   DELCKHD FE_PHC2321_n4312 (.O(FE_PHN2321_n4312), 
	.I(n4312));
   DELCKHD FE_PHC2320_n2672 (.O(FE_PHN2320_n2672), 
	.I(n2672));
   DELCKHD FE_PHC2319_n2550 (.O(FE_PHN2319_n2550), 
	.I(n2550));
   DELCKHD FE_PHC2318_n3476 (.O(FE_PHN2318_n3476), 
	.I(n3476));
   DELCKHD FE_PHC2317_n4620 (.O(FE_PHN2317_n4620), 
	.I(n4620));
   DELCKHD FE_PHC2316_n4513 (.O(FE_PHN2316_n4513), 
	.I(n4513));
   DELCKHD FE_PHC2315_n2541 (.O(FE_PHN2315_n2541), 
	.I(n2541));
   DELCKHD FE_PHC2314_n1243 (.O(FE_PHN2314_n1243), 
	.I(n1243));
   DELCKHD FE_PHC2313_n940 (.O(FE_PHN2313_n940), 
	.I(n940));
   DELCKHD FE_PHC2312_n685 (.O(FE_PHN2312_n685), 
	.I(n685));
   DELCKHD FE_PHC2311_n1272 (.O(FE_PHN2311_n1272), 
	.I(n1272));
   DELCKHD FE_PHC2310_n3659 (.O(FE_PHN2310_n3659), 
	.I(n3659));
   DELCKHD FE_PHC2309_n3858 (.O(FE_PHN2309_n3858), 
	.I(n3858));
   DELCKHD FE_PHC2308_n4457 (.O(FE_PHN2308_n4457), 
	.I(n4457));
   DELCKHD FE_PHC2307_n4597 (.O(FE_PHN2307_n4597), 
	.I(n4597));
   DELCKHD FE_PHC2306_n2302 (.O(FE_PHN2306_n2302), 
	.I(n2302));
   DELCKHD FE_PHC2305_n2234 (.O(FE_PHN2305_n2234), 
	.I(n2234));
   DELCKHD FE_PHC2304_n955 (.O(FE_PHN2304_n955), 
	.I(n955));
   DELCKHD FE_PHC2303_n4345 (.O(FE_PHN2303_n4345), 
	.I(n4345));
   DELCKHD FE_PHC2302_n3203 (.O(FE_PHN2302_n3203), 
	.I(n3203));
   DELCKHD FE_PHC2301_n1303 (.O(FE_PHN2301_n1303), 
	.I(n1303));
   DELCKHD FE_PHC2300_n2662 (.O(FE_PHN2300_n2662), 
	.I(n2662));
   DELCKHD FE_PHC2299_n4144 (.O(FE_PHN2299_n4144), 
	.I(n4144));
   DELCKHD FE_PHC2298_n1796 (.O(FE_PHN2298_n1796), 
	.I(n1796));
   DELCKHD FE_PHC2297_n2639 (.O(FE_PHN2297_n2639), 
	.I(n2639));
   DELCKHD FE_PHC2296_n3506 (.O(FE_PHN2296_n3506), 
	.I(n3506));
   DELCKHD FE_PHC2295_n1512 (.O(FE_PHN2295_n1512), 
	.I(n1512));
   DELCKHD FE_PHC2294_n3812 (.O(FE_PHN2294_n3812), 
	.I(n3812));
   DELCKHD FE_PHC2293_n3400 (.O(FE_PHN2293_n3400), 
	.I(n3400));
   DELCKHD FE_PHC2292_n1591 (.O(FE_PHN2292_n1591), 
	.I(n1591));
   DELCKHD FE_PHC2291_n1592 (.O(FE_PHN2291_n1592), 
	.I(n1592));
   DELCKHD FE_PHC2290_n3897 (.O(FE_PHN2290_n3897), 
	.I(n3897));
   DELCKHD FE_PHC2289_n1441 (.O(FE_PHN2289_n1441), 
	.I(n1441));
   DELCKHD FE_PHC2288_ram_45__8_ (.O(FE_PHN2288_ram_45__8_), 
	.I(\ram[45][8] ));
   DELCKHD FE_PHC2287_n2824 (.O(FE_PHN2287_n2824), 
	.I(n2824));
   DELCKHD FE_PHC2286_ram_217__3_ (.O(FE_PHN2286_ram_217__3_), 
	.I(\ram[217][3] ));
   DELCKHD FE_PHC2285_n3731 (.O(FE_PHN2285_n3731), 
	.I(n3731));
   DELCKHD FE_PHC2284_n632 (.O(FE_PHN2284_n632), 
	.I(n632));
   DELCKHD FE_PHC2283_n1520 (.O(FE_PHN2283_n1520), 
	.I(n1520));
   DELCKHD FE_PHC2282_n1208 (.O(FE_PHN2282_n1208), 
	.I(n1208));
   DELCKHD FE_PHC2281_n2865 (.O(FE_PHN2281_n2865), 
	.I(n2865));
   DELCKHD FE_PHC2280_n4075 (.O(FE_PHN2280_n4075), 
	.I(n4075));
   DELCKHD FE_PHC2279_n1294 (.O(FE_PHN2279_n1294), 
	.I(n1294));
   DELCKHD FE_PHC2278_n739 (.O(FE_PHN2278_n739), 
	.I(n739));
   DELCKHD FE_PHC2277_n1223 (.O(FE_PHN2277_n1223), 
	.I(n1223));
   DELCKHD FE_PHC2276_n3840 (.O(FE_PHN2276_n3840), 
	.I(n3840));
   DELCKHD FE_PHC2275_n3413 (.O(FE_PHN2275_n3413), 
	.I(n3413));
   DELCKHD FE_PHC2274_n3701 (.O(FE_PHN2274_n3701), 
	.I(n3701));
   DELCKHD FE_PHC2273_n2339 (.O(FE_PHN2273_n2339), 
	.I(n2339));
   DELCKHD FE_PHC2272_n1598 (.O(FE_PHN2272_n1598), 
	.I(n1598));
   DELCKHD FE_PHC2271_n1788 (.O(FE_PHN2271_n1788), 
	.I(n1788));
   DELCKHD FE_PHC2270_n1684 (.O(FE_PHN2270_n1684), 
	.I(n1684));
   DELCKHD FE_PHC2269_n2607 (.O(FE_PHN2269_n2607), 
	.I(n2607));
   DELCKHD FE_PHC2268_n3779 (.O(FE_PHN2268_n3779), 
	.I(n3779));
   DELCKHD FE_PHC2267_n4149 (.O(FE_PHN2267_n4149), 
	.I(n4149));
   DELCKHD FE_PHC2266_n705 (.O(FE_PHN2266_n705), 
	.I(n705));
   DELCKHD FE_PHC2265_n2100 (.O(FE_PHN2265_n2100), 
	.I(n2100));
   DELCKHD FE_PHC2264_n1096 (.O(FE_PHN2264_n1096), 
	.I(n1096));
   DELCKHD FE_PHC2263_n4301 (.O(FE_PHN2263_n4301), 
	.I(n4301));
   DELCKHD FE_PHC2262_n677 (.O(FE_PHN2262_n677), 
	.I(n677));
   DELCKHD FE_PHC2261_n1638 (.O(FE_PHN2261_n1638), 
	.I(n1638));
   DELCKHD FE_PHC2260_n744 (.O(FE_PHN2260_n744), 
	.I(n744));
   DELCKHD FE_PHC2259_n1482 (.O(FE_PHN2259_n1482), 
	.I(n1482));
   DELCKHD FE_PHC2258_n1315 (.O(FE_PHN2258_n1315), 
	.I(n1315));
   DELCKHD FE_PHC2257_n3186 (.O(FE_PHN2257_n3186), 
	.I(n3186));
   DELCKHD FE_PHC2256_n1201 (.O(FE_PHN2256_n1201), 
	.I(n1201));
   DELCKHD FE_PHC2255_n701 (.O(FE_PHN2255_n701), 
	.I(n701));
   DELCKHD FE_PHC2254_n1224 (.O(FE_PHN2254_n1224), 
	.I(n1224));
   DELCKHD FE_PHC2253_n589 (.O(FE_PHN2253_n589), 
	.I(n589));
   DELCKHD FE_PHC2252_n2755 (.O(FE_PHN2252_n2755), 
	.I(n2755));
   DELCKHD FE_PHC2251_n1221 (.O(FE_PHN2251_n1221), 
	.I(n1221));
   DELCKHD FE_PHC2250_n1262 (.O(FE_PHN2250_n1262), 
	.I(n1262));
   DELCKHD FE_PHC2249_n1517 (.O(FE_PHN2249_n1517), 
	.I(n1517));
   DELCKHD FE_PHC2248_n3686 (.O(FE_PHN2248_n3686), 
	.I(n3686));
   DELCKHD FE_PHC2247_n2813 (.O(FE_PHN2247_n2813), 
	.I(n2813));
   DELCKHD FE_PHC2246_n1660 (.O(FE_PHN2246_n1660), 
	.I(n1660));
   DELCKHD FE_PHC2245_n1926 (.O(FE_PHN2245_n1926), 
	.I(n1926));
   DELCKHD FE_PHC2244_n1362 (.O(FE_PHN2244_n1362), 
	.I(n1362));
   DELCKHD FE_PHC2243_n586 (.O(FE_PHN2243_n586), 
	.I(n586));
   DELCKHD FE_PHC2242_n760 (.O(FE_PHN2242_n760), 
	.I(n760));
   DELCKHD FE_PHC2241_n829 (.O(FE_PHN2241_n829), 
	.I(n829));
   DELCKHD FE_PHC2240_n2528 (.O(FE_PHN2240_n2528), 
	.I(n2528));
   DELCKHD FE_PHC2239_n2867 (.O(FE_PHN2239_n2867), 
	.I(n2867));
   DELCKHD FE_PHC2238_n4536 (.O(FE_PHN2238_n4536), 
	.I(n4536));
   DELCKHD FE_PHC2237_n1120 (.O(FE_PHN2237_n1120), 
	.I(n1120));
   DELCKHD FE_PHC2236_n2203 (.O(FE_PHN2236_n2203), 
	.I(n2203));
   DELCKHD FE_PHC2235_n2232 (.O(FE_PHN2235_n2232), 
	.I(n2232));
   DELCKHD FE_PHC2234_n4100 (.O(FE_PHN2234_n4100), 
	.I(n4100));
   DELCKHD FE_PHC2233_n3751 (.O(FE_PHN2233_n3751), 
	.I(n3751));
   DELCKHD FE_PHC2232_n604 (.O(FE_PHN2232_n604), 
	.I(n604));
   DELCKHD FE_PHC2231_n2009 (.O(FE_PHN2231_n2009), 
	.I(n2009));
   DELCKHD FE_PHC2230_n2485 (.O(FE_PHN2230_n2485), 
	.I(n2485));
   DELCKHD FE_PHC2229_n752 (.O(FE_PHN2229_n752), 
	.I(n752));
   DELCKHD FE_PHC2228_n2091 (.O(FE_PHN2228_n2091), 
	.I(n2091));
   DELCKHD FE_PHC2227_n3237 (.O(FE_PHN2227_n3237), 
	.I(n3237));
   DELCKHD FE_PHC2226_n1357 (.O(FE_PHN2226_n1357), 
	.I(n1357));
   DELCKHD FE_PHC2225_n747 (.O(FE_PHN2225_n747), 
	.I(n747));
   DELCKHD FE_PHC2224_n2861 (.O(FE_PHN2224_n2861), 
	.I(n2861));
   DELCKHD FE_PHC2223_n716 (.O(FE_PHN2223_n716), 
	.I(n716));
   DELCKHD FE_PHC2222_n2061 (.O(FE_PHN2222_n2061), 
	.I(n2061));
   DELCKHD FE_PHC2221_n3889 (.O(FE_PHN2221_n3889), 
	.I(n3889));
   DELCKHD FE_PHC2220_n1677 (.O(FE_PHN2220_n1677), 
	.I(n1677));
   DELCKHD FE_PHC2219_n1036 (.O(FE_PHN2219_n1036), 
	.I(n1036));
   DELCKHD FE_PHC2218_n1968 (.O(FE_PHN2218_n1968), 
	.I(n1968));
   DELCKHD FE_PHC2217_n2322 (.O(FE_PHN2217_n2322), 
	.I(n2322));
   DELCKHD FE_PHC2216_n4621 (.O(FE_PHN2216_n4621), 
	.I(n4621));
   DELCKHD FE_PHC2215_n599 (.O(FE_PHN2215_n599), 
	.I(n599));
   DELCKHD FE_PHC2214_n686 (.O(FE_PHN2214_n686), 
	.I(n686));
   DELCKHD FE_PHC2213_n4042 (.O(FE_PHN2213_n4042), 
	.I(n4042));
   DELCKHD FE_PHC2212_n675 (.O(FE_PHN2212_n675), 
	.I(n675));
   DELCKHD FE_PHC2211_n3405 (.O(FE_PHN2211_n3405), 
	.I(n3405));
   DELCKHD FE_PHC2210_n1632 (.O(FE_PHN2210_n1632), 
	.I(n1632));
   DELCKHD FE_PHC2209_n2328 (.O(FE_PHN2209_n2328), 
	.I(n2328));
   DELCKHD FE_PHC2208_n4654 (.O(FE_PHN2208_n4654), 
	.I(n4654));
   DELCKHD FE_PHC2207_n1314 (.O(FE_PHN2207_n1314), 
	.I(n1314));
   DELCKHD FE_PHC2206_n3599 (.O(FE_PHN2206_n3599), 
	.I(n3599));
   DELCKHD FE_PHC2205_n654 (.O(FE_PHN2205_n654), 
	.I(n654));
   DELCKHD FE_PHC2204_n1402 (.O(FE_PHN2204_n1402), 
	.I(n1402));
   DELCKHD FE_PHC2203_n2239 (.O(FE_PHN2203_n2239), 
	.I(n2239));
   DELCKHD FE_PHC2202_n1915 (.O(FE_PHN2202_n1915), 
	.I(n1915));
   DELCKHD FE_PHC2201_n1706 (.O(FE_PHN2201_n1706), 
	.I(n1706));
   DELCKHD FE_PHC2200_n1794 (.O(FE_PHN2200_n1794), 
	.I(n1794));
   DELCKHD FE_PHC2199_n3442 (.O(FE_PHN2199_n3442), 
	.I(n3442));
   DELCKHD FE_PHC2198_n2627 (.O(FE_PHN2198_n2627), 
	.I(n2627));
   DELCKHD FE_PHC2197_n1291 (.O(FE_PHN2197_n1291), 
	.I(n1291));
   DELCKHD FE_PHC2196_n2512 (.O(FE_PHN2196_n2512), 
	.I(n2512));
   DELCKHD FE_PHC2195_ram_199__5_ (.O(FE_PHN2195_ram_199__5_), 
	.I(\ram[199][5] ));
   DELCKHD FE_PHC2194_n3597 (.O(FE_PHN2194_n3597), 
	.I(n3597));
   DELCKHD FE_PHC2193_ram_132__8_ (.O(FE_PHN2193_ram_132__8_), 
	.I(\ram[132][8] ));
   DELCKHD FE_PHC2192_n3716 (.O(FE_PHN2192_n3716), 
	.I(n3716));
   DELCKHD FE_PHC2191_n2730 (.O(FE_PHN2191_n2730), 
	.I(n2730));
   DELCKHD FE_PHC2190_n1397 (.O(FE_PHN2190_n1397), 
	.I(n1397));
   DELCKHD FE_PHC2189_n2854 (.O(FE_PHN2189_n2854), 
	.I(n2854));
   DELCKHD FE_PHC2188_n1534 (.O(FE_PHN2188_n1534), 
	.I(n1534));
   DELCKHD FE_PHC2187_n2492 (.O(FE_PHN2187_n2492), 
	.I(n2492));
   DELCKHD FE_PHC2186_n4314 (.O(FE_PHN2186_n4314), 
	.I(n4314));
   DELCKHD FE_PHC2185_n1250 (.O(FE_PHN2185_n1250), 
	.I(n1250));
   DELCKHD FE_PHC2184_n3664 (.O(FE_PHN2184_n3664), 
	.I(n3664));
   DELCKHD FE_PHC2183_n2319 (.O(FE_PHN2183_n2319), 
	.I(n2319));
   DELCKHD FE_PHC2182_n3727 (.O(FE_PHN2182_n3727), 
	.I(n3727));
   DELCKHD FE_PHC2181_n1585 (.O(FE_PHN2181_n1585), 
	.I(n1585));
   DELCKHD FE_PHC2180_n2293 (.O(FE_PHN2180_n2293), 
	.I(n2293));
   DELCKHD FE_PHC2179_n1292 (.O(FE_PHN2179_n1292), 
	.I(n1292));
   DELCKHD FE_PHC2178_n1033 (.O(FE_PHN2178_n1033), 
	.I(n1033));
   DELCKHD FE_PHC2177_n1755 (.O(FE_PHN2177_n1755), 
	.I(n1755));
   DELCKHD FE_PHC2176_n2688 (.O(FE_PHN2176_n2688), 
	.I(n2688));
   DELCKHD FE_PHC2175_n4610 (.O(FE_PHN2175_n4610), 
	.I(n4610));
   DELCKHD FE_PHC2174_n2551 (.O(FE_PHN2174_n2551), 
	.I(n2551));
   DELCKHD FE_PHC2173_n2806 (.O(FE_PHN2173_n2806), 
	.I(n2806));
   DELCKHD FE_PHC2172_n2671 (.O(FE_PHN2172_n2671), 
	.I(n2671));
   DELCKHD FE_PHC2171_n2558 (.O(FE_PHN2171_n2558), 
	.I(n2558));
   DELCKHD FE_PHC2170_n783 (.O(FE_PHN2170_n783), 
	.I(n783));
   DELCKHD FE_PHC2169_n2694 (.O(FE_PHN2169_n2694), 
	.I(n2694));
   DELCKHD FE_PHC2168_n2661 (.O(FE_PHN2168_n2661), 
	.I(n2661));
   DELCKHD FE_PHC2167_n1610 (.O(FE_PHN2167_n1610), 
	.I(n1610));
   DELCKHD FE_PHC2166_n3345 (.O(FE_PHN2166_n3345), 
	.I(n3345));
   DELCKHD FE_PHC2165_n1193 (.O(FE_PHN2165_n1193), 
	.I(n1193));
   DELCKHD FE_PHC2164_n1323 (.O(FE_PHN2164_n1323), 
	.I(n1323));
   DELCKHD FE_PHC2163_n3602 (.O(FE_PHN2163_n3602), 
	.I(n3602));
   DELCKHD FE_PHC2162_n1712 (.O(FE_PHN2162_n1712), 
	.I(n1712));
   DELCKHD FE_PHC2161_n1514 (.O(FE_PHN2161_n1514), 
	.I(n1514));
   DELCKHD FE_PHC2160_n2707 (.O(FE_PHN2160_n2707), 
	.I(n2707));
   DELCKHD FE_PHC2159_n4221 (.O(FE_PHN2159_n4221), 
	.I(n4221));
   DELCKHD FE_PHC2158_n1639 (.O(FE_PHN2158_n1639), 
	.I(n1639));
   DELCKHD FE_PHC2157_n1199 (.O(FE_PHN2157_n1199), 
	.I(n1199));
   DELCKHD FE_PHC2156_n1338 (.O(FE_PHN2156_n1338), 
	.I(n1338));
   DELDKHD FE_PHC2155_n3385 (.O(FE_PHN2155_n3385), 
	.I(n3385));
   DELDKHD FE_PHC2154_n3799 (.O(FE_PHN2154_n3799), 
	.I(n3799));
   DELDKHD FE_PHC2153_n1304 (.O(FE_PHN2153_n1304), 
	.I(n1304));
   DELDKHD FE_PHC2152_n4649 (.O(FE_PHN2152_n4649), 
	.I(n4649));
   DELDKHD FE_PHC2151_n1658 (.O(FE_PHN2151_n1658), 
	.I(n1658));
   DELDKHD FE_PHC2150_n3770 (.O(FE_PHN2150_n3770), 
	.I(n3770));
   DELDKHD FE_PHC2149_n745 (.O(FE_PHN2149_n745), 
	.I(n745));
   DELDKHD FE_PHC2148_n4321 (.O(FE_PHN2148_n4321), 
	.I(n4321));
   DELDKHD FE_PHC2147_n3517 (.O(FE_PHN2147_n3517), 
	.I(n3517));
   DELDKHD FE_PHC2146_n2606 (.O(FE_PHN2146_n2606), 
	.I(n2606));
   DELDKHD FE_PHC2145_n1617 (.O(FE_PHN2145_n1617), 
	.I(n1617));
   DELDKHD FE_PHC2144_n4671 (.O(FE_PHN2144_n4671), 
	.I(n4671));
   DELDKHD FE_PHC2143_n1636 (.O(FE_PHN2143_n1636), 
	.I(n1636));
   DELDKHD FE_PHC2142_n3474 (.O(FE_PHN2142_n3474), 
	.I(n3474));
   DELDKHD FE_PHC2141_n1095 (.O(FE_PHN2141_n1095), 
	.I(n1095));
   DELDKHD FE_PHC2140_n2814 (.O(FE_PHN2140_n2814), 
	.I(n2814));
   DELDKHD FE_PHC2139_n1265 (.O(FE_PHN2139_n1265), 
	.I(n1265));
   DELDKHD FE_PHC2138_n668 (.O(FE_PHN2138_n668), 
	.I(n668));
   DELDKHD FE_PHC2137_n1606 (.O(FE_PHN2137_n1606), 
	.I(n1606));
   DELDKHD FE_PHC2136_n1297 (.O(FE_PHN2136_n1297), 
	.I(n1297));
   DELDKHD FE_PHC2135_n725 (.O(FE_PHN2135_n725), 
	.I(n725));
   DELDKHD FE_PHC2134_n2475 (.O(FE_PHN2134_n2475), 
	.I(n2475));
   DELDKHD FE_PHC2133_n3901 (.O(FE_PHN2133_n3901), 
	.I(n3901));
   DELDKHD FE_PHC2132_n1973 (.O(FE_PHN2132_n1973), 
	.I(n1973));
   DELDKHD FE_PHC2131_n1749 (.O(FE_PHN2131_n1749), 
	.I(n1749));
   DELDKHD FE_PHC2130_n2513 (.O(FE_PHN2130_n2513), 
	.I(n2513));
   DELDKHD FE_PHC2129_n3309 (.O(FE_PHN2129_n3309), 
	.I(n3309));
   DELDKHD FE_PHC2128_n1775 (.O(FE_PHN2128_n1775), 
	.I(n1775));
   DELDKHD FE_PHC2127_n1246 (.O(FE_PHN2127_n1246), 
	.I(n1246));
   DELDKHD FE_PHC2126_n3872 (.O(FE_PHN2126_n3872), 
	.I(n3872));
   DELDKHD FE_PHC2125_n4082 (.O(FE_PHN2125_n4082), 
	.I(n4082));
   DELDKHD FE_PHC2124_n1557 (.O(FE_PHN2124_n1557), 
	.I(n1557));
   DELDKHD FE_PHC2123_n1947 (.O(FE_PHN2123_n1947), 
	.I(n1947));
   DELDKHD FE_PHC2122_n2013 (.O(FE_PHN2122_n2013), 
	.I(n2013));
   DELDKHD FE_PHC2121_n1594 (.O(FE_PHN2121_n1594), 
	.I(n1594));
   DELDKHD FE_PHC2120_n2324 (.O(FE_PHN2120_n2324), 
	.I(n2324));
   DELDKHD FE_PHC2119_n2497 (.O(FE_PHN2119_n2497), 
	.I(n2497));
   DELDKHD FE_PHC2118_n2291 (.O(FE_PHN2118_n2291), 
	.I(n2291));
   DELDKHD FE_PHC2117_n637 (.O(FE_PHN2117_n637), 
	.I(n637));
   DELDKHD FE_PHC2116_n1270 (.O(FE_PHN2116_n1270), 
	.I(n1270));
   DELDKHD FE_PHC2115_n1346 (.O(FE_PHN2115_n1346), 
	.I(n1346));
   DELDKHD FE_PHC2114_n1391 (.O(FE_PHN2114_n1391), 
	.I(n1391));
   DELDKHD FE_PHC2113_n2216 (.O(FE_PHN2113_n2216), 
	.I(n2216));
   DELDKHD FE_PHC2112_n628 (.O(FE_PHN2112_n628), 
	.I(n628));
   DELDKHD FE_PHC2111_n2646 (.O(FE_PHN2111_n2646), 
	.I(n2646));
   DELDKHD FE_PHC2110_n1583 (.O(FE_PHN2110_n1583), 
	.I(n1583));
   DELDKHD FE_PHC2109_n3700 (.O(FE_PHN2109_n3700), 
	.I(n3700));
   DELDKHD FE_PHC2108_n1151 (.O(FE_PHN2108_n1151), 
	.I(n1151));
   DELDKHD FE_PHC2107_n2268 (.O(FE_PHN2107_n2268), 
	.I(n2268));
   DELDKHD FE_PHC2106_n1108 (.O(FE_PHN2106_n1108), 
	.I(n1108));
   DELDKHD FE_PHC2105_n636 (.O(FE_PHN2105_n636), 
	.I(n636));
   DELDKHD FE_PHC2104_n2199 (.O(FE_PHN2104_n2199), 
	.I(n2199));
   DELDKHD FE_PHC2103_n2096 (.O(FE_PHN2103_n2096), 
	.I(n2096));
   DELDKHD FE_PHC2102_n1635 (.O(FE_PHN2102_n1635), 
	.I(n1635));
   DELDKHD FE_PHC2101_n4637 (.O(FE_PHN2101_n4637), 
	.I(n4637));
   DELDKHD FE_PHC2100_n2202 (.O(FE_PHN2100_n2202), 
	.I(n2202));
   DELDKHD FE_PHC2099_n667 (.O(FE_PHN2099_n667), 
	.I(n667));
   DELDKHD FE_PHC2098_n2509 (.O(FE_PHN2098_n2509), 
	.I(n2509));
   DELDKHD FE_PHC2097_n1232 (.O(FE_PHN2097_n1232), 
	.I(n1232));
   DELDKHD FE_PHC2096_n1567 (.O(FE_PHN2096_n1567), 
	.I(n1567));
   DELDKHD FE_PHC2095_n2249 (.O(FE_PHN2095_n2249), 
	.I(n2249));
   DELDKHD FE_PHC2094_n3357 (.O(FE_PHN2094_n3357), 
	.I(n3357));
   DELDKHD FE_PHC2093_n4165 (.O(FE_PHN2093_n4165), 
	.I(n4165));
   DELDKHD FE_PHC2092_n2062 (.O(FE_PHN2092_n2062), 
	.I(n2062));
   DELDKHD FE_PHC2091_n2821 (.O(FE_PHN2091_n2821), 
	.I(n2821));
   DELDKHD FE_PHC2090_n2734 (.O(FE_PHN2090_n2734), 
	.I(n2734));
   DELDKHD FE_PHC2089_n3431 (.O(FE_PHN2089_n3431), 
	.I(n3431));
   DELDKHD FE_PHC2088_n669 (.O(FE_PHN2088_n669), 
	.I(n669));
   DELDKHD FE_PHC2087_n2318 (.O(FE_PHN2087_n2318), 
	.I(n2318));
   DELDKHD FE_PHC2086_n3390 (.O(FE_PHN2086_n3390), 
	.I(n3390));
   DELDKHD FE_PHC2085_n3655 (.O(FE_PHN2085_n3655), 
	.I(n3655));
   DELDKHD FE_PHC2084_n1168 (.O(FE_PHN2084_n1168), 
	.I(n1168));
   DELDKHD FE_PHC2083_n1981 (.O(FE_PHN2083_n1981), 
	.I(n1981));
   DELDKHD FE_PHC2082_n1220 (.O(FE_PHN2082_n1220), 
	.I(n1220));
   DELDKHD FE_PHC2081_n3594 (.O(FE_PHN2081_n3594), 
	.I(n3594));
   DELDKHD FE_PHC2080_n1179 (.O(FE_PHN2080_n1179), 
	.I(n1179));
   DELDKHD FE_PHC2079_n2843 (.O(FE_PHN2079_n2843), 
	.I(n2843));
   DELDKHD FE_PHC2078_n680 (.O(FE_PHN2078_n680), 
	.I(n680));
   DELDKHD FE_PHC2077_n2292 (.O(FE_PHN2077_n2292), 
	.I(n2292));
   DELDKHD FE_PHC2076_n656 (.O(FE_PHN2076_n656), 
	.I(n656));
   DELDKHD FE_PHC2075_n1169 (.O(FE_PHN2075_n1169), 
	.I(n1169));
   DELDKHD FE_PHC2074_n1424 (.O(FE_PHN2074_n1424), 
	.I(n1424));
   DELDKHD FE_PHC2073_n600 (.O(FE_PHN2073_n600), 
	.I(n600));
   DELDKHD FE_PHC2072_n2731 (.O(FE_PHN2072_n2731), 
	.I(n2731));
   DELDKHD FE_PHC2071_n1498 (.O(FE_PHN2071_n1498), 
	.I(n1498));
   DELDKHD FE_PHC2070_n1210 (.O(FE_PHN2070_n1210), 
	.I(n1210));
   DELDKHD FE_PHC2069_n1646 (.O(FE_PHN2069_n1646), 
	.I(n1646));
   DELDKHD FE_PHC2068_n956 (.O(FE_PHN2068_n956), 
	.I(n956));
   DELDKHD FE_PHC2067_n1414 (.O(FE_PHN2067_n1414), 
	.I(n1414));
   DELDKHD FE_PHC2066_n1990 (.O(FE_PHN2066_n1990), 
	.I(n1990));
   DELDKHD FE_PHC2065_n3410 (.O(FE_PHN2065_n3410), 
	.I(n3410));
   DELDKHD FE_PHC2064_n1537 (.O(FE_PHN2064_n1537), 
	.I(n1537));
   DELDKHD FE_PHC2063_n3477 (.O(FE_PHN2063_n3477), 
	.I(n3477));
   DELDKHD FE_PHC2062_n4661 (.O(FE_PHN2062_n4661), 
	.I(n4661));
   DELDKHD FE_PHC2061_n2056 (.O(FE_PHN2061_n2056), 
	.I(n2056));
   DELDKHD FE_PHC2060_n1768 (.O(FE_PHN2060_n1768), 
	.I(n1768));
   DELDKHD FE_PHC2059_n1312 (.O(FE_PHN2059_n1312), 
	.I(n1312));
   DELDKHD FE_PHC2058_n2547 (.O(FE_PHN2058_n2547), 
	.I(n2547));
   DELDKHD FE_PHC2057_n2287 (.O(FE_PHN2057_n2287), 
	.I(n2287));
   DELDKHD FE_PHC2056_n3204 (.O(FE_PHN2056_n3204), 
	.I(n3204));
   DELDKHD FE_PHC2055_n4117 (.O(FE_PHN2055_n4117), 
	.I(n4117));
   DELDKHD FE_PHC2054_n2080 (.O(FE_PHN2054_n2080), 
	.I(n2080));
   DELDKHD FE_PHC2053_n3729 (.O(FE_PHN2053_n3729), 
	.I(n3729));
   DELDKHD FE_PHC2052_n2690 (.O(FE_PHN2052_n2690), 
	.I(n2690));
   DELDKHD FE_PHC2051_n1995 (.O(FE_PHN2051_n1995), 
	.I(n1995));
   DELDKHD FE_PHC2050_n3174 (.O(FE_PHN2050_n3174), 
	.I(n3174));
   DELDKHD FE_PHC2049_n4585 (.O(FE_PHN2049_n4585), 
	.I(n4585));
   DELDKHD FE_PHC2048_n621 (.O(FE_PHN2048_n621), 
	.I(n621));
   DELDKHD FE_PHC2047_n3253 (.O(FE_PHN2047_n3253), 
	.I(n3253));
   DELDKHD FE_PHC2046_n3158 (.O(FE_PHN2046_n3158), 
	.I(n3158));
   DELDKHD FE_PHC2045_n3653 (.O(FE_PHN2045_n3653), 
	.I(n3653));
   DELDKHD FE_PHC2044_n1659 (.O(FE_PHN2044_n1659), 
	.I(n1659));
   DELDKHD FE_PHC2043_n2782 (.O(FE_PHN2043_n2782), 
	.I(n2782));
   DELDKHD FE_PHC2042_n4558 (.O(FE_PHN2042_n4558), 
	.I(n4558));
   DELDKHD FE_PHC2041_n1415 (.O(FE_PHN2041_n1415), 
	.I(n1415));
   DELDKHD FE_PHC2040_n2033 (.O(FE_PHN2040_n2033), 
	.I(n2033));
   DELDKHD FE_PHC2039_n2466 (.O(FE_PHN2039_n2466), 
	.I(n2466));
   DELDKHD FE_PHC2038_n2529 (.O(FE_PHN2038_n2529), 
	.I(n2529));
   DELDKHD FE_PHC2037_n661 (.O(FE_PHN2037_n661), 
	.I(n661));
   DELDKHD FE_PHC2036_n3764 (.O(FE_PHN2036_n3764), 
	.I(n3764));
   DELDKHD FE_PHC2035_n709 (.O(FE_PHN2035_n709), 
	.I(n709));
   DELDKHD FE_PHC2034_n2237 (.O(FE_PHN2034_n2237), 
	.I(n2237));
   DELDKHD FE_PHC2033_n3736 (.O(FE_PHN2033_n3736), 
	.I(n3736));
   DELDKHD FE_PHC2032_n1339 (.O(FE_PHN2032_n1339), 
	.I(n1339));
   DELDKHD FE_PHC2031_n703 (.O(FE_PHN2031_n703), 
	.I(n703));
   DELDKHD FE_PHC2030_n2768 (.O(FE_PHN2030_n2768), 
	.I(n2768));
   DELDKHD FE_PHC2029_n1209 (.O(FE_PHN2029_n1209), 
	.I(n1209));
   DELDKHD FE_PHC2028_n759 (.O(FE_PHN2028_n759), 
	.I(n759));
   DELDKHD FE_PHC2027_n2350 (.O(FE_PHN2027_n2350), 
	.I(n2350));
   DELDKHD FE_PHC2026_n1299 (.O(FE_PHN2026_n1299), 
	.I(n1299));
   DELDKHD FE_PHC2025_n4224 (.O(FE_PHN2025_n4224), 
	.I(n4224));
   DELDKHD FE_PHC2024_n815 (.O(FE_PHN2024_n815), 
	.I(n815));
   DELDKHD FE_PHC2023_n1736 (.O(FE_PHN2023_n1736), 
	.I(n1736));
   DELDKHD FE_PHC2022_n3590 (.O(FE_PHN2022_n3590), 
	.I(n3590));
   DELDKHD FE_PHC2021_n4562 (.O(FE_PHN2021_n4562), 
	.I(n4562));
   DELDKHD FE_PHC2020_n1967 (.O(FE_PHN2020_n1967), 
	.I(n1967));
   DELDKHD FE_PHC2019_n3269 (.O(FE_PHN2019_n3269), 
	.I(n3269));
   DELDKHD FE_PHC2018_n4628 (.O(FE_PHN2018_n4628), 
	.I(n4628));
   DELDKHD FE_PHC2017_n4647 (.O(FE_PHN2017_n4647), 
	.I(n4647));
   DELDKHD FE_PHC2016_n2449 (.O(FE_PHN2016_n2449), 
	.I(n2449));
   DELDKHD FE_PHC2015_n2884 (.O(FE_PHN2015_n2884), 
	.I(n2884));
   DELDKHD FE_PHC2014_n2099 (.O(FE_PHN2014_n2099), 
	.I(n2099));
   DELDKHD FE_PHC2013_n1590 (.O(FE_PHN2013_n1590), 
	.I(n1590));
   DELDKHD FE_PHC2012_n1766 (.O(FE_PHN2012_n1766), 
	.I(n1766));
   DELDKHD FE_PHC2011_n2110 (.O(FE_PHN2011_n2110), 
	.I(n2110));
   DELDKHD FE_PHC2010_n597 (.O(FE_PHN2010_n597), 
	.I(n597));
   DELDKHD FE_PHC2009_n1377 (.O(FE_PHN2009_n1377), 
	.I(n1377));
   DELDKHD FE_PHC2008_n2832 (.O(FE_PHN2008_n2832), 
	.I(n2832));
   DELDKHD FE_PHC2007_n4648 (.O(FE_PHN2007_n4648), 
	.I(n4648));
   DELDKHD FE_PHC2006_n4640 (.O(FE_PHN2006_n4640), 
	.I(n4640));
   DELDKHD FE_PHC2005_ram_202__13_ (.O(FE_PHN2005_ram_202__13_), 
	.I(\ram[202][13] ));
   DELDKHD FE_PHC2004_n1319 (.O(FE_PHN2004_n1319), 
	.I(n1319));
   DELDKHD FE_PHC2003_n648 (.O(FE_PHN2003_n648), 
	.I(n648));
   DELDKHD FE_PHC2002_n1966 (.O(FE_PHN2002_n1966), 
	.I(n1966));
   DELDKHD FE_PHC2001_n4346 (.O(FE_PHN2001_n4346), 
	.I(n4346));
   DELDKHD FE_PHC2000_n1998 (.O(FE_PHN2000_n1998), 
	.I(n1998));
   DELDKHD FE_PHC1999_n2252 (.O(FE_PHN1999_n2252), 
	.I(n2252));
   DELDKHD FE_PHC1998_n1091 (.O(FE_PHN1998_n1091), 
	.I(n1091));
   DELDKHD FE_PHC1997_n2556 (.O(FE_PHN1997_n2556), 
	.I(n2556));
   DELDKHD FE_PHC1996_n762 (.O(FE_PHN1996_n762), 
	.I(n762));
   DELDKHD FE_PHC1995_n2874 (.O(FE_PHN1995_n2874), 
	.I(n2874));
   DELDKHD FE_PHC1994_n3824 (.O(FE_PHN1994_n3824), 
	.I(n3824));
   DELDKHD FE_PHC1993_n1285 (.O(FE_PHN1993_n1285), 
	.I(n1285));
   DELDKHD FE_PHC1992_n3775 (.O(FE_PHN1992_n3775), 
	.I(n3775));
   DELDKHD FE_PHC1991_n3382 (.O(FE_PHN1991_n3382), 
	.I(n3382));
   DELDKHD FE_PHC1990_n1586 (.O(FE_PHN1990_n1586), 
	.I(n1586));
   DELDKHD FE_PHC1989_n1756 (.O(FE_PHN1989_n1756), 
	.I(n1756));
   DELDKHD FE_PHC1988_n4298 (.O(FE_PHN1988_n4298), 
	.I(n4298));
   DELDKHD FE_PHC1987_n1159 (.O(FE_PHN1987_n1159), 
	.I(n1159));
   DELDKHD FE_PHC1986_n1605 (.O(FE_PHN1986_n1605), 
	.I(n1605));
   DELDKHD FE_PHC1985_n3420 (.O(FE_PHN1985_n3420), 
	.I(n3420));
   DELDKHD FE_PHC1984_n3671 (.O(FE_PHN1984_n3671), 
	.I(n3671));
   DELDKHD FE_PHC1983_n1396 (.O(FE_PHN1983_n1396), 
	.I(n1396));
   DELDKHD FE_PHC1982_n2014 (.O(FE_PHN1982_n2014), 
	.I(n2014));
   DELDKHD FE_PHC1981_n1620 (.O(FE_PHN1981_n1620), 
	.I(n1620));
   DELDKHD FE_PHC1980_n2076 (.O(FE_PHN1980_n2076), 
	.I(n2076));
   DELDKHD FE_PHC1979_n1648 (.O(FE_PHN1979_n1648), 
	.I(n1648));
   DELDKHD FE_PHC1978_n2298 (.O(FE_PHN1978_n2298), 
	.I(n2298));
   DELDKHD FE_PHC1977_n1334 (.O(FE_PHN1977_n1334), 
	.I(n1334));
   DELDKHD FE_PHC1976_n3715 (.O(FE_PHN1976_n3715), 
	.I(n3715));
   DELDKHD FE_PHC1975_n822 (.O(FE_PHN1975_n822), 
	.I(n822));
   DELDKHD FE_PHC1974_n2357 (.O(FE_PHN1974_n2357), 
	.I(n2357));
   DELDKHD FE_PHC1973_n2552 (.O(FE_PHN1973_n2552), 
	.I(n2552));
   DELDKHD FE_PHC1972_n2058 (.O(FE_PHN1972_n2058), 
	.I(n2058));
   DELDKHD FE_PHC1971_n3416 (.O(FE_PHN1971_n3416), 
	.I(n3416));
   DELDKHD FE_PHC1970_n3902 (.O(FE_PHN1970_n3902), 
	.I(n3902));
   DELDKHD FE_PHC1969_n1999 (.O(FE_PHN1969_n1999), 
	.I(n1999));
   DELDKHD FE_PHC1968_n2748 (.O(FE_PHN1968_n2748), 
	.I(n2748));
   DELDKHD FE_PHC1967_n1527 (.O(FE_PHN1967_n1527), 
	.I(n1527));
   DELDKHD FE_PHC1966_n1393 (.O(FE_PHN1966_n1393), 
	.I(n1393));
   DELDKHD FE_PHC1965_n4074 (.O(FE_PHN1965_n4074), 
	.I(n4074));
   DELCKHD FE_PHC1964_n2650 (.O(FE_PHN1964_n2650), 
	.I(n2650));
   DELCKHD FE_PHC1963_n3790 (.O(FE_PHN1963_n3790), 
	.I(n3790));
   DELCKHD FE_PHC1962_ram_85__10_ (.O(FE_PHN1962_ram_85__10_), 
	.I(\ram[85][10] ));
   DELCKHD FE_PHC1961_n4115 (.O(FE_PHN1961_n4115), 
	.I(n4115));
   DELCKHD FE_PHC1960_n3221 (.O(FE_PHN1960_n3221), 
	.I(n3221));
   DELCKHD FE_PHC1959_n1136 (.O(FE_PHN1959_n1136), 
	.I(n1136));
   DELCKHD FE_PHC1958_n4489 (.O(FE_PHN1958_n4489), 
	.I(n4489));
   DELCKHD FE_PHC1957_n3516 (.O(FE_PHN1957_n3516), 
	.I(n3516));
   DELCKHD FE_PHC1956_n695 (.O(FE_PHN1956_n695), 
	.I(n695));
   DELCKHD FE_PHC1955_n1839 (.O(FE_PHN1955_n1839), 
	.I(n1839));
   DELCKHD FE_PHC1954_n720 (.O(FE_PHN1954_n720), 
	.I(n720));
   DELCKHD FE_PHC1953_n2286 (.O(FE_PHN1953_n2286), 
	.I(n2286));
   DELCKHD FE_PHC1952_n714 (.O(FE_PHN1952_n714), 
	.I(n714));
   DELCKHD FE_PHC1951_n2645 (.O(FE_PHN1951_n2645), 
	.I(n2645));
   DELCKHD FE_PHC1950_n2329 (.O(FE_PHN1950_n2329), 
	.I(n2329));
   DELCKHD FE_PHC1949_n3496 (.O(FE_PHN1949_n3496), 
	.I(n3496));
   DELCKHD FE_PHC1948_n1141 (.O(FE_PHN1948_n1141), 
	.I(n1141));
   DELCKHD FE_PHC1947_n2752 (.O(FE_PHN1947_n2752), 
	.I(n2752));
   DELCKHD FE_PHC1946_n4101 (.O(FE_PHN1946_n4101), 
	.I(n4101));
   DELCKHD FE_PHC1945_n2064 (.O(FE_PHN1945_n2064), 
	.I(n2064));
   DELCKHD FE_PHC1944_n2372 (.O(FE_PHN1944_n2372), 
	.I(n2372));
   DELCKHD FE_PHC1943_n1928 (.O(FE_PHN1943_n1928), 
	.I(n1928));
   DELCKHD FE_PHC1942_n2482 (.O(FE_PHN1942_n2482), 
	.I(n2482));
   DELCKHD FE_PHC1941_n1418 (.O(FE_PHN1941_n1418), 
	.I(n1418));
   DELCKHD FE_PHC1940_n718 (.O(FE_PHN1940_n718), 
	.I(n718));
   DELCKHD FE_PHC1939_n1979 (.O(FE_PHN1939_n1979), 
	.I(n1979));
   DELCKHD FE_PHC1938_n2010 (.O(FE_PHN1938_n2010), 
	.I(n2010));
   DELCKHD FE_PHC1937_n1497 (.O(FE_PHN1937_n1497), 
	.I(n1497));
   DELCKHD FE_PHC1936_n3852 (.O(FE_PHN1936_n3852), 
	.I(n3852));
   DELCKHD FE_PHC1935_n3884 (.O(FE_PHN1935_n3884), 
	.I(n3884));
   DELCKHD FE_PHC1934_n722 (.O(FE_PHN1934_n722), 
	.I(n722));
   DELCKHD FE_PHC1933_n4357 (.O(FE_PHN1933_n4357), 
	.I(n4357));
   DELCKHD FE_PHC1932_n1261 (.O(FE_PHN1932_n1261), 
	.I(n1261));
   DELCKHD FE_PHC1931_n1678 (.O(FE_PHN1931_n1678), 
	.I(n1678));
   DELCKHD FE_PHC1930_n3719 (.O(FE_PHN1930_n3719), 
	.I(n3719));
   DELCKHD FE_PHC1929_n4303 (.O(FE_PHN1929_n4303), 
	.I(n4303));
   DELCKHD FE_PHC1928_n2515 (.O(FE_PHN1928_n2515), 
	.I(n2515));
   DELCKHD FE_PHC1927_n3247 (.O(FE_PHN1927_n3247), 
	.I(n3247));
   DELCKHD FE_PHC1926_n3637 (.O(FE_PHN1926_n3637), 
	.I(n3637));
   DELCKHD FE_PHC1925_n1582 (.O(FE_PHN1925_n1582), 
	.I(n1582));
   DELCKHD FE_PHC1924_n2676 (.O(FE_PHN1924_n2676), 
	.I(n2676));
   DELCKHD FE_PHC1923_n4131 (.O(FE_PHN1923_n4131), 
	.I(n4131));
   DELCKHD FE_PHC1922_n682 (.O(FE_PHN1922_n682), 
	.I(n682));
   DELCKHD FE_PHC1921_n2106 (.O(FE_PHN1921_n2106), 
	.I(n2106));
   DELCKHD FE_PHC1920_n1041 (.O(FE_PHN1920_n1041), 
	.I(n1041));
   DELCKHD FE_PHC1919_n1564 (.O(FE_PHN1919_n1564), 
	.I(n1564));
   DELCKHD FE_PHC1918_n1237 (.O(FE_PHN1918_n1237), 
	.I(n1237));
   DELCKHD FE_PHC1917_n1954 (.O(FE_PHN1917_n1954), 
	.I(n1954));
   DELCKHD FE_PHC1916_n4200 (.O(FE_PHN1916_n4200), 
	.I(n4200));
   DELCKHD FE_PHC1915_n4559 (.O(FE_PHN1915_n4559), 
	.I(n4559));
   DELCKHD FE_PHC1914_n3225 (.O(FE_PHN1914_n3225), 
	.I(n3225));
   DELCKHD FE_PHC1913_n2316 (.O(FE_PHN1913_n2316), 
	.I(n2316));
   DELCKHD FE_PHC1912_n3833 (.O(FE_PHN1912_n3833), 
	.I(n3833));
   DELCKHD FE_PHC1911_n2347 (.O(FE_PHN1911_n2347), 
	.I(n2347));
   DELCKHD FE_PHC1910_n3381 (.O(FE_PHN1910_n3381), 
	.I(n3381));
   DELCKHD FE_PHC1909_n3290 (.O(FE_PHN1909_n3290), 
	.I(n3290));
   DELCKHD FE_PHC1908_n2698 (.O(FE_PHN1908_n2698), 
	.I(n2698));
   DELCKHD FE_PHC1907_n808 (.O(FE_PHN1907_n808), 
	.I(n808));
   DELCKHD FE_PHC1906_n2689 (.O(FE_PHN1906_n2689), 
	.I(n2689));
   DELCKHD FE_PHC1905_n1884 (.O(FE_PHN1905_n1884), 
	.I(n1884));
   DELCKHD FE_PHC1904_n3181 (.O(FE_PHN1904_n3181), 
	.I(n3181));
   DELCKHD FE_PHC1903_n1860 (.O(FE_PHN1903_n1860), 
	.I(n1860));
   DELCKHD FE_PHC1902_n2810 (.O(FE_PHN1902_n2810), 
	.I(n2810));
   DELCKHD FE_PHC1901_n3211 (.O(FE_PHN1901_n3211), 
	.I(n3211));
   DELCKHD FE_PHC1900_n3177 (.O(FE_PHN1900_n3177), 
	.I(n3177));
   DELCKHD FE_PHC1899_n923 (.O(FE_PHN1899_n923), 
	.I(n923));
   DELCKHD FE_PHC1898_n2709 (.O(FE_PHN1898_n2709), 
	.I(n2709));
   DELCKHD FE_PHC1897_n1410 (.O(FE_PHN1897_n1410), 
	.I(n1410));
   DELCKHD FE_PHC1896_n4490 (.O(FE_PHN1896_n4490), 
	.I(n4490));
   DELCKHD FE_PHC1895_n3502 (.O(FE_PHN1895_n3502), 
	.I(n3502));
   DELCKHD FE_PHC1894_n1258 (.O(FE_PHN1894_n1258), 
	.I(n1258));
   DELCKHD FE_PHC1893_n1679 (.O(FE_PHN1893_n1679), 
	.I(n1679));
   DELCKHD FE_PHC1892_n1372 (.O(FE_PHN1892_n1372), 
	.I(n1372));
   DELCKHD FE_PHC1891_n2830 (.O(FE_PHN1891_n2830), 
	.I(n2830));
   DELCKHD FE_PHC1890_n3904 (.O(FE_PHN1890_n3904), 
	.I(n3904));
   DELCKHD FE_PHC1889_n1729 (.O(FE_PHN1889_n1729), 
	.I(n1729));
   DELCKHD FE_PHC1888_n1925 (.O(FE_PHN1888_n1925), 
	.I(n1925));
   DELCKHD FE_PHC1887_n1986 (.O(FE_PHN1887_n1986), 
	.I(n1986));
   DELCKHD FE_PHC1886_n2451 (.O(FE_PHN1886_n2451), 
	.I(n2451));
   DELCKHD FE_PHC1885_n4454 (.O(FE_PHN1885_n4454), 
	.I(n4454));
   DELCKHD FE_PHC1884_n3601 (.O(FE_PHN1884_n3601), 
	.I(n3601));
   DELCKHD FE_PHC1883_n2450 (.O(FE_PHN1883_n2450), 
	.I(n2450));
   DELCKHD FE_PHC1882_n1641 (.O(FE_PHN1882_n1641), 
	.I(n1641));
   DELCKHD FE_PHC1881_n817 (.O(FE_PHN1881_n817), 
	.I(n817));
   DELCKHD FE_PHC1880_n4336 (.O(FE_PHN1880_n4336), 
	.I(n4336));
   DELCKHD FE_PHC1879_n1139 (.O(FE_PHN1879_n1139), 
	.I(n1139));
   DELCKHD FE_PHC1878_n1388 (.O(FE_PHN1878_n1388), 
	.I(n1388));
   DELCKHD FE_PHC1877_n3667 (.O(FE_PHN1877_n3667), 
	.I(n3667));
   DELCKHD FE_PHC1876_n3906 (.O(FE_PHN1876_n3906), 
	.I(n3906));
   DELCKHD FE_PHC1875_n2301 (.O(FE_PHN1875_n2301), 
	.I(n2301));
   DELCKHD FE_PHC1874_n883 (.O(FE_PHN1874_n883), 
	.I(n883));
   DELCKHD FE_PHC1873_n4351 (.O(FE_PHN1873_n4351), 
	.I(n4351));
   DELCKHD FE_PHC1872_n787 (.O(FE_PHN1872_n787), 
	.I(n787));
   DELCKHD FE_PHC1871_n3193 (.O(FE_PHN1871_n3193), 
	.I(n3193));
   DELCKHD FE_PHC1870_n4650 (.O(FE_PHN1870_n4650), 
	.I(n4650));
   DELCKHD FE_PHC1869_n4526 (.O(FE_PHN1869_n4526), 
	.I(n4526));
   DELCKHD FE_PHC1868_n1539 (.O(FE_PHN1868_n1539), 
	.I(n1539));
   DELCKHD FE_PHC1867_n1933 (.O(FE_PHN1867_n1933), 
	.I(n1933));
   DELCKHD FE_PHC1866_n3559 (.O(FE_PHN1866_n3559), 
	.I(n3559));
   DELCKHD FE_PHC1865_n4551 (.O(FE_PHN1865_n4551), 
	.I(n4551));
   DELCKHD FE_PHC1864_n1234 (.O(FE_PHN1864_n1234), 
	.I(n1234));
   DELCKHD FE_PHC1863_n2225 (.O(FE_PHN1863_n2225), 
	.I(n2225));
   DELCKHD FE_PHC1862_n2290 (.O(FE_PHN1862_n2290), 
	.I(n2290));
   DELCKHD FE_PHC1861_n2045 (.O(FE_PHN1861_n2045), 
	.I(n2045));
   DELCKHD FE_PHC1860_n2371 (.O(FE_PHN1860_n2371), 
	.I(n2371));
   DELCKHD FE_PHC1859_n2263 (.O(FE_PHN1859_n2263), 
	.I(n2263));
   DELCKHD FE_PHC1858_n3605 (.O(FE_PHN1858_n3605), 
	.I(n3605));
   DELCKHD FE_PHC1857_n3661 (.O(FE_PHN1857_n3661), 
	.I(n3661));
   DELCKHD FE_PHC1856_n792 (.O(FE_PHN1856_n792), 
	.I(n792));
   DELCKHD FE_PHC1855_n2772 (.O(FE_PHN1855_n2772), 
	.I(n2772));
   DELCKHD FE_PHC1854_n2295 (.O(FE_PHN1854_n2295), 
	.I(n2295));
   DELCKHD FE_PHC1853_n1516 (.O(FE_PHN1853_n1516), 
	.I(n1516));
   DELCKHD FE_PHC1852_n4189 (.O(FE_PHN1852_n4189), 
	.I(n4189));
   DELCKHD FE_PHC1851_n3369 (.O(FE_PHN1851_n3369), 
	.I(n3369));
   DELCKHD FE_PHC1850_n1333 (.O(FE_PHN1850_n1333), 
	.I(n1333));
   DELCKHD FE_PHC1849_n3240 (.O(FE_PHN1849_n3240), 
	.I(n3240));
   DELCKHD FE_PHC1848_n1852 (.O(FE_PHN1848_n1852), 
	.I(n1852));
   DELCKHD FE_PHC1847_n4674 (.O(FE_PHN1847_n4674), 
	.I(n4674));
   DELCKHD FE_PHC1846_n2353 (.O(FE_PHN1846_n2353), 
	.I(n2353));
   DELCKHD FE_PHC1845_n3407 (.O(FE_PHN1845_n3407), 
	.I(n3407));
   DELCKHD FE_PHC1844_n3850 (.O(FE_PHN1844_n3850), 
	.I(n3850));
   DELCKHD FE_PHC1843_n3642 (.O(FE_PHN1843_n3642), 
	.I(n3642));
   DELCKHD FE_PHC1842_n2878 (.O(FE_PHN1842_n2878), 
	.I(n2878));
   DELCKHD FE_PHC1841_n2114 (.O(FE_PHN1841_n2114), 
	.I(n2114));
   DELCKHD FE_PHC1840_n4619 (.O(FE_PHN1840_n4619), 
	.I(n4619));
   DELCKHD FE_PHC1839_n1649 (.O(FE_PHN1839_n1649), 
	.I(n1649));
   DELCKHD FE_PHC1838_n3184 (.O(FE_PHN1838_n3184), 
	.I(n3184));
   DELCKHD FE_PHC1837_n630 (.O(FE_PHN1837_n630), 
	.I(n630));
   DELCKHD FE_PHC1836_n1535 (.O(FE_PHN1836_n1535), 
	.I(n1535));
   DELCKHD FE_PHC1835_n1664 (.O(FE_PHN1835_n1664), 
	.I(n1664));
   DELCKHD FE_PHC1834_n1011 (.O(FE_PHN1834_n1011), 
	.I(n1011));
   DELCKHD FE_PHC1833_n2847 (.O(FE_PHN1833_n2847), 
	.I(n2847));
   DELCKHD FE_PHC1832_n3460 (.O(FE_PHN1832_n3460), 
	.I(n3460));
   DELCKHD FE_PHC1831_n3436 (.O(FE_PHN1831_n3436), 
	.I(n3436));
   DELCKHD FE_PHC1830_n3444 (.O(FE_PHN1830_n3444), 
	.I(n3444));
   DELCKHD FE_PHC1829_n1412 (.O(FE_PHN1829_n1412), 
	.I(n1412));
   DELCKHD FE_PHC1828_n3869 (.O(FE_PHN1828_n3869), 
	.I(n3869));
   DELCKHD FE_PHC1827_n2729 (.O(FE_PHN1827_n2729), 
	.I(n2729));
   DELCKHD FE_PHC1826_n1473 (.O(FE_PHN1826_n1473), 
	.I(n1473));
   DELCKHD FE_PHC1825_n3278 (.O(FE_PHN1825_n3278), 
	.I(n3278));
   DELCKHD FE_PHC1824_n824 (.O(FE_PHN1824_n824), 
	.I(n824));
   DELCKHD FE_PHC1823_n3585 (.O(FE_PHN1823_n3585), 
	.I(n3585));
   DELCKHD FE_PHC1822_n1738 (.O(FE_PHN1822_n1738), 
	.I(n1738));
   DELCKHD FE_PHC1821_n2742 (.O(FE_PHN1821_n2742), 
	.I(n2742));
   DELCKHD FE_PHC1820_n1495 (.O(FE_PHN1820_n1495), 
	.I(n1495));
   DELCKHD FE_PHC1819_n1810 (.O(FE_PHN1819_n1810), 
	.I(n1810));
   DELCKHD FE_PHC1818_n3527 (.O(FE_PHN1818_n3527), 
	.I(n3527));
   DELCKHD FE_PHC1817_n2182 (.O(FE_PHN1817_n2182), 
	.I(n2182));
   DELCKHD FE_PHC1816_n2913 (.O(FE_PHN1816_n2913), 
	.I(n2913));
   DELCKHD FE_PHC1815_n1122 (.O(FE_PHN1815_n1122), 
	.I(n1122));
   DELCKHD FE_PHC1814_n2373 (.O(FE_PHN1814_n2373), 
	.I(n2373));
   DELCKHD FE_PHC1813_n3787 (.O(FE_PHN1813_n3787), 
	.I(n3787));
   DELCKHD FE_PHC1812_n1039 (.O(FE_PHN1812_n1039), 
	.I(n1039));
   DELCKHD FE_PHC1811_n3178 (.O(FE_PHN1811_n3178), 
	.I(n3178));
   DELCKHD FE_PHC1810_n2827 (.O(FE_PHN1810_n2827), 
	.I(n2827));
   DELCKHD FE_PHC1809_n4491 (.O(FE_PHN1809_n4491), 
	.I(n4491));
   DELCKHD FE_PHC1808_n2108 (.O(FE_PHN1808_n2108), 
	.I(n2108));
   DELCKHD FE_PHC1807_n2469 (.O(FE_PHN1807_n2469), 
	.I(n2469));
   DELCKHD FE_PHC1806_n3160 (.O(FE_PHN1806_n3160), 
	.I(n3160));
   DELCKHD FE_PHC1805_n4520 (.O(FE_PHN1805_n4520), 
	.I(n4520));
   DELCKHD FE_PHC1804_n690 (.O(FE_PHN1804_n690), 
	.I(n690));
   DELCKHD FE_PHC1803_n726 (.O(FE_PHN1803_n726), 
	.I(n726));
   DELCKHD FE_PHC1802_n3293 (.O(FE_PHN1802_n3293), 
	.I(n3293));
   DELCKHD FE_PHC1801_n807 (.O(FE_PHN1801_n807), 
	.I(n807));
   DELCKHD FE_PHC1800_n3900 (.O(FE_PHN1800_n3900), 
	.I(n3900));
   DELCKHD FE_PHC1799_n1275 (.O(FE_PHN1799_n1275), 
	.I(n1275));
   DELCKHD FE_PHC1798_n3593 (.O(FE_PHN1798_n3593), 
	.I(n3593));
   DELCKHD FE_PHC1797_n1560 (.O(FE_PHN1797_n1560), 
	.I(n1560));
   DELCKHD FE_PHC1796_n1836 (.O(FE_PHN1796_n1836), 
	.I(n1836));
   DELCKHD FE_PHC1795_n2668 (.O(FE_PHN1795_n2668), 
	.I(n2668));
   DELCKHD FE_PHC1794_n1173 (.O(FE_PHN1794_n1173), 
	.I(n1173));
   DELCKHD FE_PHC1793_n2595 (.O(FE_PHN1793_n2595), 
	.I(n2595));
   DELCKHD FE_PHC1792_n1321 (.O(FE_PHN1792_n1321), 
	.I(n1321));
   DELCKHD FE_PHC1791_n772 (.O(FE_PHN1791_n772), 
	.I(n772));
   DELCKHD FE_PHC1790_n3662 (.O(FE_PHN1790_n3662), 
	.I(n3662));
   DELCKHD FE_PHC1789_n1305 (.O(FE_PHN1789_n1305), 
	.I(n1305));
   DELCKHD FE_PHC1788_n1960 (.O(FE_PHN1788_n1960), 
	.I(n1960));
   DELCKHD FE_PHC1787_n3412 (.O(FE_PHN1787_n3412), 
	.I(n3412));
   DELCKHD FE_PHC1786_n704 (.O(FE_PHN1786_n704), 
	.I(n704));
   DELCKHD FE_PHC1785_n3428 (.O(FE_PHN1785_n3428), 
	.I(n3428));
   DELCKHD FE_PHC1784_n2028 (.O(FE_PHN1784_n2028), 
	.I(n2028));
   DELCKHD FE_PHC1783_n4237 (.O(FE_PHN1783_n4237), 
	.I(n4237));
   DELDKHD FE_PHC1782_n3612 (.O(FE_PHN1782_n3612), 
	.I(n3612));
   DELDKHD FE_PHC1781_ram_63__5_ (.O(FE_PHN1781_ram_63__5_), 
	.I(\ram[63][5] ));
   DELDKHD FE_PHC1780_n1842 (.O(FE_PHN1780_n1842), 
	.I(n1842));
   DELDKHD FE_PHC1779_n4045 (.O(FE_PHN1779_n4045), 
	.I(n4045));
   DELDKHD FE_PHC1778_ram_61__13_ (.O(FE_PHN1778_ram_61__13_), 
	.I(\ram[61][13] ));
   DELDKHD FE_PHC1777_n3270 (.O(FE_PHN1777_n3270), 
	.I(n3270));
   DELDKHD FE_PHC1776_n2686 (.O(FE_PHN1776_n2686), 
	.I(n2686));
   DELDKHD FE_PHC1775_n1793 (.O(FE_PHN1775_n1793), 
	.I(n1793));
   DELDKHD FE_PHC1774_n3146 (.O(FE_PHN1774_n3146), 
	.I(n3146));
   DELDKHD FE_PHC1773_n3718 (.O(FE_PHN1773_n3718), 
	.I(n3718));
   DELDKHD FE_PHC1772_n670 (.O(FE_PHN1772_n670), 
	.I(n670));
   DELDKHD FE_PHC1771_n3452 (.O(FE_PHN1771_n3452), 
	.I(n3452));
   DELDKHD FE_PHC1770_n4059 (.O(FE_PHN1770_n4059), 
	.I(n4059));
   DELDKHD FE_PHC1769_n4152 (.O(FE_PHN1769_n4152), 
	.I(n4152));
   DELDKHD FE_PHC1768_n3359 (.O(FE_PHN1768_n3359), 
	.I(n3359));
   DELDKHD FE_PHC1767_n4122 (.O(FE_PHN1767_n4122), 
	.I(n4122));
   DELDKHD FE_PHC1766_n4145 (.O(FE_PHN1766_n4145), 
	.I(n4145));
   DELDKHD FE_PHC1765_n3446 (.O(FE_PHN1765_n3446), 
	.I(n3446));
   DELDKHD FE_PHC1764_n3586 (.O(FE_PHN1764_n3586), 
	.I(n3586));
   DELDKHD FE_PHC1763_n1477 (.O(FE_PHN1763_n1477), 
	.I(n1477));
   DELDKHD FE_PHC1762_n4192 (.O(FE_PHN1762_n4192), 
	.I(n4192));
   DELDKHD FE_PHC1761_n4564 (.O(FE_PHN1761_n4564), 
	.I(n4564));
   DELDKHD FE_PHC1760_n4184 (.O(FE_PHN1760_n4184), 
	.I(n4184));
   DELDKHD FE_PHC1759_n608 (.O(FE_PHN1759_n608), 
	.I(n608));
   DELDKHD FE_PHC1758_n1724 (.O(FE_PHN1758_n1724), 
	.I(n1724));
   DELDKHD FE_PHC1757_n4442 (.O(FE_PHN1757_n4442), 
	.I(n4442));
   DELDKHD FE_PHC1756_n4608 (.O(FE_PHN1756_n4608), 
	.I(n4608));
   DELDKHD FE_PHC1755_n2279 (.O(FE_PHN1755_n2279), 
	.I(n2279));
   DELDKHD FE_PHC1754_n2879 (.O(FE_PHN1754_n2879), 
	.I(n2879));
   DELDKHD FE_PHC1753_n1174 (.O(FE_PHN1753_n1174), 
	.I(n1174));
   DELDKHD FE_PHC1752_n2764 (.O(FE_PHN1752_n2764), 
	.I(n2764));
   DELDKHD FE_PHC1751_n3847 (.O(FE_PHN1751_n3847), 
	.I(n3847));
   DELDKHD FE_PHC1750_n3695 (.O(FE_PHN1750_n3695), 
	.I(n3695));
   DELDKHD FE_PHC1749_n4052 (.O(FE_PHN1749_n4052), 
	.I(n4052));
   DELDKHD FE_PHC1748_n4467 (.O(FE_PHN1748_n4467), 
	.I(n4467));
   DELDKHD FE_PHC1747_n1282 (.O(FE_PHN1747_n1282), 
	.I(n1282));
   DELDKHD FE_PHC1746_n4484 (.O(FE_PHN1746_n4484), 
	.I(n4484));
   DELDKHD FE_PHC1745_n2034 (.O(FE_PHN1745_n2034), 
	.I(n2034));
   DELDKHD FE_PHC1744_n591 (.O(FE_PHN1744_n591), 
	.I(n591));
   DELDKHD FE_PHC1743_n1368 (.O(FE_PHN1743_n1368), 
	.I(n1368));
   DELDKHD FE_PHC1742_n3206 (.O(FE_PHN1742_n3206), 
	.I(n3206));
   DELDKHD FE_PHC1741_n3256 (.O(FE_PHN1741_n3256), 
	.I(n3256));
   DELDKHD FE_PHC1740_n1971 (.O(FE_PHN1740_n1971), 
	.I(n1971));
   DELDKHD FE_PHC1739_n2000 (.O(FE_PHN1739_n2000), 
	.I(n2000));
   DELDKHD FE_PHC1738_n3281 (.O(FE_PHN1738_n3281), 
	.I(n3281));
   DELDKHD FE_PHC1737_n674 (.O(FE_PHN1737_n674), 
	.I(n674));
   DELDKHD FE_PHC1736_n1549 (.O(FE_PHN1736_n1549), 
	.I(n1549));
   DELDKHD FE_PHC1735_n4584 (.O(FE_PHN1735_n4584), 
	.I(n4584));
   DELDKHD FE_PHC1734_n3666 (.O(FE_PHN1734_n3666), 
	.I(n3666));
   DELDKHD FE_PHC1733_n2255 (.O(FE_PHN1733_n2255), 
	.I(n2255));
   DELDKHD FE_PHC1732_n1244 (.O(FE_PHN1732_n1244), 
	.I(n1244));
   DELDKHD FE_PHC1731_n2737 (.O(FE_PHN1731_n2737), 
	.I(n2737));
   DELDKHD FE_PHC1730_n3627 (.O(FE_PHN1730_n3627), 
	.I(n3627));
   DELDKHD FE_PHC1729_n2026 (.O(FE_PHN1729_n2026), 
	.I(n2026));
   DELDKHD FE_PHC1728_n3439 (.O(FE_PHN1728_n3439), 
	.I(n3439));
   DELDKHD FE_PHC1727_n644 (.O(FE_PHN1727_n644), 
	.I(n644));
   DELDKHD FE_PHC1726_n1226 (.O(FE_PHN1726_n1226), 
	.I(n1226));
   DELDKHD FE_PHC1725_n1295 (.O(FE_PHN1725_n1295), 
	.I(n1295));
   DELDKHD FE_PHC1724_n1459 (.O(FE_PHN1724_n1459), 
	.I(n1459));
   DELDKHD FE_PHC1723_n2097 (.O(FE_PHN1723_n2097), 
	.I(n2097));
   DELDKHD FE_PHC1722_n3450 (.O(FE_PHN1722_n3450), 
	.I(n3450));
   DELDKHD FE_PHC1721_n4476 (.O(FE_PHN1721_n4476), 
	.I(n4476));
   DELDKHD FE_PHC1720_ram_117__6_ (.O(FE_PHN1720_ram_117__6_), 
	.I(\ram[117][6] ));
   DELDKHD FE_PHC1719_n4041 (.O(FE_PHN1719_n4041), 
	.I(n4041));
   DELDKHD FE_PHC1718_n4530 (.O(FE_PHN1718_n4530), 
	.I(n4530));
   DELDKHD FE_PHC1717_n2596 (.O(FE_PHN1717_n2596), 
	.I(n2596));
   DELDKHD FE_PHC1716_n2855 (.O(FE_PHN1716_n2855), 
	.I(n2855));
   DELDKHD FE_PHC1715_n2015 (.O(FE_PHN1715_n2015), 
	.I(n2015));
   DELDKHD FE_PHC1714_n836 (.O(FE_PHN1714_n836), 
	.I(n836));
   DELDKHD FE_PHC1713_n1390 (.O(FE_PHN1713_n1390), 
	.I(n1390));
   DELDKHD FE_PHC1712_n4586 (.O(FE_PHN1712_n4586), 
	.I(n4586));
   DELDKHD FE_PHC1711_n2828 (.O(FE_PHN1711_n2828), 
	.I(n2828));
   DELDKHD FE_PHC1710_n4591 (.O(FE_PHN1710_n4591), 
	.I(n4591));
   DELDKHD FE_PHC1709_n757 (.O(FE_PHN1709_n757), 
	.I(n757));
   DELDKHD FE_PHC1708_n3316 (.O(FE_PHN1708_n3316), 
	.I(n3316));
   DELDKHD FE_PHC1707_n4223 (.O(FE_PHN1707_n4223), 
	.I(n4223));
   DELDKHD FE_PHC1706_n3361 (.O(FE_PHN1706_n3361), 
	.I(n3361));
   DELDKHD FE_PHC1705_n4529 (.O(FE_PHN1705_n4529), 
	.I(n4529));
   DELDKHD FE_PHC1704_n3249 (.O(FE_PHN1704_n3249), 
	.I(n3249));
   DELDKHD FE_PHC1703_n2452 (.O(FE_PHN1703_n2452), 
	.I(n2452));
   DELDKHD FE_PHC1702_n3232 (.O(FE_PHN1702_n3232), 
	.I(n3232));
   DELDKHD FE_PHC1701_n2496 (.O(FE_PHN1701_n2496), 
	.I(n2496));
   DELDKHD FE_PHC1700_n3216 (.O(FE_PHN1700_n3216), 
	.I(n3216));
   DELDKHD FE_PHC1699_n3495 (.O(FE_PHN1699_n3495), 
	.I(n3495));
   DELDKHD FE_PHC1698_n1869 (.O(FE_PHN1698_n1869), 
	.I(n1869));
   DELDKHD FE_PHC1697_n4463 (.O(FE_PHN1697_n4463), 
	.I(n4463));
   DELDKHD FE_PHC1696_n676 (.O(FE_PHN1696_n676), 
	.I(n676));
   DELDKHD FE_PHC1695_n3180 (.O(FE_PHN1695_n3180), 
	.I(n3180));
   DELDKHD FE_PHC1694_n4563 (.O(FE_PHN1694_n4563), 
	.I(n4563));
   DELDKHD FE_PHC1693_n693 (.O(FE_PHN1693_n693), 
	.I(n693));
   DELDKHD FE_PHC1692_n3709 (.O(FE_PHN1692_n3709), 
	.I(n3709));
   DELDKHD FE_PHC1691_n1252 (.O(FE_PHN1691_n1252), 
	.I(n1252));
   DELDKHD FE_PHC1690_n3711 (.O(FE_PHN1690_n3711), 
	.I(n3711));
   DELDKHD FE_PHC1689_n4468 (.O(FE_PHN1689_n4468), 
	.I(n4468));
   DELDKHD FE_PHC1688_n1942 (.O(FE_PHN1688_n1942), 
	.I(n1942));
   DELDKHD FE_PHC1687_n2088 (.O(FE_PHN1687_n2088), 
	.I(n2088));
   DELDKHD FE_PHC1686_n2345 (.O(FE_PHN1686_n2345), 
	.I(n2345));
   DELDKHD FE_PHC1685_n4677 (.O(FE_PHN1685_n4677), 
	.I(n4677));
   DELDKHD FE_PHC1684_n696 (.O(FE_PHN1684_n696), 
	.I(n696));
   DELDKHD FE_PHC1683_n1181 (.O(FE_PHN1683_n1181), 
	.I(n1181));
   DELDKHD FE_PHC1682_n1276 (.O(FE_PHN1682_n1276), 
	.I(n1276));
   DELDKHD FE_PHC1681_n821 (.O(FE_PHN1681_n821), 
	.I(n821));
   DELDKHD FE_PHC1680_n1909 (.O(FE_PHN1680_n1909), 
	.I(n1909));
   DELDKHD FE_PHC1679_n4234 (.O(FE_PHN1679_n4234), 
	.I(n4234));
   DELDKHD FE_PHC1678_n2305 (.O(FE_PHN1678_n2305), 
	.I(n2305));
   DELDKHD FE_PHC1677_n4069 (.O(FE_PHN1677_n4069), 
	.I(n4069));
   DELDKHD FE_PHC1676_n2834 (.O(FE_PHN1676_n2834), 
	.I(n2834));
   DELDKHD FE_PHC1675_n1599 (.O(FE_PHN1675_n1599), 
	.I(n1599));
   DELDKHD FE_PHC1674_n1944 (.O(FE_PHN1674_n1944), 
	.I(n1944));
   DELDKHD FE_PHC1673_n665 (.O(FE_PHN1673_n665), 
	.I(n665));
   DELDKHD FE_PHC1672_n3620 (.O(FE_PHN1672_n3620), 
	.I(n3620));
   DELDKHD FE_PHC1671_n1853 (.O(FE_PHN1671_n1853), 
	.I(n1853));
   DELDKHD FE_PHC1670_n3371 (.O(FE_PHN1670_n3371), 
	.I(n3371));
   DELDKHD FE_PHC1669_n764 (.O(FE_PHN1669_n764), 
	.I(n764));
   DELDKHD FE_PHC1668_n1717 (.O(FE_PHN1668_n1717), 
	.I(n1717));
   DELDKHD FE_PHC1667_n3199 (.O(FE_PHN1667_n3199), 
	.I(n3199));
   DELDKHD FE_PHC1666_n1939 (.O(FE_PHN1666_n1939), 
	.I(n1939));
   DELDKHD FE_PHC1665_n3613 (.O(FE_PHN1665_n3613), 
	.I(n3613));
   DELDKHD FE_PHC1664_n1826 (.O(FE_PHN1664_n1826), 
	.I(n1826));
   DELDKHD FE_PHC1663_n2191 (.O(FE_PHN1663_n2191), 
	.I(n2191));
   DELDKHD FE_PHC1662_n2664 (.O(FE_PHN1662_n2664), 
	.I(n2664));
   DELDKHD FE_PHC1661_n1746 (.O(FE_PHN1661_n1746), 
	.I(n1746));
   DELDKHD FE_PHC1660_n3785 (.O(FE_PHN1660_n3785), 
	.I(n3785));
   DELDKHD FE_PHC1659_n2095 (.O(FE_PHN1659_n2095), 
	.I(n2095));
   DELDKHD FE_PHC1658_n771 (.O(FE_PHN1658_n771), 
	.I(n771));
   DELDKHD FE_PHC1657_n3287 (.O(FE_PHN1657_n3287), 
	.I(n3287));
   DELDKHD FE_PHC1656_n1989 (.O(FE_PHN1656_n1989), 
	.I(n1989));
   DELDKHD FE_PHC1655_n2640 (.O(FE_PHN1655_n2640), 
	.I(n2640));
   DELDKHD FE_PHC1654_n3419 (.O(FE_PHN1654_n3419), 
	.I(n3419));
   DELDKHD FE_PHC1653_n1499 (.O(FE_PHN1653_n1499), 
	.I(n1499));
   DELDKHD FE_PHC1652_n3825 (.O(FE_PHN1652_n3825), 
	.I(n3825));
   DELDKHD FE_PHC1651_n4039 (.O(FE_PHN1651_n4039), 
	.I(n4039));
   DELDKHD FE_PHC1650_n1129 (.O(FE_PHN1650_n1129), 
	.I(n1129));
   DELDKHD FE_PHC1649_n1098 (.O(FE_PHN1649_n1098), 
	.I(n1098));
   DELDKHD FE_PHC1648_n1317 (.O(FE_PHN1648_n1317), 
	.I(n1317));
   DELDKHD FE_PHC1647_n1504 (.O(FE_PHN1647_n1504), 
	.I(n1504));
   DELDKHD FE_PHC1646_n2666 (.O(FE_PHN1646_n2666), 
	.I(n2666));
   DELDKHD FE_PHC1645_n1682 (.O(FE_PHN1645_n1682), 
	.I(n1682));
   DELDKHD FE_PHC1644_n1253 (.O(FE_PHN1644_n1253), 
	.I(n1253));
   DELDKHD FE_PHC1643_n2311 (.O(FE_PHN1643_n2311), 
	.I(n2311));
   DELDKHD FE_PHC1642_n2327 (.O(FE_PHN1642_n2327), 
	.I(n2327));
   DELDKHD FE_PHC1641_n2635 (.O(FE_PHN1641_n2635), 
	.I(n2635));
   DELDKHD FE_PHC1640_n2660 (.O(FE_PHN1640_n2660), 
	.I(n2660));
   DELDKHD FE_PHC1639_n678 (.O(FE_PHN1639_n678), 
	.I(n678));
   DELDKHD FE_PHC1638_n708 (.O(FE_PHN1638_n708), 
	.I(n708));
   DELDKHD FE_PHC1637_n1521 (.O(FE_PHN1637_n1521), 
	.I(n1521));
   DELDKHD FE_PHC1636_n1631 (.O(FE_PHN1636_n1631), 
	.I(n1631));
   DELDKHD FE_PHC1635_n3600 (.O(FE_PHN1635_n3600), 
	.I(n3600));
   DELDKHD FE_PHC1634_n4487 (.O(FE_PHN1634_n4487), 
	.I(n4487));
   DELDKHD FE_PHC1633_n2548 (.O(FE_PHN1633_n2548), 
	.I(n2548));
   DELDKHD FE_PHC1632_n2007 (.O(FE_PHN1632_n2007), 
	.I(n2007));
   DELDKHD FE_PHC1631_n2246 (.O(FE_PHN1631_n2246), 
	.I(n2246));
   DELDKHD FE_PHC1630_n3187 (.O(FE_PHN1630_n3187), 
	.I(n3187));
   DELDKHD FE_PHC1629_n3660 (.O(FE_PHN1629_n3660), 
	.I(n3660));
   DELDKHD FE_PHC1628_n3793 (.O(FE_PHN1628_n3793), 
	.I(n3793));
   DELDKHD FE_PHC1627_n4492 (.O(FE_PHN1627_n4492), 
	.I(n4492));
   DELDKHD FE_PHC1626_n4601 (.O(FE_PHN1626_n4601), 
	.I(n4601));
   DELDKHD FE_PHC1625_n1227 (.O(FE_PHN1625_n1227), 
	.I(n1227));
   DELDKHD FE_PHC1624_n2323 (.O(FE_PHN1624_n2323), 
	.I(n2323));
   DELDKHD FE_PHC1623_n2364 (.O(FE_PHN1623_n2364), 
	.I(n2364));
   DELDKHD FE_PHC1622_n3335 (.O(FE_PHN1622_n3335), 
	.I(n3335));
   DELDKHD FE_PHC1621_n707 (.O(FE_PHN1621_n707), 
	.I(n707));
   DELDKHD FE_PHC1620_n1230 (.O(FE_PHN1620_n1230), 
	.I(n1230));
   DELDKHD FE_PHC1619_n1544 (.O(FE_PHN1619_n1544), 
	.I(n1544));
   DELDKHD FE_PHC1618_n1552 (.O(FE_PHN1618_n1552), 
	.I(n1552));
   DELDKHD FE_PHC1617_n1300 (.O(FE_PHN1617_n1300), 
	.I(n1300));
   DELDKHD FE_PHC1616_n2303 (.O(FE_PHN1616_n2303), 
	.I(n2303));
   DELDKHD FE_PHC1615_n1888 (.O(FE_PHN1615_n1888), 
	.I(n1888));
   DELDKHD FE_PHC1614_n2020 (.O(FE_PHN1614_n2020), 
	.I(n2020));
   DELDKHD FE_PHC1613_n2860 (.O(FE_PHN1613_n2860), 
	.I(n2860));
   DELDKHD FE_PHC1612_n2346 (.O(FE_PHN1612_n2346), 
	.I(n2346));
   DELDKHD FE_PHC1611_n671 (.O(FE_PHN1611_n671), 
	.I(n671));
   DELDKHD FE_PHC1610_n2275 (.O(FE_PHN1610_n2275), 
	.I(n2275));
   DELDKHD FE_PHC1609_n1932 (.O(FE_PHN1609_n1932), 
	.I(n1932));
   DELDKHD FE_PHC1608_n1238 (.O(FE_PHN1608_n1238), 
	.I(n1238));
   DELDKHD FE_PHC1607_n1288 (.O(FE_PHN1607_n1288), 
	.I(n1288));
   DELDKHD FE_PHC1606_n1743 (.O(FE_PHN1606_n1743), 
	.I(n1743));
   DELDKHD FE_PHC1605_n4140 (.O(FE_PHN1605_n4140), 
	.I(n4140));
   DELDKHD FE_PHC1604_n3494 (.O(FE_PHN1604_n3494), 
	.I(n3494));
   DELDKHD FE_PHC1603_n3229 (.O(FE_PHN1603_n3229), 
	.I(n3229));
   DELDKHD FE_PHC1602_n2525 (.O(FE_PHN1602_n2525), 
	.I(n2525));
   DELDKHD FE_PHC1601_n1131 (.O(FE_PHN1601_n1131), 
	.I(n1131));
   DELDKHD FE_PHC1600_n2313 (.O(FE_PHN1600_n2313), 
	.I(n2313));
   DELDKHD FE_PHC1599_n4472 (.O(FE_PHN1599_n4472), 
	.I(n4472));
   DELDKHD FE_PHC1598_n748 (.O(FE_PHN1598_n748), 
	.I(n748));
   DELDKHD FE_PHC1597_n1505 (.O(FE_PHN1597_n1505), 
	.I(n1505));
   DELDKHD FE_PHC1596_n2244 (.O(FE_PHN1596_n2244), 
	.I(n2244));
   DELDKHD FE_PHC1595_n3690 (.O(FE_PHN1595_n3690), 
	.I(n3690));
   DELDKHD FE_PHC1594_n3294 (.O(FE_PHN1594_n3294), 
	.I(n3294));
   DELDKHD FE_PHC1593_n1251 (.O(FE_PHN1593_n1251), 
	.I(n1251));
   DELDKHD FE_PHC1592_n3251 (.O(FE_PHN1592_n3251), 
	.I(n3251));
   DELDKHD FE_PHC1591_n2864 (.O(FE_PHN1591_n2864), 
	.I(n2864));
   DELDKHD FE_PHC1590_n4660 (.O(FE_PHN1590_n4660), 
	.I(n4660));
   DELDKHD FE_PHC1589_n767 (.O(FE_PHN1589_n767), 
	.I(n767));
   DELDKHD FE_PHC1588_n1172 (.O(FE_PHN1588_n1172), 
	.I(n1172));
   DELDKHD FE_PHC1587_n786 (.O(FE_PHN1587_n786), 
	.I(n786));
   DELDKHD FE_PHC1586_n1951 (.O(FE_PHN1586_n1951), 
	.I(n1951));
   DELDKHD FE_PHC1585_n2608 (.O(FE_PHN1585_n2608), 
	.I(n2608));
   DELDKHD FE_PHC1584_n4653 (.O(FE_PHN1584_n4653), 
	.I(n4653));
   DELDKHD FE_PHC1583_n3379 (.O(FE_PHN1583_n3379), 
	.I(n3379));
   DELDKHD FE_PHC1582_n3712 (.O(FE_PHN1582_n3712), 
	.I(n3712));
   DELDKHD FE_PHC1581_n1655 (.O(FE_PHN1581_n1655), 
	.I(n1655));
   DELDKHD FE_PHC1580_n1721 (.O(FE_PHN1580_n1721), 
	.I(n1721));
   DELDKHD FE_PHC1579_n1189 (.O(FE_PHN1579_n1189), 
	.I(n1189));
   DELDKHD FE_PHC1578_n1204 (.O(FE_PHN1578_n1204), 
	.I(n1204));
   DELDKHD FE_PHC1577_n3188 (.O(FE_PHN1577_n3188), 
	.I(n3188));
   DELDKHD FE_PHC1576_n582 (.O(FE_PHN1576_n582), 
	.I(n582));
   DELDKHD FE_PHC1575_n3208 (.O(FE_PHN1575_n3208), 
	.I(n3208));
   DELDKHD FE_PHC1574_n1637 (.O(FE_PHN1574_n1637), 
	.I(n1637));
   DELDKHD FE_PHC1573_n776 (.O(FE_PHN1573_n776), 
	.I(n776));
   DELDKHD FE_PHC1572_n835 (.O(FE_PHN1572_n835), 
	.I(n835));
   DELDKHD FE_PHC1571_n1485 (.O(FE_PHN1571_n1485), 
	.I(n1485));
   DELDKHD FE_PHC1570_n3514 (.O(FE_PHN1570_n3514), 
	.I(n3514));
   DELCKHD FE_PHC1569_n4592 (.O(FE_PHN1569_n4592), 
	.I(n4592));
   DELCKHD FE_PHC1568_n647 (.O(FE_PHN1568_n647), 
	.I(n647));
   DELCKHD FE_PHC1567_n1822 (.O(FE_PHN1567_n1822), 
	.I(n1822));
   DELCKHD FE_PHC1566_n1689 (.O(FE_PHN1566_n1689), 
	.I(n1689));
   DELCKHD FE_PHC1565_n3317 (.O(FE_PHN1565_n3317), 
	.I(n3317));
   DELCKHD FE_PHC1564_n2233 (.O(FE_PHN1564_n2233), 
	.I(n2233));
   DELCKHD FE_PHC1563_n2468 (.O(FE_PHN1563_n2468), 
	.I(n2468));
   DELCKHD FE_PHC1562_n3836 (.O(FE_PHN1562_n3836), 
	.I(n3836));
   DELCKHD FE_PHC1561_n2725 (.O(FE_PHN1561_n2725), 
	.I(n2725));
   DELCKHD FE_PHC1560_n4630 (.O(FE_PHN1560_n4630), 
	.I(n4630));
   DELCKHD FE_PHC1559_n2762 (.O(FE_PHN1559_n2762), 
	.I(n2762));
   DELCKHD FE_PHC1558_n1114 (.O(FE_PHN1558_n1114), 
	.I(n1114));
   DELCKHD FE_PHC1557_n3424 (.O(FE_PHN1557_n3424), 
	.I(n3424));
   DELCKHD FE_PHC1556_n1490 (.O(FE_PHN1556_n1490), 
	.I(n1490));
   DELCKHD FE_PHC1555_n3314 (.O(FE_PHN1555_n3314), 
	.I(n3314));
   DELCKHD FE_PHC1554_n4594 (.O(FE_PHN1554_n4594), 
	.I(n4594));
   DELCKHD FE_PHC1553_n1803 (.O(FE_PHN1553_n1803), 
	.I(n1803));
   DELCKHD FE_PHC1552_n2025 (.O(FE_PHN1552_n2025), 
	.I(n2025));
   DELCKHD FE_PHC1551_n4126 (.O(FE_PHN1551_n4126), 
	.I(n4126));
   DELCKHD FE_PHC1550_n698 (.O(FE_PHN1550_n698), 
	.I(n698));
   DELCKHD FE_PHC1549_n3569 (.O(FE_PHN1549_n3569), 
	.I(n3569));
   DELCKHD FE_PHC1548_n3183 (.O(FE_PHN1548_n3183), 
	.I(n3183));
   DELCKHD FE_PHC1547_n1548 (.O(FE_PHN1547_n1548), 
	.I(n1548));
   DELCKHD FE_PHC1546_n611 (.O(FE_PHN1546_n611), 
	.I(n611));
   DELCKHD FE_PHC1545_n825 (.O(FE_PHN1545_n825), 
	.I(n825));
   DELCKHD FE_PHC1544_n2568 (.O(FE_PHN1544_n2568), 
	.I(n2568));
   DELCKHD FE_PHC1543_n3330 (.O(FE_PHN1543_n3330), 
	.I(n3330));
   DELCKHD FE_PHC1542_n2092 (.O(FE_PHN1542_n2092), 
	.I(n2092));
   DELCKHD FE_PHC1541_n3789 (.O(FE_PHN1541_n3789), 
	.I(n3789));
   DELCKHD FE_PHC1540_n1478 (.O(FE_PHN1540_n1478), 
	.I(n1478));
   DELCKHD FE_PHC1539_n2289 (.O(FE_PHN1539_n2289), 
	.I(n2289));
   DELCKHD FE_PHC1538_n1709 (.O(FE_PHN1538_n1709), 
	.I(n1709));
   DELCKHD FE_PHC1537_n3305 (.O(FE_PHN1537_n3305), 
	.I(n3305));
   DELCKHD FE_PHC1536_n3173 (.O(FE_PHN1536_n3173), 
	.I(n3173));
   DELCKHD FE_PHC1535_n2187 (.O(FE_PHN1535_n2187), 
	.I(n2187));
   DELCKHD FE_PHC1534_n3539 (.O(FE_PHN1534_n3539), 
	.I(n3539));
   DELCKHD FE_PHC1533_n1783 (.O(FE_PHN1533_n1783), 
	.I(n1783));
   DELCKHD FE_PHC1532_n2593 (.O(FE_PHN1532_n2593), 
	.I(n2593));
   DELCKHD FE_PHC1531_n3652 (.O(FE_PHN1531_n3652), 
	.I(n3652));
   DELCKHD FE_PHC1530_n660 (.O(FE_PHN1530_n660), 
	.I(n660));
   DELCKHD FE_PHC1529_n1307 (.O(FE_PHN1529_n1307), 
	.I(n1307));
   DELCKHD FE_PHC1528_n1353 (.O(FE_PHN1528_n1353), 
	.I(n1353));
   DELCKHD FE_PHC1527_n1542 (.O(FE_PHN1527_n1542), 
	.I(n1542));
   DELCKHD FE_PHC1526_n2881 (.O(FE_PHN1526_n2881), 
	.I(n2881));
   DELCKHD FE_PHC1525_n3596 (.O(FE_PHN1525_n3596), 
	.I(n3596));
   DELCKHD FE_PHC1524_n1471 (.O(FE_PHN1524_n1471), 
	.I(n1471));
   DELCKHD FE_PHC1523_n2539 (.O(FE_PHN1523_n2539), 
	.I(n2539));
   DELCKHD FE_PHC1522_n3753 (.O(FE_PHN1522_n3753), 
	.I(n3753));
   DELCKHD FE_PHC1521_n1835 (.O(FE_PHN1521_n1835), 
	.I(n1835));
   DELCKHD FE_PHC1520_n1623 (.O(FE_PHN1520_n1623), 
	.I(n1623));
   DELCKHD FE_PHC1519_n2780 (.O(FE_PHN1519_n2780), 
	.I(n2780));
   DELCKHD FE_PHC1518_n3773 (.O(FE_PHN1518_n3773), 
	.I(n3773));
   DELCKHD FE_PHC1517_n3867 (.O(FE_PHN1517_n3867), 
	.I(n3867));
   DELCKHD FE_PHC1516_n4160 (.O(FE_PHN1516_n4160), 
	.I(n4160));
   DELCKHD FE_PHC1515_n3425 (.O(FE_PHN1515_n3425), 
	.I(n3425));
   DELCKHD FE_PHC1514_n3696 (.O(FE_PHN1514_n3696), 
	.I(n3696));
   DELCKHD FE_PHC1513_n3276 (.O(FE_PHN1513_n3276), 
	.I(n3276));
   DELCKHD FE_PHC1512_n1182 (.O(FE_PHN1512_n1182), 
	.I(n1182));
   DELCKHD FE_PHC1511_n1556 (.O(FE_PHN1511_n1556), 
	.I(n1556));
   DELCKHD FE_PHC1510_n4485 (.O(FE_PHN1510_n4485), 
	.I(n4485));
   DELCKHD FE_PHC1509_n4060 (.O(FE_PHN1509_n4060), 
	.I(n4060));
   DELCKHD FE_PHC1508_n1895 (.O(FE_PHN1508_n1895), 
	.I(n1895));
   DELCKHD FE_PHC1507_n2321 (.O(FE_PHN1507_n2321), 
	.I(n2321));
   DELCKHD FE_PHC1506_n816 (.O(FE_PHN1506_n816), 
	.I(n816));
   DELCKHD FE_PHC1505_n1092 (.O(FE_PHN1505_n1092), 
	.I(n1092));
   DELCKHD FE_PHC1504_n3482 (.O(FE_PHN1504_n3482), 
	.I(n3482));
   DELCKHD FE_PHC1503_n4154 (.O(FE_PHN1503_n4154), 
	.I(n4154));
   DELCKHD FE_PHC1502_n2840 (.O(FE_PHN1502_n2840), 
	.I(n2840));
   DELCKHD FE_PHC1501_n1273 (.O(FE_PHN1501_n1273), 
	.I(n1273));
   DELCKHD FE_PHC1500_n2006 (.O(FE_PHN1500_n2006), 
	.I(n2006));
   DELCKHD FE_PHC1499_n2498 (.O(FE_PHN1499_n2498), 
	.I(n2498));
   DELCKHD FE_PHC1498_n626 (.O(FE_PHN1498_n626), 
	.I(n626));
   DELCKHD FE_PHC1497_n3282 (.O(FE_PHN1497_n3282), 
	.I(n3282));
   DELCKHD FE_PHC1496_n1207 (.O(FE_PHN1496_n1207), 
	.I(n1207));
   DELCKHD FE_PHC1495_n1335 (.O(FE_PHN1495_n1335), 
	.I(n1335));
   DELCKHD FE_PHC1494_n2617 (.O(FE_PHN1494_n2617), 
	.I(n2617));
   DELCKHD FE_PHC1493_n587 (.O(FE_PHN1493_n587), 
	.I(n587));
   DELCKHD FE_PHC1492_n2877 (.O(FE_PHN1492_n2877), 
	.I(n2877));
   DELCKHD FE_PHC1491_n3876 (.O(FE_PHN1491_n3876), 
	.I(n3876));
   DELCKHD FE_PHC1490_n2198 (.O(FE_PHN1490_n2198), 
	.I(n2198));
   DELCKHD FE_PHC1489_n2011 (.O(FE_PHN1489_n2011), 
	.I(n2011));
   DELCKHD FE_PHC1488_n3399 (.O(FE_PHN1488_n3399), 
	.I(n3399));
   DELCKHD FE_PHC1487_n3672 (.O(FE_PHN1487_n3672), 
	.I(n3672));
   DELCKHD FE_PHC1486_n4481 (.O(FE_PHN1486_n4481), 
	.I(n4481));
   DELCKHD FE_PHC1485_n1965 (.O(FE_PHN1485_n1965), 
	.I(n1965));
   DELCKHD FE_PHC1484_n1830 (.O(FE_PHN1484_n1830), 
	.I(n1830));
   DELCKHD FE_PHC1483_n3732 (.O(FE_PHN1483_n3732), 
	.I(n3732));
   DELCKHD FE_PHC1482_n780 (.O(FE_PHN1482_n780), 
	.I(n780));
   DELCKHD FE_PHC1481_n1797 (.O(FE_PHN1481_n1797), 
	.I(n1797));
   DELCKHD FE_PHC1480_n1812 (.O(FE_PHN1480_n1812), 
	.I(n1812));
   DELCKHD FE_PHC1479_n2656 (.O(FE_PHN1479_n2656), 
	.I(n2656));
   DELCKHD FE_PHC1478_n3658 (.O(FE_PHN1478_n3658), 
	.I(n3658));
   DELCKHD FE_PHC1477_n1844 (.O(FE_PHN1477_n1844), 
	.I(n1844));
   DELCKHD FE_PHC1476_n3933 (.O(FE_PHN1476_n3933), 
	.I(n3933));
   DELCKHD FE_PHC1475_n3336 (.O(FE_PHN1475_n3336), 
	.I(n3336));
   DELCKHD FE_PHC1474_n4447 (.O(FE_PHN1474_n4447), 
	.I(n4447));
   DELCKHD FE_PHC1473_n1308 (.O(FE_PHN1473_n1308), 
	.I(n1308));
   DELCKHD FE_PHC1472_n4335 (.O(FE_PHN1472_n4335), 
	.I(n4335));
   DELCKHD FE_PHC1471_n2774 (.O(FE_PHN1471_n2774), 
	.I(n2774));
   DELCKHD FE_PHC1470_ram_122__2_ (.O(FE_PHN1470_ram_122__2_), 
	.I(\ram[122][2] ));
   DELCKHD FE_PHC1469_n1071 (.O(FE_PHN1469_n1071), 
	.I(n1071));
   DELCKHD FE_PHC1468_n2634 (.O(FE_PHN1468_n2634), 
	.I(n2634));
   DELCKHD FE_PHC1467_n1819 (.O(FE_PHN1467_n1819), 
	.I(n1819));
   DELCKHD FE_PHC1466_n3268 (.O(FE_PHN1466_n3268), 
	.I(n3268));
   DELCKHD FE_PHC1465_n3578 (.O(FE_PHN1465_n3578), 
	.I(n3578));
   DELCKHD FE_PHC1464_n3684 (.O(FE_PHN1464_n3684), 
	.I(n3684));
   DELCKHD FE_PHC1463_n1625 (.O(FE_PHN1463_n1625), 
	.I(n1625));
   DELCKHD FE_PHC1462_n2563 (.O(FE_PHN1462_n2563), 
	.I(n2563));
   DELCKHD FE_PHC1461_n1332 (.O(FE_PHN1461_n1332), 
	.I(n1332));
   DELCKHD FE_PHC1460_n4543 (.O(FE_PHN1460_n4543), 
	.I(n4543));
   DELCKHD FE_PHC1459_n1854 (.O(FE_PHN1459_n1854), 
	.I(n1854));
   DELCKHD FE_PHC1458_n3163 (.O(FE_PHN1458_n3163), 
	.I(n3163));
   DELCKHD FE_PHC1457_n2315 (.O(FE_PHN1457_n2315), 
	.I(n2315));
   DELCKHD FE_PHC1456_n4500 (.O(FE_PHN1456_n4500), 
	.I(n4500));
   DELCKHD FE_PHC1455_n614 (.O(FE_PHN1455_n614), 
	.I(n614));
   DELCKHD FE_PHC1454_n788 (.O(FE_PHN1454_n788), 
	.I(n788));
   DELCKHD FE_PHC1453_n2490 (.O(FE_PHN1453_n2490), 
	.I(n2490));
   DELCKHD FE_PHC1452_n2494 (.O(FE_PHN1452_n2494), 
	.I(n2494));
   DELCKHD FE_PHC1451_n2486 (.O(FE_PHN1451_n2486), 
	.I(n2486));
   DELCKHD FE_PHC1450_n3347 (.O(FE_PHN1450_n3347), 
	.I(n3347));
   DELCKHD FE_PHC1449_n3334 (.O(FE_PHN1449_n3334), 
	.I(n3334));
   DELCKHD FE_PHC1448_n2218 (.O(FE_PHN1448_n2218), 
	.I(n2218));
   DELCKHD FE_PHC1447_n2705 (.O(FE_PHN1447_n2705), 
	.I(n2705));
   DELCKHD FE_PHC1446_n3147 (.O(FE_PHN1446_n3147), 
	.I(n3147));
   DELCKHD FE_PHC1445_n3755 (.O(FE_PHN1445_n3755), 
	.I(n3755));
   DELCKHD FE_PHC1444_n1125 (.O(FE_PHN1444_n1125), 
	.I(n1125));
   DELCKHD FE_PHC1443_n3774 (.O(FE_PHN1443_n3774), 
	.I(n3774));
   DELCKHD FE_PHC1442_n1955 (.O(FE_PHN1442_n1955), 
	.I(n1955));
   DELCKHD FE_PHC1441_n3393 (.O(FE_PHN1441_n3393), 
	.I(n3393));
   DELCKHD FE_PHC1440_n4347 (.O(FE_PHN1440_n4347), 
	.I(n4347));
   DELCKHD FE_PHC1439_n2800 (.O(FE_PHN1439_n2800), 
	.I(n2800));
   DELCKHD FE_PHC1438_n3582 (.O(FE_PHN1438_n3582), 
	.I(n3582));
   DELCKHD FE_PHC1437_n3383 (.O(FE_PHN1437_n3383), 
	.I(n3383));
   DELCKHD FE_PHC1436_n3515 (.O(FE_PHN1436_n3515), 
	.I(n3515));
   DELCKHD FE_PHC1435_n3823 (.O(FE_PHN1435_n3823), 
	.I(n3823));
   DELCKHD FE_PHC1434_n4488 (.O(FE_PHN1434_n4488), 
	.I(n4488));
   DELCKHD FE_PHC1433_n1423 (.O(FE_PHN1433_n1423), 
	.I(n1423));
   DELCKHD FE_PHC1432_n712 (.O(FE_PHN1432_n712), 
	.I(n712));
   DELCKHD FE_PHC1431_n1985 (.O(FE_PHN1431_n1985), 
	.I(n1985));
   DELCKHD FE_PHC1430_n2557 (.O(FE_PHN1430_n2557), 
	.I(n2557));
   DELCKHD FE_PHC1429_n2767 (.O(FE_PHN1429_n2767), 
	.I(n2767));
   DELCKHD FE_PHC1428_n3713 (.O(FE_PHN1428_n3713), 
	.I(n3713));
   DELCKHD FE_PHC1427_n3705 (.O(FE_PHN1427_n3705), 
	.I(n3705));
   DELCKHD FE_PHC1426_n2272 (.O(FE_PHN1426_n2272), 
	.I(n2272));
   DELCKHD FE_PHC1425_n4452 (.O(FE_PHN1425_n4452), 
	.I(n4452));
   DELCKHD FE_PHC1424_n1138 (.O(FE_PHN1424_n1138), 
	.I(n1138));
   DELCKHD FE_PHC1423_n3218 (.O(FE_PHN1423_n3218), 
	.I(n3218));
   DELCKHD FE_PHC1422_n1633 (.O(FE_PHN1422_n1633), 
	.I(n1633));
   DELCKHD FE_PHC1421_n3414 (.O(FE_PHN1421_n3414), 
	.I(n3414));
   DELCKHD FE_PHC1420_n995 (.O(FE_PHN1420_n995), 
	.I(n995));
   DELCKHD FE_PHC1419_n3886 (.O(FE_PHN1419_n3886), 
	.I(n3886));
   DELCKHD FE_PHC1418_n1067 (.O(FE_PHN1418_n1067), 
	.I(n1067));
   DELCKHD FE_PHC1417_n826 (.O(FE_PHN1417_n826), 
	.I(n826));
   DELCKHD FE_PHC1416_n1837 (.O(FE_PHN1416_n1837), 
	.I(n1837));
   DELCKHD FE_PHC1415_n3801 (.O(FE_PHN1415_n3801), 
	.I(n3801));
   DELCKHD FE_PHC1414_n730 (.O(FE_PHN1414_n730), 
	.I(n730));
   DELCKHD FE_PHC1413_n3741 (.O(FE_PHN1413_n3741), 
	.I(n3741));
   DELCKHD FE_PHC1412_n2822 (.O(FE_PHN1412_n2822), 
	.I(n2822));
   DELCKHD FE_PHC1411_n3198 (.O(FE_PHN1411_n3198), 
	.I(n3198));
   DELCKHD FE_PHC1410_n4444 (.O(FE_PHN1410_n4444), 
	.I(n4444));
   DELCKHD FE_PHC1409_n1541 (.O(FE_PHN1409_n1541), 
	.I(n1541));
   DELCKHD FE_PHC1408_n1575 (.O(FE_PHN1408_n1575), 
	.I(n1575));
   DELCKHD FE_PHC1407_n1892 (.O(FE_PHN1407_n1892), 
	.I(n1892));
   DELCKHD FE_PHC1406_n3415 (.O(FE_PHN1406_n3415), 
	.I(n3415));
   DELCKHD FE_PHC1405_n4657 (.O(FE_PHN1405_n4657), 
	.I(n4657));
   DELCKHD FE_PHC1404_n2784 (.O(FE_PHN1404_n2784), 
	.I(n2784));
   DELCKHD FE_PHC1403_n3529 (.O(FE_PHN1403_n3529), 
	.I(n3529));
   DELCKHD FE_PHC1402_n2844 (.O(FE_PHN1402_n2844), 
	.I(n2844));
   DELCKHD FE_PHC1401_n1327 (.O(FE_PHN1401_n1327), 
	.I(n1327));
   DELCKHD FE_PHC1400_n790 (.O(FE_PHN1400_n790), 
	.I(n790));
   DELCKHD FE_PHC1399_n774 (.O(FE_PHN1399_n774), 
	.I(n774));
   DELCKHD FE_PHC1398_n624 (.O(FE_PHN1398_n624), 
	.I(n624));
   DELCKHD FE_PHC1397_n2530 (.O(FE_PHN1397_n2530), 
	.I(n2530));
   DELCKHD FE_PHC1396_n1566 (.O(FE_PHN1396_n1566), 
	.I(n1566));
   DELCKHD FE_PHC1395_n4453 (.O(FE_PHN1395_n4453), 
	.I(n4453));
   DELCKHD FE_PHC1394_n1211 (.O(FE_PHN1394_n1211), 
	.I(n1211));
   DELCKHD FE_PHC1393_n2584 (.O(FE_PHN1393_n2584), 
	.I(n2584));
   DELCKHD FE_PHC1392_n3644 (.O(FE_PHN1392_n3644), 
	.I(n3644));
   DELCKHD FE_PHC1391_n1180 (.O(FE_PHN1391_n1180), 
	.I(n1180));
   DELCKHD FE_PHC1390_n4306 (.O(FE_PHN1390_n4306), 
	.I(n4306));
   DELCKHD FE_PHC1389_n4458 (.O(FE_PHN1389_n4458), 
	.I(n4458));
   DELCKHD FE_PHC1388_n1763 (.O(FE_PHN1388_n1763), 
	.I(n1763));
   DELCKHD FE_PHC1387_n1833 (.O(FE_PHN1387_n1833), 
	.I(n1833));
   DELCKHD FE_PHC1386_n3397 (.O(FE_PHN1386_n3397), 
	.I(n3397));
   DELCKHD FE_PHC1385_n765 (.O(FE_PHN1385_n765), 
	.I(n765));
   DELCKHD FE_PHC1384_n3571 (.O(FE_PHN1384_n3571), 
	.I(n3571));
   DELCKHD FE_PHC1383_n4089 (.O(FE_PHN1383_n4089), 
	.I(n4089));
   DELCKHD FE_PHC1382_n4652 (.O(FE_PHN1382_n4652), 
	.I(n4652));
   DELCKHD FE_PHC1381_n3266 (.O(FE_PHN1381_n3266), 
	.I(n3266));
   DELCKHD FE_PHC1380_n3395 (.O(FE_PHN1380_n3395), 
	.I(n3395));
   DELCKHD FE_PHC1379_n1733 (.O(FE_PHN1379_n1733), 
	.I(n1733));
   DELCKHD FE_PHC1378_n1900 (.O(FE_PHN1378_n1900), 
	.I(n1900));
   DELCKHD FE_PHC1377_n2537 (.O(FE_PHN1377_n2537), 
	.I(n2537));
   DELCKHD FE_PHC1376_n4431 (.O(FE_PHN1376_n4431), 
	.I(n4431));
   DELCKHD FE_PHC1375_n4433 (.O(FE_PHN1375_n4433), 
	.I(n4433));
   DELCKHD FE_PHC1374_n1185 (.O(FE_PHN1374_n1185), 
	.I(n1185));
   DELCKHD FE_PHC1373_n1858 (.O(FE_PHN1373_n1858), 
	.I(n1858));
   DELCKHD FE_PHC1372_n2812 (.O(FE_PHN1372_n2812), 
	.I(n2812));
   DELCKHD FE_PHC1371_n3703 (.O(FE_PHN1371_n3703), 
	.I(n3703));
   DELCKHD FE_PHC1370_n3890 (.O(FE_PHN1370_n3890), 
	.I(n3890));
   DELDKHD FE_PHC1369_n2230 (.O(FE_PHN1369_n2230), 
	.I(n2230));
   DELDKHD FE_PHC1368_n4108 (.O(FE_PHN1368_n4108), 
	.I(n4108));
   DELDKHD FE_PHC1367_n3342 (.O(FE_PHN1367_n3342), 
	.I(n3342));
   DELDKHD FE_PHC1366_n3809 (.O(FE_PHN1366_n3809), 
	.I(n3809));
   DELDKHD FE_PHC1365_n1202 (.O(FE_PHN1365_n1202), 
	.I(n1202));
   DELDKHD FE_PHC1364_n1871 (.O(FE_PHN1364_n1871), 
	.I(n1871));
   DELDKHD FE_PHC1363_n3492 (.O(FE_PHN1363_n3492), 
	.I(n3492));
   DELDKHD FE_PHC1362_n3391 (.O(FE_PHN1362_n3391), 
	.I(n3391));
   DELDKHD FE_PHC1361_n2503 (.O(FE_PHN1361_n2503), 
	.I(n2503));
   DELDKHD FE_PHC1360_n2194 (.O(FE_PHN1360_n2194), 
	.I(n2194));
   DELDKHD FE_PHC1359_n3196 (.O(FE_PHN1359_n3196), 
	.I(n3196));
   DELDKHD FE_PHC1358_n3780 (.O(FE_PHN1358_n3780), 
	.I(n3780));
   DELDKHD FE_PHC1357_n1515 (.O(FE_PHN1357_n1515), 
	.I(n1515));
   DELDKHD FE_PHC1356_n3691 (.O(FE_PHN1356_n3691), 
	.I(n3691));
   DELDKHD FE_PHC1355_n2082 (.O(FE_PHN1355_n2082), 
	.I(n2082));
   DELDKHD FE_PHC1354_n3322 (.O(FE_PHN1354_n3322), 
	.I(n3322));
   DELDKHD FE_PHC1353_n4432 (.O(FE_PHN1353_n4432), 
	.I(n4432));
   DELDKHD FE_PHC1352_n1510 (.O(FE_PHN1352_n1510), 
	.I(n1510));
   DELDKHD FE_PHC1351_n1805 (.O(FE_PHN1351_n1805), 
	.I(n1805));
   DELDKHD FE_PHC1350_n4051 (.O(FE_PHN1350_n4051), 
	.I(n4051));
   DELDKHD FE_PHC1349_n1847 (.O(FE_PHN1349_n1847), 
	.I(n1847));
   DELDKHD FE_PHC1348_n2538 (.O(FE_PHN1348_n2538), 
	.I(n2538));
   DELDKHD FE_PHC1347_n1907 (.O(FE_PHN1347_n1907), 
	.I(n1907));
   DELDKHD FE_PHC1346_n3607 (.O(FE_PHN1346_n3607), 
	.I(n3607));
   DELDKHD FE_PHC1345_n3837 (.O(FE_PHN1345_n3837), 
	.I(n3837));
   DELDKHD FE_PHC1344_n2643 (.O(FE_PHN1344_n2643), 
	.I(n2643));
   DELDKHD FE_PHC1343_n1378 (.O(FE_PHN1343_n1378), 
	.I(n1378));
   DELDKHD FE_PHC1342_n3283 (.O(FE_PHN1342_n3283), 
	.I(n3283));
   DELDKHD FE_PHC1341_n3834 (.O(FE_PHN1341_n3834), 
	.I(n3834));
   DELDKHD FE_PHC1340_n2680 (.O(FE_PHN1340_n2680), 
	.I(n2680));
   DELDKHD FE_PHC1339_n2514 (.O(FE_PHN1339_n2514), 
	.I(n2514));
   DELDKHD FE_PHC1338_n1466 (.O(FE_PHN1338_n1466), 
	.I(n1466));
   DELDKHD FE_PHC1337_n3949 (.O(FE_PHN1337_n3949), 
	.I(n3949));
   DELDKHD FE_PHC1336_n4078 (.O(FE_PHN1336_n4078), 
	.I(n4078));
   DELDKHD FE_PHC1335_n2819 (.O(FE_PHN1335_n2819), 
	.I(n2819));
   DELDKHD FE_PHC1334_n4552 (.O(FE_PHN1334_n4552), 
	.I(n4552));
   DELDKHD FE_PHC1333_n3811 (.O(FE_PHN1333_n3811), 
	.I(n3811));
   DELDKHD FE_PHC1332_n1073 (.O(FE_PHN1332_n1073), 
	.I(n1073));
   DELDKHD FE_PHC1331_n3318 (.O(FE_PHN1331_n3318), 
	.I(n3318));
   DELDKHD FE_PHC1330_n1411 (.O(FE_PHN1330_n1411), 
	.I(n1411));
   DELDKHD FE_PHC1329_n697 (.O(FE_PHN1329_n697), 
	.I(n697));
   DELDKHD FE_PHC1328_n1982 (.O(FE_PHN1328_n1982), 
	.I(n1982));
   DELDKHD FE_PHC1327_n1364 (.O(FE_PHN1327_n1364), 
	.I(n1364));
   DELDKHD FE_PHC1326_n2046 (.O(FE_PHN1326_n2046), 
	.I(n2046));
   DELDKHD FE_PHC1325_n2520 (.O(FE_PHN1325_n2520), 
	.I(n2520));
   DELDKHD FE_PHC1324_n2940 (.O(FE_PHN1324_n2940), 
	.I(n2940));
   DELDKHD FE_PHC1323_n4626 (.O(FE_PHN1323_n4626), 
	.I(n4626));
   DELDKHD FE_PHC1322_ram_129__7_ (.O(FE_PHN1322_ram_129__7_), 
	.I(\ram[129][7] ));
   DELDKHD FE_PHC1321_ram_65__8_ (.O(FE_PHN1321_ram_65__8_), 
	.I(\ram[65][8] ));
   DELDKHD FE_PHC1320_n3650 (.O(FE_PHN1320_n3650), 
	.I(n3650));
   DELDKHD FE_PHC1319_n3303 (.O(FE_PHN1319_n3303), 
	.I(n3303));
   DELDKHD FE_PHC1318_ram_81__13_ (.O(FE_PHN1318_ram_81__13_), 
	.I(\ram[81][13] ));
   DELDKHD FE_PHC1317_n679 (.O(FE_PHN1317_n679), 
	.I(n679));
   DELDKHD FE_PHC1316_n605 (.O(FE_PHN1316_n605), 
	.I(n605));
   DELDKHD FE_PHC1315_n3698 (.O(FE_PHN1315_n3698), 
	.I(n3698));
   DELDKHD FE_PHC1314_n3488 (.O(FE_PHN1314_n3488), 
	.I(n3488));
   DELDKHD FE_PHC1313_n1769 (.O(FE_PHN1313_n1769), 
	.I(n1769));
   DELDKHD FE_PHC1312_n2363 (.O(FE_PHN1312_n2363), 
	.I(n2363));
   DELDKHD FE_PHC1311_n1217 (.O(FE_PHN1311_n1217), 
	.I(n1217));
   DELDKHD FE_PHC1310_n1214 (.O(FE_PHN1310_n1214), 
	.I(n1214));
   DELDKHD FE_PHC1309_n3333 (.O(FE_PHN1309_n3333), 
	.I(n3333));
   DELDKHD FE_PHC1308_n1075 (.O(FE_PHN1308_n1075), 
	.I(n1075));
   DELDKHD FE_PHC1307_n1248 (.O(FE_PHN1307_n1248), 
	.I(n1248));
   DELDKHD FE_PHC1306_n3464 (.O(FE_PHN1306_n3464), 
	.I(n3464));
   DELDKHD FE_PHC1305_n798 (.O(FE_PHN1305_n798), 
	.I(n798));
   DELDKHD FE_PHC1304_n1643 (.O(FE_PHN1304_n1643), 
	.I(n1643));
   DELDKHD FE_PHC1303_n4455 (.O(FE_PHN1303_n4455), 
	.I(n4455));
   DELDKHD FE_PHC1302_n4535 (.O(FE_PHN1302_n4535), 
	.I(n4535));
   DELDKHD FE_PHC1301_n2267 (.O(FE_PHN1301_n2267), 
	.I(n2267));
   DELDKHD FE_PHC1300_n3145 (.O(FE_PHN1300_n3145), 
	.I(n3145));
   DELDKHD FE_PHC1299_n2853 (.O(FE_PHN1299_n2853), 
	.I(n2853));
   DELDKHD FE_PHC1298_n3480 (.O(FE_PHN1298_n3480), 
	.I(n3480));
   DELDKHD FE_PHC1297_n3717 (.O(FE_PHN1297_n3717), 
	.I(n3717));
   DELDKHD FE_PHC1296_n1218 (.O(FE_PHN1296_n1218), 
	.I(n1218));
   DELDKHD FE_PHC1295_n2081 (.O(FE_PHN1295_n2081), 
	.I(n2081));
   DELDKHD FE_PHC1294_n3788 (.O(FE_PHN1294_n3788), 
	.I(n3788));
   DELDKHD FE_PHC1293_n4612 (.O(FE_PHN1293_n4612), 
	.I(n4612));
   DELDKHD FE_PHC1292_n3815 (.O(FE_PHN1292_n3815), 
	.I(n3815));
   DELDKHD FE_PHC1291_n1409 (.O(FE_PHN1291_n1409), 
	.I(n1409));
   DELDKHD FE_PHC1290_n2250 (.O(FE_PHN1290_n2250), 
	.I(n2250));
   DELDKHD FE_PHC1289_n3880 (.O(FE_PHN1289_n3880), 
	.I(n3880));
   DELDKHD FE_PHC1288_n659 (.O(FE_PHN1288_n659), 
	.I(n659));
   DELDKHD FE_PHC1287_n1123 (.O(FE_PHN1287_n1123), 
	.I(n1123));
   DELDKHD FE_PHC1286_n1846 (.O(FE_PHN1286_n1846), 
	.I(n1846));
   DELDKHD FE_PHC1285_n3725 (.O(FE_PHN1285_n3725), 
	.I(n3725));
   DELDKHD FE_PHC1284_n3162 (.O(FE_PHN1284_n3162), 
	.I(n3162));
   DELDKHD FE_PHC1283_n1930 (.O(FE_PHN1283_n1930), 
	.I(n1930));
   DELDKHD FE_PHC1282_n2160 (.O(FE_PHN1282_n2160), 
	.I(n2160));
   DELDKHD FE_PHC1281_n4627 (.O(FE_PHN1281_n4627), 
	.I(n4627));
   DELDKHD FE_PHC1280_n4157 (.O(FE_PHN1280_n4157), 
	.I(n4157));
   DELDKHD FE_PHC1279_n3154 (.O(FE_PHN1279_n3154), 
	.I(n3154));
   DELDKHD FE_PHC1278_n4556 (.O(FE_PHN1278_n4556), 
	.I(n4556));
   DELDKHD FE_PHC1277_n1240 (.O(FE_PHN1277_n1240), 
	.I(n1240));
   DELDKHD FE_PHC1276_n4531 (.O(FE_PHN1276_n4531), 
	.I(n4531));
   DELDKHD FE_PHC1275_n1607 (.O(FE_PHN1275_n1607), 
	.I(n1607));
   DELDKHD FE_PHC1274_n827 (.O(FE_PHN1274_n827), 
	.I(n827));
   DELDKHD FE_PHC1273_n1233 (.O(FE_PHN1273_n1233), 
	.I(n1233));
   DELDKHD FE_PHC1272_n1241 (.O(FE_PHN1272_n1241), 
	.I(n1241));
   DELDKHD FE_PHC1271_n1340 (.O(FE_PHN1271_n1340), 
	.I(n1340));
   DELDKHD FE_PHC1270_n1394 (.O(FE_PHN1270_n1394), 
	.I(n1394));
   DELDKHD FE_PHC1269_n1550 (.O(FE_PHN1269_n1550), 
	.I(n1550));
   DELDKHD FE_PHC1268_n4348 (.O(FE_PHN1268_n4348), 
	.I(n4348));
   DELDKHD FE_PHC1267_n4656 (.O(FE_PHN1267_n4656), 
	.I(n4656));
   DELDKHD FE_PHC1266_n2658 (.O(FE_PHN1266_n2658), 
	.I(n2658));
   DELDKHD FE_PHC1265_n2837 (.O(FE_PHN1265_n2837), 
	.I(n2837));
   DELDKHD FE_PHC1264_n810 (.O(FE_PHN1264_n810), 
	.I(n810));
   DELDKHD FE_PHC1263_n2684 (.O(FE_PHN1263_n2684), 
	.I(n2684));
   DELDKHD FE_PHC1262_n2296 (.O(FE_PHN1262_n2296), 
	.I(n2296));
   DELDKHD FE_PHC1261_n3368 (.O(FE_PHN1261_n3368), 
	.I(n3368));
   DELDKHD FE_PHC1260_n3521 (.O(FE_PHN1260_n3521), 
	.I(n3521));
   DELDKHD FE_PHC1259_n3215 (.O(FE_PHN1259_n3215), 
	.I(n3215));
   DELDKHD FE_PHC1258_n4127 (.O(FE_PHN1258_n4127), 
	.I(n4127));
   DELDKHD FE_PHC1257_n1668 (.O(FE_PHN1257_n1668), 
	.I(n1668));
   DELDKHD FE_PHC1256_n4483 (.O(FE_PHN1256_n4483), 
	.I(n4483));
   DELDKHD FE_PHC1255_n3315 (.O(FE_PHN1255_n3315), 
	.I(n3315));
   DELDKHD FE_PHC1254_n1140 (.O(FE_PHN1254_n1140), 
	.I(n1140));
   DELDKHD FE_PHC1253_n2342 (.O(FE_PHN1253_n2342), 
	.I(n2342));
   DELDKHD FE_PHC1252_n2792 (.O(FE_PHN1252_n2792), 
	.I(n2792));
   DELDKHD FE_PHC1251_n1651 (.O(FE_PHN1251_n1651), 
	.I(n1651));
   DELDKHD FE_PHC1250_n4354 (.O(FE_PHN1250_n4354), 
	.I(n4354));
   DELDKHD FE_PHC1249_n1728 (.O(FE_PHN1249_n1728), 
	.I(n1728));
   DELDKHD FE_PHC1248_n4534 (.O(FE_PHN1248_n4534), 
	.I(n4534));
   DELDKHD FE_PHC1247_n4264 (.O(FE_PHN1247_n4264), 
	.I(n4264));
   DELDKHD FE_PHC1246_n4611 (.O(FE_PHN1246_n4611), 
	.I(n4611));
   DELDKHD FE_PHC1245_n2823 (.O(FE_PHN1245_n2823), 
	.I(n2823));
   DELDKHD FE_PHC1244_n2591 (.O(FE_PHN1244_n2591), 
	.I(n2591));
   DELDKHD FE_PHC1243_n2283 (.O(FE_PHN1243_n2283), 
	.I(n2283));
   DELDKHD FE_PHC1242_n1758 (.O(FE_PHN1242_n1758), 
	.I(n1758));
   DELDKHD FE_PHC1241_n4061 (.O(FE_PHN1241_n4061), 
	.I(n4061));
   DELDKHD FE_PHC1240_n1666 (.O(FE_PHN1240_n1666), 
	.I(n1666));
   DELDKHD FE_PHC1239_n2228 (.O(FE_PHN1239_n2228), 
	.I(n2228));
   DELDKHD FE_PHC1238_n2620 (.O(FE_PHN1238_n2620), 
	.I(n2620));
   DELDKHD FE_PHC1237_n3806 (.O(FE_PHN1237_n3806), 
	.I(n3806));
   DELDKHD FE_PHC1236_n1379 (.O(FE_PHN1236_n1379), 
	.I(n1379));
   DELDKHD FE_PHC1235_n1903 (.O(FE_PHN1235_n1903), 
	.I(n1903));
   DELDKHD FE_PHC1234_n2641 (.O(FE_PHN1234_n2641), 
	.I(n2641));
   DELDKHD FE_PHC1233_n2931 (.O(FE_PHN1233_n2931), 
	.I(n2931));
   DELDKHD FE_PHC1232_n2657 (.O(FE_PHN1232_n2657), 
	.I(n2657));
   DELDKHD FE_PHC1231_n3227 (.O(FE_PHN1231_n3227), 
	.I(n3227));
   DELDKHD FE_PHC1230_n805 (.O(FE_PHN1230_n805), 
	.I(n805));
   DELDKHD FE_PHC1229_n2745 (.O(FE_PHN1229_n2745), 
	.I(n2745));
   DELDKHD FE_PHC1228_n3189 (.O(FE_PHN1228_n3189), 
	.I(n3189));
   DELDKHD FE_PHC1227_n2687 (.O(FE_PHN1227_n2687), 
	.I(n2687));
   DELDKHD FE_PHC1226_n1867 (.O(FE_PHN1226_n1867), 
	.I(n1867));
   DELDKHD FE_PHC1225_n2491 (.O(FE_PHN1225_n2491), 
	.I(n2491));
   DELDKHD FE_PHC1224_n2763 (.O(FE_PHN1224_n2763), 
	.I(n2763));
   DELDKHD FE_PHC1223_n683 (.O(FE_PHN1223_n683), 
	.I(n683));
   DELDKHD FE_PHC1222_n1849 (.O(FE_PHN1222_n1849), 
	.I(n1849));
   DELDKHD FE_PHC1221_n1348 (.O(FE_PHN1221_n1348), 
	.I(n1348));
   DELDKHD FE_PHC1220_n2699 (.O(FE_PHN1220_n2699), 
	.I(n2699));
   DELDKHD FE_PHC1219_n2838 (.O(FE_PHN1219_n2838), 
	.I(n2838));
   DELDKHD FE_PHC1218_n4505 (.O(FE_PHN1218_n4505), 
	.I(n4505));
   DELDKHD FE_PHC1217_n3581 (.O(FE_PHN1217_n3581), 
	.I(n3581));
   DELDKHD FE_PHC1216_n3615 (.O(FE_PHN1216_n3615), 
	.I(n3615));
   DELDKHD FE_PHC1215_n3831 (.O(FE_PHN1215_n3831), 
	.I(n3831));
   DELDKHD FE_PHC1214_n4177 (.O(FE_PHN1214_n4177), 
	.I(n4177));
   DELDKHD FE_PHC1213_n2457 (.O(FE_PHN1213_n2457), 
	.I(n2457));
   DELDKHD FE_PHC1212_n4546 (.O(FE_PHN1212_n4546), 
	.I(n4546));
   DELDKHD FE_PHC1211_n3406 (.O(FE_PHN1211_n3406), 
	.I(n3406));
   DELDKHD FE_PHC1210_n3291 (.O(FE_PHN1210_n3291), 
	.I(n3291));
   DELDKHD FE_PHC1209_n4550 (.O(FE_PHN1209_n4550), 
	.I(n4550));
   DELDKHD FE_PHC1208_n2794 (.O(FE_PHN1208_n2794), 
	.I(n2794));
   DELDKHD FE_PHC1207_n1192 (.O(FE_PHN1207_n1192), 
	.I(n1192));
   DELDKHD FE_PHC1206_n2300 (.O(FE_PHN1206_n2300), 
	.I(n2300));
   DELDKHD FE_PHC1205_n1670 (.O(FE_PHN1205_n1670), 
	.I(n1670));
   DELDKHD FE_PHC1204_n3200 (.O(FE_PHN1204_n3200), 
	.I(n3200));
   DELDKHD FE_PHC1203_n3845 (.O(FE_PHN1203_n3845), 
	.I(n3845));
   DELDKHD FE_PHC1202_n1881 (.O(FE_PHN1202_n1881), 
	.I(n1881));
   DELDKHD FE_PHC1201_n3841 (.O(FE_PHN1201_n3841), 
	.I(n3841));
   DELDKHD FE_PHC1200_n1685 (.O(FE_PHN1200_n1685), 
	.I(n1685));
   DELDKHD FE_PHC1199_n3583 (.O(FE_PHN1199_n3583), 
	.I(n3583));
   DELDKHD FE_PHC1198_n3161 (.O(FE_PHN1198_n3161), 
	.I(n3161));
   DELDKHD FE_PHC1197_n2644 (.O(FE_PHN1197_n2644), 
	.I(n2644));
   DELDKHD FE_PHC1196_n1385 (.O(FE_PHN1196_n1385), 
	.I(n1385));
   DELDKHD FE_PHC1195_n3264 (.O(FE_PHN1195_n3264), 
	.I(n3264));
   DELDKHD FE_PHC1194_n1953 (.O(FE_PHN1194_n1953), 
	.I(n1953));
   DELDKHD FE_PHC1193_n2862 (.O(FE_PHN1193_n2862), 
	.I(n2862));
   DELDKHD FE_PHC1192_n2579 (.O(FE_PHN1192_n2579), 
	.I(n2579));
   DELDKHD FE_PHC1191_n1862 (.O(FE_PHN1191_n1862), 
	.I(n1862));
   DELDKHD FE_PHC1190_n2679 (.O(FE_PHN1190_n2679), 
	.I(n2679));
   DELDKHD FE_PHC1189_n2831 (.O(FE_PHN1189_n2831), 
	.I(n2831));
   DELDKHD FE_PHC1188_n2677 (.O(FE_PHN1188_n2677), 
	.I(n2677));
   DELDKHD FE_PHC1187_n3398 (.O(FE_PHN1187_n3398), 
	.I(n3398));
   DELDKHD FE_PHC1186_n1231 (.O(FE_PHN1186_n1231), 
	.I(n1231));
   DELCKHD FE_PHC1185_n1371 (.O(FE_PHN1185_n1371), 
	.I(n1371));
   DELCKHD FE_PHC1184_n4617 (.O(FE_PHN1184_n4617), 
	.I(n4617));
   DELCKHD FE_PHC1183_n963 (.O(FE_PHN1183_n963), 
	.I(n963));
   DELCKHD FE_PHC1182_n2777 (.O(FE_PHN1182_n2777), 
	.I(n2777));
   DELCKHD FE_PHC1181_n2018 (.O(FE_PHN1181_n2018), 
	.I(n2018));
   DELCKHD FE_PHC1180_n2724 (.O(FE_PHN1180_n2724), 
	.I(n2724));
   DELCKHD FE_PHC1179_n3851 (.O(FE_PHN1179_n3851), 
	.I(n3851));
   DELCKHD FE_PHC1178_n2190 (.O(FE_PHN1178_n2190), 
	.I(n2190));
   DELCKHD FE_PHC1177_n3636 (.O(FE_PHN1177_n3636), 
	.I(n3636));
   DELCKHD FE_PHC1176_n3299 (.O(FE_PHN1176_n3299), 
	.I(n3299));
   DELCKHD FE_PHC1175_n3873 (.O(FE_PHN1175_n3873), 
	.I(n3873));
   DELCKHD FE_PHC1174_n3859 (.O(FE_PHN1174_n3859), 
	.I(n3859));
   DELCKHD FE_PHC1173_n2308 (.O(FE_PHN1173_n2308), 
	.I(n2308));
   DELCKHD FE_PHC1172_n2524 (.O(FE_PHN1172_n2524), 
	.I(n2524));
   DELCKHD FE_PHC1171_n3197 (.O(FE_PHN1171_n3197), 
	.I(n3197));
   DELCKHD FE_PHC1170_n1603 (.O(FE_PHN1170_n1603), 
	.I(n1603));
   DELCKHD FE_PHC1169_n2567 (.O(FE_PHN1169_n2567), 
	.I(n2567));
   DELCKHD FE_PHC1168_n1698 (.O(FE_PHN1168_n1698), 
	.I(n1698));
   DELCKHD FE_PHC1167_n3728 (.O(FE_PHN1167_n3728), 
	.I(n3728));
   DELCKHD FE_PHC1166_n3899 (.O(FE_PHN1166_n3899), 
	.I(n3899));
   DELCKHD FE_PHC1165_n833 (.O(FE_PHN1165_n833), 
	.I(n833));
   DELCKHD FE_PHC1164_n3566 (.O(FE_PHN1164_n3566), 
	.I(n3566));
   DELCKHD FE_PHC1163_n3752 (.O(FE_PHN1163_n3752), 
	.I(n3752));
   DELCKHD FE_PHC1162_n1840 (.O(FE_PHN1162_n1840), 
	.I(n1840));
   DELCKHD FE_PHC1161_n2825 (.O(FE_PHN1161_n2825), 
	.I(n2825));
   DELCKHD FE_PHC1160_n3821 (.O(FE_PHN1160_n3821), 
	.I(n3821));
   DELCKHD FE_PHC1159_n3340 (.O(FE_PHN1159_n3340), 
	.I(n3340));
   DELCKHD FE_PHC1158_n2833 (.O(FE_PHN1158_n2833), 
	.I(n2833));
   DELCKHD FE_PHC1157_n3813 (.O(FE_PHN1157_n3813), 
	.I(n3813));
   DELCKHD FE_PHC1156_n4470 (.O(FE_PHN1156_n4470), 
	.I(n4470));
   DELCKHD FE_PHC1155_n3304 (.O(FE_PHN1155_n3304), 
	.I(n3304));
   DELCKHD FE_PHC1154_n3325 (.O(FE_PHN1154_n3325), 
	.I(n3325));
   DELCKHD FE_PHC1153_n3411 (.O(FE_PHN1153_n3411), 
	.I(n3411));
   DELCKHD FE_PHC1152_n2685 (.O(FE_PHN1152_n2685), 
	.I(n2685));
   DELCKHD FE_PHC1151_n3802 (.O(FE_PHN1151_n3802), 
	.I(n3802));
   DELCKHD FE_PHC1150_n1732 (.O(FE_PHN1150_n1732), 
	.I(n1732));
   DELCKHD FE_PHC1149_n2231 (.O(FE_PHN1149_n2231), 
	.I(n2231));
   DELCKHD FE_PHC1148_n1196 (.O(FE_PHN1148_n1196), 
	.I(n1196));
   DELCKHD FE_PHC1147_n3808 (.O(FE_PHN1147_n3808), 
	.I(n3808));
   DELCKHD FE_PHC1146_n1370 (.O(FE_PHN1146_n1370), 
	.I(n1370));
   DELCKHD FE_PHC1145_n3766 (.O(FE_PHN1145_n3766), 
	.I(n3766));
   DELCKHD FE_PHC1144_n1084 (.O(FE_PHN1144_n1084), 
	.I(n1084));
   DELCKHD FE_PHC1143_n3820 (.O(FE_PHN1143_n3820), 
	.I(n3820));
   DELCKHD FE_PHC1142_n1588 (.O(FE_PHN1142_n1588), 
	.I(n1588));
   DELCKHD FE_PHC1141_n4607 (.O(FE_PHN1141_n4607), 
	.I(n4607));
   DELCKHD FE_PHC1140_n2325 (.O(FE_PHN1140_n2325), 
	.I(n2325));
   DELCKHD FE_PHC1139_n2816 (.O(FE_PHN1139_n2816), 
	.I(n2816));
   DELCKHD FE_PHC1138_n2472 (.O(FE_PHN1138_n2472), 
	.I(n2472));
   DELCKHD FE_PHC1137_n1581 (.O(FE_PHN1137_n1581), 
	.I(n1581));
   DELCKHD FE_PHC1136_n3214 (.O(FE_PHN1136_n3214), 
	.I(n3214));
   DELCKHD FE_PHC1135_n2791 (.O(FE_PHN1135_n2791), 
	.I(n2791));
   DELCKHD FE_PHC1134_n4673 (.O(FE_PHN1134_n4673), 
	.I(n4673));
   DELCKHD FE_PHC1133_n4511 (.O(FE_PHN1133_n4511), 
	.I(n4511));
   DELCKHD FE_PHC1132_n3346 (.O(FE_PHN1132_n3346), 
	.I(n3346));
   DELCKHD FE_PHC1131_n3835 (.O(FE_PHN1131_n3835), 
	.I(n3835));
   DELCKHD FE_PHC1130_n2738 (.O(FE_PHN1130_n2738), 
	.I(n2738));
   DELCKHD FE_PHC1129_n3687 (.O(FE_PHN1129_n3687), 
	.I(n3687));
   DELCKHD FE_PHC1128_n2442 (.O(FE_PHN1128_n2442), 
	.I(n2442));
   DELCKHD FE_PHC1127_n2072 (.O(FE_PHN1127_n2072), 
	.I(n2072));
   DELCKHD FE_PHC1126_n1877 (.O(FE_PHN1126_n1877), 
	.I(n1877));
   DELCKHD FE_PHC1125_n1563 (.O(FE_PHN1125_n1563), 
	.I(n1563));
   DELCKHD FE_PHC1124_n1661 (.O(FE_PHN1124_n1661), 
	.I(n1661));
   DELCKHD FE_PHC1123_n2681 (.O(FE_PHN1123_n2681), 
	.I(n2681));
   DELCKHD FE_PHC1122_n4133 (.O(FE_PHN1122_n4133), 
	.I(n4133));
   DELCKHD FE_PHC1121_n3874 (.O(FE_PHN1121_n3874), 
	.I(n3874));
   DELCKHD FE_PHC1120_n1673 (.O(FE_PHN1120_n1673), 
	.I(n1673));
   DELCKHD FE_PHC1119_n3057 (.O(FE_PHN1119_n3057), 
	.I(n3057));
   DELCKHD FE_PHC1118_n3192 (.O(FE_PHN1118_n3192), 
	.I(n3192));
   DELCKHD FE_PHC1117_n1387 (.O(FE_PHN1117_n1387), 
	.I(n1387));
   DELCKHD FE_PHC1116_n1503 (.O(FE_PHN1116_n1503), 
	.I(n1503));
   DELCKHD FE_PHC1115_n1621 (.O(FE_PHN1115_n1621), 
	.I(n1621));
   DELCKHD FE_PHC1114_n1558 (.O(FE_PHN1114_n1558), 
	.I(n1558));
   DELCKHD FE_PHC1113_n672 (.O(FE_PHN1113_n672), 
	.I(n672));
   DELCKHD FE_PHC1112_n1976 (.O(FE_PHN1112_n1976), 
	.I(n1976));
   DELCKHD FE_PHC1111_n2704 (.O(FE_PHN1111_n2704), 
	.I(n2704));
   DELCKHD FE_PHC1110_n3595 (.O(FE_PHN1110_n3595), 
	.I(n3595));
   DELCKHD FE_PHC1109_n1949 (.O(FE_PHN1109_n1949), 
	.I(n1949));
   DELCKHD FE_PHC1108_n3228 (.O(FE_PHN1108_n3228), 
	.I(n3228));
   DELCKHD FE_PHC1107_n1554 (.O(FE_PHN1107_n1554), 
	.I(n1554));
   DELCKHD FE_PHC1106_n1910 (.O(FE_PHN1106_n1910), 
	.I(n1910));
   DELCKHD FE_PHC1105_n2188 (.O(FE_PHN1105_n2188), 
	.I(n2188));
   DELCKHD FE_PHC1104_n2858 (.O(FE_PHN1104_n2858), 
	.I(n2858));
   DELCKHD FE_PHC1103_n4250 (.O(FE_PHN1103_n4250), 
	.I(n4250));
   DELCKHD FE_PHC1102_n3045 (.O(FE_PHN1102_n3045), 
	.I(n3045));
   DELCKHD FE_PHC1101_n1386 (.O(FE_PHN1101_n1386), 
	.I(n1386));
   DELCKHD FE_PHC1100_n2807 (.O(FE_PHN1100_n2807), 
	.I(n2807));
   DELCKHD FE_PHC1099_n4124 (.O(FE_PHN1099_n4124), 
	.I(n4124));
   DELCKHD FE_PHC1098_n3279 (.O(FE_PHN1098_n3279), 
	.I(n3279));
   DELCKHD FE_PHC1097_n1245 (.O(FE_PHN1097_n1245), 
	.I(n1245));
   DELCKHD FE_PHC1096_n3623 (.O(FE_PHN1096_n3623), 
	.I(n3623));
   DELCKHD FE_PHC1095_n2713 (.O(FE_PHN1095_n2713), 
	.I(n2713));
   DELCKHD FE_PHC1094_n3373 (.O(FE_PHN1094_n3373), 
	.I(n3373));
   DELCKHD FE_PHC1093_n3588 (.O(FE_PHN1093_n3588), 
	.I(n3588));
   DELCKHD FE_PHC1092_n2070 (.O(FE_PHN1092_n2070), 
	.I(n2070));
   DELCKHD FE_PHC1091_n2193 (.O(FE_PHN1091_n2193), 
	.I(n2193));
   DELCKHD FE_PHC1090_n2481 (.O(FE_PHN1090_n2481), 
	.I(n2481));
   DELCKHD FE_PHC1089_n3348 (.O(FE_PHN1089_n3348), 
	.I(n3348));
   DELCKHD FE_PHC1088_n4445 (.O(FE_PHN1088_n4445), 
	.I(n4445));
   DELCKHD FE_PHC1087_n4593 (.O(FE_PHN1087_n4593), 
	.I(n4593));
   DELCKHD FE_PHC1086_n2195 (.O(FE_PHN1086_n2195), 
	.I(n2195));
   DELCKHD FE_PHC1085_n3039 (.O(FE_PHN1085_n3039), 
	.I(n3039));
   DELCKHD FE_PHC1084_n1130 (.O(FE_PHN1084_n1130), 
	.I(n1130));
   DELCKHD FE_PHC1083_n1444 (.O(FE_PHN1083_n1444), 
	.I(n1444));
   DELCKHD FE_PHC1082_n908 (.O(FE_PHN1082_n908), 
	.I(n908));
   DELCKHD FE_PHC1081_n1500 (.O(FE_PHN1081_n1500), 
	.I(n1500));
   DELCKHD FE_PHC1080_n2785 (.O(FE_PHN1080_n2785), 
	.I(n2785));
   DELCKHD FE_PHC1079_n1113 (.O(FE_PHN1079_n1113), 
	.I(n1113));
   DELCKHD FE_PHC1078_n3758 (.O(FE_PHN1078_n3758), 
	.I(n3758));
   DELCKHD FE_PHC1077_n4666 (.O(FE_PHN1077_n4666), 
	.I(n4666));
   DELCKHD FE_PHC1076_n2226 (.O(FE_PHN1076_n2226), 
	.I(n2226));
   DELCKHD FE_PHC1075_n2924 (.O(FE_PHN1075_n2924), 
	.I(n2924));
   DELCKHD FE_PHC1074_n1360 (.O(FE_PHN1074_n1360), 
	.I(n1360));
   DELCKHD FE_PHC1073_n1923 (.O(FE_PHN1073_n1923), 
	.I(n1923));
   DELCKHD FE_PHC1072_n2682 (.O(FE_PHN1072_n2682), 
	.I(n2682));
   DELCKHD FE_PHC1071_n1260 (.O(FE_PHN1071_n1260), 
	.I(n1260));
   DELCKHD FE_PHC1070_n1522 (.O(FE_PHN1070_n1522), 
	.I(n1522));
   DELCKHD FE_PHC1069_n1742 (.O(FE_PHN1069_n1742), 
	.I(n1742));
   DELCKHD FE_PHC1068_n2189 (.O(FE_PHN1068_n2189), 
	.I(n2189));
   DELCKHD FE_PHC1067_n3604 (.O(FE_PHN1067_n3604), 
	.I(n3604));
   DELCKHD FE_PHC1066_n607 (.O(FE_PHN1066_n607), 
	.I(n607));
   DELCKHD FE_PHC1065_n4537 (.O(FE_PHN1065_n4537), 
	.I(n4537));
   DELCKHD FE_PHC1064_n784 (.O(FE_PHN1064_n784), 
	.I(n784));
   DELCKHD FE_PHC1063_n1102 (.O(FE_PHN1063_n1102), 
	.I(n1102));
   DELCKHD FE_PHC1062_n3721 (.O(FE_PHN1062_n3721), 
	.I(n3721));
   DELCKHD FE_PHC1061_n4588 (.O(FE_PHN1061_n4588), 
	.I(n4588));
   DELCKHD FE_PHC1060_n4598 (.O(FE_PHN1060_n4598), 
	.I(n4598));
   DELCKHD FE_PHC1059_n689 (.O(FE_PHN1059_n689), 
	.I(n689));
   DELCKHD FE_PHC1058_ram_201__5_ (.O(FE_PHN1058_ram_201__5_), 
	.I(\ram[201][5] ));
   DELCKHD FE_PHC1057_n4427 (.O(FE_PHN1057_n4427), 
	.I(n4427));
   DELCKHD FE_PHC1056_n4322 (.O(FE_PHN1056_n4322), 
	.I(n4322));
   DELCKHD FE_PHC1055_n2917 (.O(FE_PHN1055_n2917), 
	.I(n2917));
   DELCKHD FE_PHC1054_n1785 (.O(FE_PHN1054_n1785), 
	.I(n1785));
   DELCKHD FE_PHC1053_n2027 (.O(FE_PHN1053_n2027), 
	.I(n2027));
   DELCKHD FE_PHC1052_n4197 (.O(FE_PHN1052_n4197), 
	.I(n4197));
   DELCKHD FE_PHC1051_n618 (.O(FE_PHN1051_n618), 
	.I(n618));
   DELCKHD FE_PHC1050_n3814 (.O(FE_PHN1050_n3814), 
	.I(n3814));
   DELCKHD FE_PHC1049_n4048 (.O(FE_PHN1049_n4048), 
	.I(n4048));
   DELCKHD FE_PHC1048_n3706 (.O(FE_PHN1048_n3706), 
	.I(n3706));
   DELCKHD FE_PHC1047_n3155 (.O(FE_PHN1047_n3155), 
	.I(n3155));
   DELCKHD FE_PHC1046_n663 (.O(FE_PHN1046_n663), 
	.I(n663));
   DELCKHD FE_PHC1045_n615 (.O(FE_PHN1045_n615), 
	.I(n615));
   DELCKHD FE_PHC1044_n4040 (.O(FE_PHN1044_n4040), 
	.I(n4040));
   DELCKHD FE_PHC1043_n926 (.O(FE_PHN1043_n926), 
	.I(n926));
   DELCKHD FE_PHC1042_n1855 (.O(FE_PHN1042_n1855), 
	.I(n1855));
   DELCKHD FE_PHC1041_n2493 (.O(FE_PHN1041_n2493), 
	.I(n2493));
   DELCKHD FE_PHC1040_n3339 (.O(FE_PHN1040_n3339), 
	.I(n3339));
   DELCKHD FE_PHC1039_n2474 (.O(FE_PHN1039_n2474), 
	.I(n2474));
   DELCKHD FE_PHC1038_n3403 (.O(FE_PHN1038_n3403), 
	.I(n3403));
   DELCKHD FE_PHC1037_n3396 (.O(FE_PHN1037_n3396), 
	.I(n3396));
   DELCKHD FE_PHC1036_n4499 (.O(FE_PHN1036_n4499), 
	.I(n4499));
   DELCKHD FE_PHC1035_n1824 (.O(FE_PHN1035_n1824), 
	.I(n1824));
   DELCKHD FE_PHC1034_n2649 (.O(FE_PHN1034_n2649), 
	.I(n2649));
   DELCKHD FE_PHC1033_n3449 (.O(FE_PHN1033_n3449), 
	.I(n3449));
   DELCKHD FE_PHC1032_n4088 (.O(FE_PHN1032_n4088), 
	.I(n4088));
   DELCKHD FE_PHC1031_n4086 (.O(FE_PHN1031_n4086), 
	.I(n4086));
   DELCKHD FE_PHC1030_n4478 (.O(FE_PHN1030_n4478), 
	.I(n4478));
   DELCKHD FE_PHC1029_n4429 (.O(FE_PHN1029_n4429), 
	.I(n4429));
   DELCKHD FE_PHC1028_n2416 (.O(FE_PHN1028_n2416), 
	.I(n2416));
   DELCKHD FE_PHC1027_n2526 (.O(FE_PHN1027_n2526), 
	.I(n2526));
   DELCKHD FE_PHC1026_n823 (.O(FE_PHN1026_n823), 
	.I(n823));
   DELCKHD FE_PHC1025_n1843 (.O(FE_PHN1025_n1843), 
	.I(n1843));
   DELCKHD FE_PHC1024_n2075 (.O(FE_PHN1024_n2075), 
	.I(n2075));
   DELCKHD FE_PHC1023_n2213 (.O(FE_PHN1023_n2213), 
	.I(n2213));
   DELCKHD FE_PHC1022_n2387 (.O(FE_PHN1022_n2387), 
	.I(n2387));
   DELCKHD FE_PHC1021_n4067 (.O(FE_PHN1021_n4067), 
	.I(n4067));
   DELCKHD FE_PHC1020_n4112 (.O(FE_PHN1020_n4112), 
	.I(n4112));
   DELCKHD FE_PHC1019_n1384 (.O(FE_PHN1019_n1384), 
	.I(n1384));
   DELDKHD FE_PHC1018_n1628 (.O(FE_PHN1018_n1628), 
	.I(n1628));
   DELDKHD FE_PHC1017_n3681 (.O(FE_PHN1017_n3681), 
	.I(n3681));
   DELDKHD FE_PHC1016_n1718 (.O(FE_PHN1016_n1718), 
	.I(n1718));
   DELDKHD FE_PHC1015_n2851 (.O(FE_PHN1015_n2851), 
	.I(n2851));
   DELDKHD FE_PHC1014_n2477 (.O(FE_PHN1014_n2477), 
	.I(n2477));
   DELDKHD FE_PHC1013_n3740 (.O(FE_PHN1013_n3740), 
	.I(n3740));
   DELDKHD FE_PHC1012_n4672 (.O(FE_PHN1012_n4672), 
	.I(n4672));
   DELDKHD FE_PHC1011_n1507 (.O(FE_PHN1011_n1507), 
	.I(n1507));
   DELDKHD FE_PHC1010_n1943 (.O(FE_PHN1010_n1943), 
	.I(n1943));
   DELDKHD FE_PHC1009_n4071 (.O(FE_PHN1009_n4071), 
	.I(n4071));
   DELDKHD FE_PHC1008_n617 (.O(FE_PHN1008_n617), 
	.I(n617));
   DELDKHD FE_PHC1007_n1432 (.O(FE_PHN1007_n1432), 
	.I(n1432));
   DELDKHD FE_PHC1006_n2192 (.O(FE_PHN1006_n2192), 
	.I(n2192));
   DELDKHD FE_PHC1005_n1442 (.O(FE_PHN1005_n1442), 
	.I(n1442));
   DELDKHD FE_PHC1004_n3273 (.O(FE_PHN1004_n3273), 
	.I(n3273));
   DELDKHD FE_PHC1003_n2019 (.O(FE_PHN1003_n2019), 
	.I(n2019));
   DELDKHD FE_PHC1002_n3326 (.O(FE_PHN1002_n3326), 
	.I(n3326));
   DELDKHD FE_PHC1001_n1893 (.O(FE_PHN1001_n1893), 
	.I(n1893));
   DELDKHD FE_PHC1000_n3646 (.O(FE_PHN1000_n3646), 
	.I(n3646));
   DELDKHD FE_PHC999_n4616 (.O(FE_PHN999_n4616), 
	.I(n4616));
   DELDKHD FE_PHC998_n1809 (.O(FE_PHN998_n1809), 
	.I(n1809));
   DELDKHD FE_PHC997_n2846 (.O(FE_PHN997_n2846), 
	.I(n2846));
   DELDKHD FE_PHC996_n4486 (.O(FE_PHN996_n4486), 
	.I(n4486));
   DELDKHD FE_PHC995_n1832 (.O(FE_PHN995_n1832), 
	.I(n1832));
   DELDKHD FE_PHC994_n3384 (.O(FE_PHN994_n3384), 
	.I(n3384));
   DELDKHD FE_PHC993_n3794 (.O(FE_PHN993_n3794), 
	.I(n3794));
   DELDKHD FE_PHC992_n1669 (.O(FE_PHN992_n1669), 
	.I(n1669));
   DELDKHD FE_PHC991_n4646 (.O(FE_PHN991_n4646), 
	.I(n4646));
   DELDKHD FE_PHC990_n1528 (.O(FE_PHN990_n1528), 
	.I(n1528));
   DELDKHD FE_PHC989_n3553 (.O(FE_PHN989_n3553), 
	.I(n3553));
   DELDKHD FE_PHC988_n3865 (.O(FE_PHN988_n3865), 
	.I(n3865));
   DELDKHD FE_PHC987_n3726 (.O(FE_PHN987_n3726), 
	.I(n3726));
   DELDKHD FE_PHC986_n2332 (.O(FE_PHN986_n2332), 
	.I(n2332));
   DELDKHD FE_PHC985_n1124 (.O(FE_PHN985_n1124), 
	.I(n1124));
   DELDKHD FE_PHC984_n1506 (.O(FE_PHN984_n1506), 
	.I(n1506));
   DELDKHD FE_PHC983_n1980 (.O(FE_PHN983_n1980), 
	.I(n1980));
   DELDKHD FE_PHC982_n694 (.O(FE_PHN982_n694), 
	.I(n694));
   DELDKHD FE_PHC981_n1408 (.O(FE_PHN981_n1408), 
	.I(n1408));
   DELDKHD FE_PHC980_n2042 (.O(FE_PHN980_n2042), 
	.I(n2042));
   DELDKHD FE_PHC979_n2836 (.O(FE_PHN979_n2836), 
	.I(n2836));
   DELDKHD FE_PHC978_n1351 (.O(FE_PHN978_n1351), 
	.I(n1351));
   DELDKHD FE_PHC977_n4053 (.O(FE_PHN977_n4053), 
	.I(n4053));
   DELDKHD FE_PHC976_n4063 (.O(FE_PHN976_n4063), 
	.I(n4063));
   DELDKHD FE_PHC975_n2856 (.O(FE_PHN975_n2856), 
	.I(n2856));
   DELDKHD FE_PHC974_n2866 (.O(FE_PHN974_n2866), 
	.I(n2866));
   DELDKHD FE_PHC973_n4664 (.O(FE_PHN973_n4664), 
	.I(n4664));
   DELDKHD FE_PHC972_n2440 (.O(FE_PHN972_n2440), 
	.I(n2440));
   DELDKHD FE_PHC971_n2775 (.O(FE_PHN971_n2775), 
	.I(n2775));
   DELDKHD FE_PHC970_n2243 (.O(FE_PHN970_n2243), 
	.I(n2243));
   DELDKHD FE_PHC969_n662 (.O(FE_PHN969_n662), 
	.I(n662));
   DELDKHD FE_PHC968_n1645 (.O(FE_PHN968_n1645), 
	.I(n1645));
   DELDKHD FE_PHC967_n1329 (.O(FE_PHN967_n1329), 
	.I(n1329));
   DELDKHD FE_PHC966_n1081 (.O(FE_PHN966_n1081), 
	.I(n1081));
   DELDKHD FE_PHC965_n3883 (.O(FE_PHN965_n3883), 
	.I(n3883));
   DELDKHD FE_PHC964_n2736 (.O(FE_PHN964_n2736), 
	.I(n2736));
   DELDKHD FE_PHC963_n3589 (.O(FE_PHN963_n3589), 
	.I(n3589));
   DELDKHD FE_PHC962_n2077 (.O(FE_PHN962_n2077), 
	.I(n2077));
   DELDKHD FE_PHC961_n4450 (.O(FE_PHN961_n4450), 
	.I(n4450));
   DELDKHD FE_PHC960_n3505 (.O(FE_PHN960_n3505), 
	.I(n3505));
   DELDKHD FE_PHC959_n1126 (.O(FE_PHN959_n1126), 
	.I(n1126));
   DELDKHD FE_PHC958_n4676 (.O(FE_PHN958_n4676), 
	.I(n4676));
   DELDKHD FE_PHC957_n3441 (.O(FE_PHN957_n3441), 
	.I(n3441));
   DELDKHD FE_PHC956_n1450 (.O(FE_PHN956_n1450), 
	.I(n1450));
   DELDKHD FE_PHC955_n3839 (.O(FE_PHN955_n3839), 
	.I(n3839));
   DELDKHD FE_PHC954_n4272 (.O(FE_PHN954_n4272), 
	.I(n4272));
   DELDKHD FE_PHC953_n4524 (.O(FE_PHN953_n4524), 
	.I(n4524));
   DELDKHD FE_PHC952_n3822 (.O(FE_PHN952_n3822), 
	.I(n3822));
   DELDKHD FE_PHC951_n1565 (.O(FE_PHN951_n1565), 
	.I(n1565));
   DELDKHD FE_PHC950_n1851 (.O(FE_PHN950_n1851), 
	.I(n1851));
   DELDKHD FE_PHC949_n2533 (.O(FE_PHN949_n2533), 
	.I(n2533));
   DELDKHD FE_PHC948_n3195 (.O(FE_PHN948_n3195), 
	.I(n3195));
   DELDKHD FE_PHC947_n4624 (.O(FE_PHN947_n4624), 
	.I(n4624));
   DELDKHD FE_PHC946_n2454 (.O(FE_PHN946_n2454), 
	.I(n2454));
   DELDKHD FE_PHC945_n3254 (.O(FE_PHN945_n3254), 
	.I(n3254));
   DELDKHD FE_PHC944_n3289 (.O(FE_PHN944_n3289), 
	.I(n3289));
   DELDKHD FE_PHC943_n4641 (.O(FE_PHN943_n4641), 
	.I(n4641));
   DELDKHD FE_PHC942_n3311 (.O(FE_PHN942_n3311), 
	.I(n3311));
   DELDKHD FE_PHC941_n779 (.O(FE_PHN941_n779), 
	.I(n779));
   DELDKHD FE_PHC940_n2848 (.O(FE_PHN940_n2848), 
	.I(n2848));
   DELDKHD FE_PHC939_n3202 (.O(FE_PHN939_n3202), 
	.I(n3202));
   DELDKHD FE_PHC938_n1446 (.O(FE_PHN938_n1446), 
	.I(n1446));
   DELDKHD FE_PHC937_n1152 (.O(FE_PHN937_n1152), 
	.I(n1152));
   DELDKHD FE_PHC936_n3648 (.O(FE_PHN936_n3648), 
	.I(n3648));
   DELDKHD FE_PHC935_n2128 (.O(FE_PHN935_n2128), 
	.I(n2128));
   DELDKHD FE_PHC934_n813 (.O(FE_PHN934_n813), 
	.I(n813));
   DELDKHD FE_PHC933_n942 (.O(FE_PHN933_n942), 
	.I(n942));
   DELDKHD FE_PHC932_n1165 (.O(FE_PHN932_n1165), 
	.I(n1165));
   DELDKHD FE_PHC931_n1439 (.O(FE_PHN931_n1439), 
	.I(n1439));
   DELDKHD FE_PHC930_n2518 (.O(FE_PHN930_n2518), 
	.I(n2518));
   DELDKHD FE_PHC929_n1627 (.O(FE_PHN929_n1627), 
	.I(n1627));
   DELDKHD FE_PHC928_n2094 (.O(FE_PHN928_n2094), 
	.I(n2094));
   DELDKHD FE_PHC927_n1380 (.O(FE_PHN927_n1380), 
	.I(n1380));
   DELDKHD FE_PHC926_n1845 (.O(FE_PHN926_n1845), 
	.I(n1845));
   DELDKHD FE_PHC925_n3159 (.O(FE_PHN925_n3159), 
	.I(n3159));
   DELDKHD FE_PHC924_n4156 (.O(FE_PHN924_n4156), 
	.I(n4156));
   DELDKHD FE_PHC923_n1523 (.O(FE_PHN923_n1523), 
	.I(n1523));
   DELDKHD FE_PHC922_n606 (.O(FE_PHN922_n606), 
	.I(n606));
   DELDKHD FE_PHC921_n4528 (.O(FE_PHN921_n4528), 
	.I(n4528));
   DELDKHD FE_PHC920_n2638 (.O(FE_PHN920_n2638), 
	.I(n2638));
   DELDKHD FE_PHC919_n3530 (.O(FE_PHN919_n3530), 
	.I(n3530));
   DELDKHD FE_PHC918_n1433 (.O(FE_PHN918_n1433), 
	.I(n1433));
   DELDKHD FE_PHC917_n3576 (.O(FE_PHN917_n3576), 
	.I(n3576));
   DELDKHD FE_PHC916_n1890 (.O(FE_PHN916_n1890), 
	.I(n1890));
   DELDKHD FE_PHC915_n1745 (.O(FE_PHN915_n1745), 
	.I(n1745));
   DELDKHD FE_PHC914_n1570 (.O(FE_PHN914_n1570), 
	.I(n1570));
   DELDKHD FE_PHC913_n3767 (.O(FE_PHN913_n3767), 
	.I(n3767));
   DELDKHD FE_PHC912_n3628 (.O(FE_PHN912_n3628), 
	.I(n3628));
   DELDKHD FE_PHC911_n1667 (.O(FE_PHN911_n1667), 
	.I(n1667));
   DELDKHD FE_PHC910_n2334 (.O(FE_PHN910_n2334), 
	.I(n2334));
   DELDKHD FE_PHC909_n3737 (.O(FE_PHN909_n3737), 
	.I(n3737));
   DELDKHD FE_PHC908_n1184 (.O(FE_PHN908_n1184), 
	.I(n1184));
   DELDKHD FE_PHC907_n1675 (.O(FE_PHN907_n1675), 
	.I(n1675));
   DELDKHD FE_PHC906_n3804 (.O(FE_PHN906_n3804), 
	.I(n3804));
   DELDKHD FE_PHC905_n1841 (.O(FE_PHN905_n1841), 
	.I(n1841));
   DELDKHD FE_PHC904_n3685 (.O(FE_PHN904_n3685), 
	.I(n3685));
   DELDKHD FE_PHC903_n3829 (.O(FE_PHN903_n3829), 
	.I(n3829));
   DELDKHD FE_PHC902_n4595 (.O(FE_PHN902_n4595), 
	.I(n4595));
   DELDKHD FE_PHC901_n2808 (.O(FE_PHN901_n2808), 
	.I(n2808));
   DELDKHD FE_PHC900_n4625 (.O(FE_PHN900_n4625), 
	.I(n4625));
   DELDKHD FE_PHC899_n1100 (.O(FE_PHN899_n1100), 
	.I(n1100));
   DELDKHD FE_PHC898_n3907 (.O(FE_PHN898_n3907), 
	.I(n3907));
   DELDKHD FE_PHC897_n2312 (.O(FE_PHN897_n2312), 
	.I(n2312));
   DELDKHD FE_PHC896_n2197 (.O(FE_PHN896_n2197), 
	.I(n2197));
   DELDKHD FE_PHC895_n1715 (.O(FE_PHN895_n1715), 
	.I(n1715));
   DELDKHD FE_PHC894_n3360 (.O(FE_PHN894_n3360), 
	.I(n3360));
   DELDKHD FE_PHC893_n800 (.O(FE_PHN893_n800), 
	.I(n800));
   DELDKHD FE_PHC892_n2849 (.O(FE_PHN892_n2849), 
	.I(n2849));
   DELDKHD FE_PHC891_n3761 (.O(FE_PHN891_n3761), 
	.I(n3761));
   DELDKHD FE_PHC890_n4422 (.O(FE_PHN890_n4422), 
	.I(n4422));
   DELDKHD FE_PHC889_n4498 (.O(FE_PHN889_n4498), 
	.I(n4498));
   DELDKHD FE_PHC888_n932 (.O(FE_PHN888_n932), 
	.I(n932));
   DELDKHD FE_PHC887_n2221 (.O(FE_PHN887_n2221), 
	.I(n2221));
   DELDKHD FE_PHC886_n2439 (.O(FE_PHN886_n2439), 
	.I(n2439));
   DELDKHD FE_PHC885_n1811 (.O(FE_PHN885_n1811), 
	.I(n1811));
   DELDKHD FE_PHC884_n4516 (.O(FE_PHN884_n4516), 
	.I(n4516));
   DELDKHD FE_PHC883_n2352 (.O(FE_PHN883_n2352), 
	.I(n2352));
   DELDKHD FE_PHC882_n3248 (.O(FE_PHN882_n3248), 
	.I(n3248));
   DELDKHD FE_PHC881_n2484 (.O(FE_PHN881_n2484), 
	.I(n2484));
   DELDKHD FE_PHC880_n2751 (.O(FE_PHN880_n2751), 
	.I(n2751));
   DELDKHD FE_PHC879_n3832 (.O(FE_PHN879_n3832), 
	.I(n3832));
   DELDKHD FE_PHC878_n4572 (.O(FE_PHN878_n4572), 
	.I(n4572));
   DELDKHD FE_PHC877_n818 (.O(FE_PHN877_n818), 
	.I(n818));
   DELDKHD FE_PHC876_n612 (.O(FE_PHN876_n612), 
	.I(n612));
   DELDKHD FE_PHC875_n1188 (.O(FE_PHN875_n1188), 
	.I(n1188));
   DELDKHD FE_PHC874_n775 (.O(FE_PHN874_n775), 
	.I(n775));
   DELDKHD FE_PHC873_n1801 (.O(FE_PHN873_n1801), 
	.I(n1801));
   DELDKHD FE_PHC872_n2809 (.O(FE_PHN872_n2809), 
	.I(n2809));
   DELCKHD FE_PHC871_ram_249__12_ (.O(FE_PHN871_ram_249__12_), 
	.I(\ram[249][12] ));
   DELCKHD FE_PHC870_n1128 (.O(FE_PHN870_n1128), 
	.I(n1128));
   DELCKHD FE_PHC869_n3745 (.O(FE_PHN869_n3745), 
	.I(n3745));
   DELCKHD FE_PHC868_n4253 (.O(FE_PHN868_n4253), 
	.I(n4253));
   DELCKHD FE_PHC867_n2776 (.O(FE_PHN867_n2776), 
	.I(n2776));
   DELCKHD FE_PHC866_n3828 (.O(FE_PHN866_n3828), 
	.I(n3828));
   DELCKHD FE_PHC865_n1777 (.O(FE_PHN865_n1777), 
	.I(n1777));
   DELCKHD FE_PHC864_n3404 (.O(FE_PHN864_n3404), 
	.I(n3404));
   DELCKHD FE_PHC863_n4136 (.O(FE_PHN863_n4136), 
	.I(n4136));
   DELCKHD FE_PHC862_n3879 (.O(FE_PHN862_n3879), 
	.I(n3879));
   DELCKHD FE_PHC861_n4545 (.O(FE_PHN861_n4545), 
	.I(n4545));
   DELCKHD FE_PHC860_n3486 (.O(FE_PHN860_n3486), 
	.I(n3486));
   DELCKHD FE_PHC859_n3176 (.O(FE_PHN859_n3176), 
	.I(n3176));
   DELCKHD FE_PHC858_n4293 (.O(FE_PHN858_n4293), 
	.I(n4293));
   DELCKHD FE_PHC857_n1191 (.O(FE_PHN857_n1191), 
	.I(n1191));
   DELCKHD FE_PHC856_n2253 (.O(FE_PHN856_n2253), 
	.I(n2253));
   DELCKHD FE_PHC855_n4337 (.O(FE_PHN855_n4337), 
	.I(n4337));
   DELCKHD FE_PHC854_n741 (.O(FE_PHN854_n741), 
	.I(n741));
   DELCKHD FE_PHC853_n3720 (.O(FE_PHN853_n3720), 
	.I(n3720));
   DELCKHD FE_PHC852_n3760 (.O(FE_PHN852_n3760), 
	.I(n3760));
   DELCKHD FE_PHC851_n3307 (.O(FE_PHN851_n3307), 
	.I(n3307));
   DELCKHD FE_PHC850_n4085 (.O(FE_PHN850_n4085), 
	.I(n4085));
   DELCKHD FE_PHC849_n4523 (.O(FE_PHN849_n4523), 
	.I(n4523));
   DELCKHD FE_PHC848_n723 (.O(FE_PHN848_n723), 
	.I(n723));
   DELCKHD FE_PHC847_n4058 (.O(FE_PHN847_n4058), 
	.I(n4058));
   DELCKHD FE_PHC846_n4198 (.O(FE_PHN846_n4198), 
	.I(n4198));
   DELCKHD FE_PHC845_n1800 (.O(FE_PHN845_n1800), 
	.I(n1800));
   DELCKHD FE_PHC844_n3288 (.O(FE_PHN844_n3288), 
	.I(n3288));
   DELCKHD FE_PHC843_n4099 (.O(FE_PHN843_n4099), 
	.I(n4099));
   DELCKHD FE_PHC842_n3296 (.O(FE_PHN842_n3296), 
	.I(n3296));
   DELCKHD FE_PHC841_n3551 (.O(FE_PHN841_n3551), 
	.I(n3551));
   DELCKHD FE_PHC840_n2899 (.O(FE_PHN840_n2899), 
	.I(n2899));
   DELCKHD FE_PHC839_n875 (.O(FE_PHN839_n875), 
	.I(n875));
   DELCKHD FE_PHC838_n3675 (.O(FE_PHN838_n3675), 
	.I(n3675));
   DELCKHD FE_PHC837_n1089 (.O(FE_PHN837_n1089), 
	.I(n1089));
   DELCKHD FE_PHC836_n3271 (.O(FE_PHN836_n3271), 
	.I(n3271));
   DELCKHD FE_PHC835_n1170 (.O(FE_PHN835_n1170), 
	.I(n1170));
   DELCKHD FE_PHC834_n1827 (.O(FE_PHN834_n1827), 
	.I(n1827));
   DELCKHD FE_PHC833_n2939 (.O(FE_PHN833_n2939), 
	.I(n2939));
   DELCKHD FE_PHC832_n1004 (.O(FE_PHN832_n1004), 
	.I(n1004));
   DELCKHD FE_PHC831_n1479 (.O(FE_PHN831_n1479), 
	.I(n1479));
   DELCKHD FE_PHC830_n2129 (.O(FE_PHN830_n2129), 
	.I(n2129));
   DELCKHD FE_PHC829_n3201 (.O(FE_PHN829_n3201), 
	.I(n3201));
   DELCKHD FE_PHC828_n3222 (.O(FE_PHN828_n3222), 
	.I(n3222));
   DELCKHD FE_PHC827_n3643 (.O(FE_PHN827_n3643), 
	.I(n3643));
   DELCKHD FE_PHC826_n2418 (.O(FE_PHN826_n2418), 
	.I(n2418));
   DELCKHD FE_PHC825_n3418 (.O(FE_PHN825_n3418), 
	.I(n3418));
   DELCKHD FE_PHC824_n3925 (.O(FE_PHN824_n3925), 
	.I(n3925));
   DELCKHD FE_PHC823_n1526 (.O(FE_PHN823_n1526), 
	.I(n1526));
   DELCKHD FE_PHC822_n1187 (.O(FE_PHN822_n1187), 
	.I(n1187));
   DELCKHD FE_PHC821_n3528 (.O(FE_PHN821_n3528), 
	.I(n3528));
   DELCKHD FE_PHC820_n2307 (.O(FE_PHN820_n2307), 
	.I(n2307));
   DELCKHD FE_PHC819_n4473 (.O(FE_PHN819_n4473), 
	.I(n4473));
   DELCKHD FE_PHC818_n2835 (.O(FE_PHN818_n2835), 
	.I(n2835));
   DELCKHD FE_PHC817_n1502 (.O(FE_PHN817_n1502), 
	.I(n1502));
   DELCKHD FE_PHC816_n859 (.O(FE_PHN816_n859), 
	.I(n859));
   DELCKHD FE_PHC815_n3423 (.O(FE_PHN815_n3423), 
	.I(n3423));
   DELCKHD FE_PHC814_n3485 (.O(FE_PHN814_n3485), 
	.I(n3485));
   DELCKHD FE_PHC813_n2717 (.O(FE_PHN813_n2717), 
	.I(n2717));
   DELCKHD FE_PHC812_n2797 (.O(FE_PHN812_n2797), 
	.I(n2797));
   DELCKHD FE_PHC811_n3724 (.O(FE_PHN811_n3724), 
	.I(n3724));
   DELCKHD FE_PHC810_n3871 (.O(FE_PHN810_n3871), 
	.I(n3871));
   DELCKHD FE_PHC809_n1440 (.O(FE_PHN809_n1440), 
	.I(n1440));
   DELCKHD FE_PHC808_n1524 (.O(FE_PHN808_n1524), 
	.I(n1524));
   DELCKHD FE_PHC807_n1882 (.O(FE_PHN807_n1882), 
	.I(n1882));
   DELCKHD FE_PHC806_n2947 (.O(FE_PHN806_n2947), 
	.I(n2947));
   DELCKHD FE_PHC805_n3168 (.O(FE_PHN805_n3168), 
	.I(n3168));
   DELCKHD FE_PHC804_n751 (.O(FE_PHN804_n751), 
	.I(n751));
   DELCKHD FE_PHC803_n1255 (.O(FE_PHN803_n1255), 
	.I(n1255));
   DELCKHD FE_PHC802_n1650 (.O(FE_PHN802_n1650), 
	.I(n1650));
   DELCKHD FE_PHC801_n4651 (.O(FE_PHN801_n4651), 
	.I(n4651));
   DELCKHD FE_PHC800_n1561 (.O(FE_PHN800_n1561), 
	.I(n1561));
   DELCKHD FE_PHC799_n1683 (.O(FE_PHN799_n1683), 
	.I(n1683));
   DELCKHD FE_PHC798_n2488 (.O(FE_PHN798_n2488), 
	.I(n2488));
   DELCKHD FE_PHC797_n1612 (.O(FE_PHN797_n1612), 
	.I(n1612));
   DELCKHD FE_PHC796_n2107 (.O(FE_PHN796_n2107), 
	.I(n2107));
   DELCKHD FE_PHC795_n2781 (.O(FE_PHN795_n2781), 
	.I(n2781));
   DELCKHD FE_PHC794_n4521 (.O(FE_PHN794_n4521), 
	.I(n4521));
   DELCKHD FE_PHC793_n2404 (.O(FE_PHN793_n2404), 
	.I(n2404));
   DELCKHD FE_PHC792_n1751 (.O(FE_PHN792_n1751), 
	.I(n1751));
   DELCKHD FE_PHC791_n2799 (.O(FE_PHN791_n2799), 
	.I(n2799));
   DELCKHD FE_PHC790_n3244 (.O(FE_PHN790_n3244), 
	.I(n3244));
   DELCKHD FE_PHC789_n4424 (.O(FE_PHN789_n4424), 
	.I(n4424));
   DELCKHD FE_PHC788_n2678 (.O(FE_PHN788_n2678), 
	.I(n2678));
   DELCKHD FE_PHC787_n1629 (.O(FE_PHN787_n1629), 
	.I(n1629));
   DELCKHD FE_PHC786_n2150 (.O(FE_PHN786_n2150), 
	.I(n2150));
   DELCKHD FE_PHC785_n3306 (.O(FE_PHN785_n3306), 
	.I(n3306));
   DELCKHD FE_PHC784_n4555 (.O(FE_PHN784_n4555), 
	.I(n4555));
   DELCKHD FE_PHC783_n4638 (.O(FE_PHN783_n4638), 
	.I(n4638));
   DELCKHD FE_PHC782_n3421 (.O(FE_PHN782_n3421), 
	.I(n3421));
   DELCKHD FE_PHC781_n4663 (.O(FE_PHN781_n4663), 
	.I(n4663));
   DELCKHD FE_PHC780_n2260 (.O(FE_PHN780_n2260), 
	.I(n2260));
   DELCKHD FE_PHC779_n3710 (.O(FE_PHN779_n3710), 
	.I(n3710));
   DELCKHD FE_PHC778_n3796 (.O(FE_PHN778_n3796), 
	.I(n3796));
   DELCKHD FE_PHC777_n4066 (.O(FE_PHN777_n4066), 
	.I(n4066));
   DELCKHD FE_PHC776_n2459 (.O(FE_PHN776_n2459), 
	.I(n2459));
   DELCKHD FE_PHC775_n619 (.O(FE_PHN775_n619), 
	.I(n619));
   DELCKHD FE_PHC774_n1597 (.O(FE_PHN774_n1597), 
	.I(n1597));
   DELCKHD FE_PHC773_n3238 (.O(FE_PHN773_n3238), 
	.I(n3238));
   DELCKHD FE_PHC772_n3708 (.O(FE_PHN772_n3708), 
	.I(n3708));
   DELCKHD FE_PHC771_n4554 (.O(FE_PHN771_n4554), 
	.I(n4554));
   DELCKHD FE_PHC770_n3366 (.O(FE_PHN770_n3366), 
	.I(n3366));
   DELCKHD FE_PHC769_n3699 (.O(FE_PHN769_n3699), 
	.I(n3699));
   DELCKHD FE_PHC768_n2597 (.O(FE_PHN768_n2597), 
	.I(n2597));
   DELCKHD FE_PHC767_n3587 (.O(FE_PHN767_n3587), 
	.I(n3587));
   DELCKHD FE_PHC766_n4425 (.O(FE_PHN766_n4425), 
	.I(n4425));
   DELCKHD FE_PHC765_n4072 (.O(FE_PHN765_n4072), 
	.I(n4072));
   DELCKHD FE_PHC764_n860 (.O(FE_PHN764_n860), 
	.I(n860));
   DELCKHD FE_PHC763_n3324 (.O(FE_PHN763_n3324), 
	.I(n3324));
   DELCKHD FE_PHC762_n3465 (.O(FE_PHN762_n3465), 
	.I(n3465));
   DELCKHD FE_PHC761_n4287 (.O(FE_PHN761_n4287), 
	.I(n4287));
   DELCKHD FE_PHC760_n1720 (.O(FE_PHN760_n1720), 
	.I(n1720));
   DELCKHD FE_PHC759_n3479 (.O(FE_PHN759_n3479), 
	.I(n3479));
   DELCKHD FE_PHC758_n4083 (.O(FE_PHN758_n4083), 
	.I(n4083));
   DELCKHD FE_PHC757_n603 (.O(FE_PHN757_n603), 
	.I(n603));
   DELCKHD FE_PHC756_n2436 (.O(FE_PHN756_n2436), 
	.I(n2436));
   DELCKHD FE_PHC755_n3349 (.O(FE_PHN755_n3349), 
	.I(n3349));
   DELCKHD FE_PHC754_n3645 (.O(FE_PHN754_n3645), 
	.I(n3645));
   DELCKHD FE_PHC753_n640 (.O(FE_PHN753_n640), 
	.I(n640));
   DELCKHD FE_PHC752_n1057 (.O(FE_PHN752_n1057), 
	.I(n1057));
   DELCKHD FE_PHC751_n1475 (.O(FE_PHN751_n1475), 
	.I(n1475));
   DELCKHD FE_PHC750_n1105 (.O(FE_PHN750_n1105), 
	.I(n1105));
   DELCKHD FE_PHC749_n1145 (.O(FE_PHN749_n1145), 
	.I(n1145));
   DELCKHD FE_PHC748_n1657 (.O(FE_PHN748_n1657), 
	.I(n1657));
   DELCKHD FE_PHC747_n2783 (.O(FE_PHN747_n2783), 
	.I(n2783));
   DELCKHD FE_PHC746_n2143 (.O(FE_PHN746_n2143), 
	.I(n2143));
   DELCKHD FE_PHC745_n750 (.O(FE_PHN745_n750), 
	.I(n750));
   DELCKHD FE_PHC744_n1680 (.O(FE_PHN744_n1680), 
	.I(n1680));
   DELCKHD FE_PHC743_n2222 (.O(FE_PHN743_n2222), 
	.I(n2222));
   DELCKHD FE_PHC742_n4113 (.O(FE_PHN742_n4113), 
	.I(n4113));
   DELCKHD FE_PHC741_n3885 (.O(FE_PHN741_n3885), 
	.I(n3885));
   DELCKHD FE_PHC740_n4302 (.O(FE_PHN740_n4302), 
	.I(n4302));
   DELCKHD FE_PHC739_n1885 (.O(FE_PHN739_n1885), 
	.I(n1885));
   DELCKHD FE_PHC738_n3277 (.O(FE_PHN738_n3277), 
	.I(n3277));
   DELCKHD FE_PHC737_n3853 (.O(FE_PHN737_n3853), 
	.I(n3853));
   DELCKHD FE_PHC736_n2085 (.O(FE_PHN736_n2085), 
	.I(n2085));
   DELCKHD FE_PHC735_n2219 (.O(FE_PHN735_n2219), 
	.I(n2219));
   DELCKHD FE_PHC734_n1604 (.O(FE_PHN734_n1604), 
	.I(n1604));
   DELCKHD FE_PHC733_n2084 (.O(FE_PHN733_n2084), 
	.I(n2084));
   DELCKHD FE_PHC732_n3194 (.O(FE_PHN732_n3194), 
	.I(n3194));
   DELCKHD FE_PHC731_n2441 (.O(FE_PHN731_n2441), 
	.I(n2441));
   DELCKHD FE_PHC730_n3356 (.O(FE_PHN730_n3356), 
	.I(n3356));
   DELCKHD FE_PHC729_n728 (.O(FE_PHN729_n728), 
	.I(n728));
   DELCKHD FE_PHC728_n1716 (.O(FE_PHN728_n1716), 
	.I(n1716));
   DELCKHD FE_PHC727_n2211 (.O(FE_PHN727_n2211), 
	.I(n2211));
   DELCKHD FE_PHC726_n3171 (.O(FE_PHN726_n3171), 
	.I(n3171));
   DELCKHD FE_PHC725_n4349 (.O(FE_PHN725_n4349), 
	.I(n4349));
   DELCKHD FE_PHC724_n4518 (.O(FE_PHN724_n4518), 
	.I(n4518));
   DELCKHD FE_PHC723_n3573 (.O(FE_PHN723_n3573), 
	.I(n3573));
   DELCKHD FE_PHC722_n4659 (.O(FE_PHN722_n4659), 
	.I(n4659));
   DELCKHD FE_PHC721_n4501 (.O(FE_PHN721_n4501), 
	.I(n4501));
   DELCKHD FE_PHC720_n4519 (.O(FE_PHN720_n4519), 
	.I(n4519));
   DELCKHD FE_PHC719_n1703 (.O(FE_PHN719_n1703), 
	.I(n1703));
   DELCKHD FE_PHC718_n733 (.O(FE_PHN718_n733), 
	.I(n733));
   DELCKHD FE_PHC717_n1052 (.O(FE_PHN717_n1052), 
	.I(n1052));
   DELCKHD FE_PHC716_n1608 (.O(FE_PHN716_n1608), 
	.I(n1608));
   DELCKHD FE_PHC715_n2173 (.O(FE_PHN715_n2173), 
	.I(n2173));
   DELCKHD FE_PHC714_n4091 (.O(FE_PHN714_n4091), 
	.I(n4091));
   DELCKHD FE_PHC713_n1144 (.O(FE_PHN713_n1144), 
	.I(n1144));
   DELCKHD FE_PHC712_n1298 (.O(FE_PHN712_n1298), 
	.I(n1298));
   DELCKHD FE_PHC711_n3511 (.O(FE_PHN711_n3511), 
	.I(n3511));
   DELDKHD FE_PHC710_n1820 (.O(FE_PHN710_n1820), 
	.I(n1820));
   DELDKHD FE_PHC709_n3733 (.O(FE_PHN709_n3733), 
	.I(n3733));
   DELDKHD FE_PHC708_n3941 (.O(FE_PHN708_n3941), 
	.I(n3941));
   DELDKHD FE_PHC707_n3651 (.O(FE_PHN707_n3651), 
	.I(n3651));
   DELDKHD FE_PHC706_n3061 (.O(FE_PHN706_n3061), 
	.I(n3061));
   DELDKHD FE_PHC705_n3267 (.O(FE_PHN705_n3267), 
	.I(n3267));
   DELDKHD FE_PHC704_n3575 (.O(FE_PHN704_n3575), 
	.I(n3575));
   DELDKHD FE_PHC703_n2739 (.O(FE_PHN703_n2739), 
	.I(n2739));
   DELDKHD FE_PHC702_n2271 (.O(FE_PHN702_n2271), 
	.I(n2271));
   DELDKHD FE_PHC701_n3875 (.O(FE_PHN701_n3875), 
	.I(n3875));
   DELDKHD FE_PHC700_n4495 (.O(FE_PHN700_n4495), 
	.I(n4495));
   DELDKHD FE_PHC699_n3759 (.O(FE_PHN699_n3759), 
	.I(n3759));
   DELDKHD FE_PHC698_n2911 (.O(FE_PHN698_n2911), 
	.I(n2911));
   DELDKHD FE_PHC697_n2905 (.O(FE_PHN697_n2905), 
	.I(n2905));
   DELDKHD FE_PHC696_n820 (.O(FE_PHN696_n820), 
	.I(n820));
   DELDKHD FE_PHC695_n4056 (.O(FE_PHN695_n4056), 
	.I(n4056));
   DELDKHD FE_PHC694_n4668 (.O(FE_PHN694_n4668), 
	.I(n4668));
   DELDKHD FE_PHC693_n1480 (.O(FE_PHN693_n1480), 
	.I(n1480));
   DELDKHD FE_PHC692_n3498 (.O(FE_PHN692_n3498), 
	.I(n3498));
   DELDKHD FE_PHC691_n1831 (.O(FE_PHN691_n1831), 
	.I(n1831));
   DELDKHD FE_PHC690_n2269 (.O(FE_PHN690_n2269), 
	.I(n2269));
   DELDKHD FE_PHC689_n2276 (.O(FE_PHN689_n2276), 
	.I(n2276));
   DELDKHD FE_PHC688_n2811 (.O(FE_PHN688_n2811), 
	.I(n2811));
   DELDKHD FE_PHC687_n1887 (.O(FE_PHN687_n1887), 
	.I(n1887));
   DELDKHD FE_PHC686_n1889 (.O(FE_PHN686_n1889), 
	.I(n1889));
   DELDKHD FE_PHC685_n4436 (.O(FE_PHN685_n4436), 
	.I(n4436));
   DELDKHD FE_PHC684_n4532 (.O(FE_PHN684_n4532), 
	.I(n4532));
   DELDKHD FE_PHC683_n1647 (.O(FE_PHN683_n1647), 
	.I(n1647));
   DELDKHD FE_PHC682_n4643 (.O(FE_PHN682_n4643), 
	.I(n4643));
   DELDKHD FE_PHC681_n1771 (.O(FE_PHN681_n1771), 
	.I(n1771));
   DELDKHD FE_PHC680_n4669 (.O(FE_PHN680_n4669), 
	.I(n4669));
   DELDKHD FE_PHC679_n4434 (.O(FE_PHN679_n4434), 
	.I(n4434));
   DELDKHD FE_PHC678_n1175 (.O(FE_PHN678_n1175), 
	.I(n1175));
   DELDKHD FE_PHC677_n1496 (.O(FE_PHN677_n1496), 
	.I(n1496));
   DELDKHD FE_PHC676_n2673 (.O(FE_PHN676_n2673), 
	.I(n2673));
   DELDKHD FE_PHC675_n3113 (.O(FE_PHN675_n3113), 
	.I(n3113));
   DELDKHD FE_PHC674_n1494 (.O(FE_PHN674_n1494), 
	.I(n1494));
   DELDKHD FE_PHC673_n2914 (.O(FE_PHN673_n2914), 
	.I(n2914));
   DELDKHD FE_PHC672_n2527 (.O(FE_PHN672_n2527), 
	.I(n2527));
   DELDKHD FE_PHC671_n2507 (.O(FE_PHN671_n2507), 
	.I(n2507));
   DELDKHD FE_PHC670_n4459 (.O(FE_PHN670_n4459), 
	.I(n4459));
   DELDKHD FE_PHC669_n4665 (.O(FE_PHN669_n4665), 
	.I(n4665));
   DELDKHD FE_PHC668_n1247 (.O(FE_PHN668_n1247), 
	.I(n1247));
   DELDKHD FE_PHC667_n1367 (.O(FE_PHN667_n1367), 
	.I(n1367));
   DELDKHD FE_PHC666_n3702 (.O(FE_PHN666_n3702), 
	.I(n3702));
   DELDKHD FE_PHC665_n4576 (.O(FE_PHN665_n4576), 
	.I(n4576));
   DELDKHD FE_PHC664_n2139 (.O(FE_PHN664_n2139), 
	.I(n2139));
   DELDKHD FE_PHC663_ram_109__5_ (.O(FE_PHN663_ram_109__5_), 
	.I(\ram[109][5] ));
   DELDKHD FE_PHC662_n4517 (.O(FE_PHN662_n4517), 
	.I(n4517));
   DELDKHD FE_PHC661_n2270 (.O(FE_PHN661_n2270), 
	.I(n2270));
   DELDKHD FE_PHC660_n1445 (.O(FE_PHN660_n1445), 
	.I(n1445));
   DELDKHD FE_PHC659_n1740 (.O(FE_PHN659_n1740), 
	.I(n1740));
   DELDKHD FE_PHC658_n3882 (.O(FE_PHN658_n3882), 
	.I(n3882));
   DELDKHD FE_PHC657_n3297 (.O(FE_PHN657_n3297), 
	.I(n3297));
   DELDKHD FE_PHC656_n2519 (.O(FE_PHN656_n2519), 
	.I(n2519));
   DELDKHD FE_PHC655_n4639 (.O(FE_PHN655_n4639), 
	.I(n4639));
   DELDKHD FE_PHC654_n1249 (.O(FE_PHN654_n1249), 
	.I(n1249));
   DELDKHD FE_PHC653_n1640 (.O(FE_PHN653_n1640), 
	.I(n1640));
   DELDKHD FE_PHC652_n1697 (.O(FE_PHN652_n1697), 
	.I(n1697));
   DELDKHD FE_PHC651_n2655 (.O(FE_PHN651_n2655), 
	.I(n2655));
   DELDKHD FE_PHC650_n2463 (.O(FE_PHN650_n2463), 
	.I(n2463));
   DELDKHD FE_PHC649_n3059 (.O(FE_PHN649_n3059), 
	.I(n3059));
   DELDKHD FE_PHC648_n1035 (.O(FE_PHN648_n1035), 
	.I(n1035));
   DELDKHD FE_PHC647_n1828 (.O(FE_PHN647_n1828), 
	.I(n1828));
   DELDKHD FE_PHC646_n2532 (.O(FE_PHN646_n2532), 
	.I(n2532));
   DELDKHD FE_PHC645_n3312 (.O(FE_PHN645_n3312), 
	.I(n3312));
   DELDKHD FE_PHC644_n3313 (.O(FE_PHN644_n3313), 
	.I(n3313));
   DELDKHD FE_PHC643_n3501 (.O(FE_PHN643_n3501), 
	.I(n3501));
   DELDKHD FE_PHC642_n2852 (.O(FE_PHN642_n2852), 
	.I(n2852));
   DELDKHD FE_PHC641_n1559 (.O(FE_PHN641_n1559), 
	.I(n1559));
   DELDKHD FE_PHC640_n3245 (.O(FE_PHN640_n3245), 
	.I(n3245));
   DELDKHD FE_PHC639_n4443 (.O(FE_PHN639_n4443), 
	.I(n4443));
   DELDKHD FE_PHC638_n3591 (.O(FE_PHN638_n3591), 
	.I(n3591));
   DELDKHD FE_PHC637_n1176 (.O(FE_PHN637_n1176), 
	.I(n1176));
   DELDKHD FE_PHC636_n3513 (.O(FE_PHN636_n3513), 
	.I(n3513));
   DELDKHD FE_PHC635_n1116 (.O(FE_PHN635_n1116), 
	.I(n1116));
   DELDKHD FE_PHC634_n2710 (.O(FE_PHN634_n2710), 
	.I(n2710));
   DELDKHD FE_PHC633_n4618 (.O(FE_PHN633_n4618), 
	.I(n4618));
   DELDKHD FE_PHC632_n666 (.O(FE_PHN632_n666), 
	.I(n666));
   DELDKHD FE_PHC631_n1493 (.O(FE_PHN631_n1493), 
	.I(n1493));
   DELDKHD FE_PHC630_n1798 (.O(FE_PHN630_n1798), 
	.I(n1798));
   DELDKHD FE_PHC629_n2444 (.O(FE_PHN629_n2444), 
	.I(n2444));
   DELDKHD FE_PHC628_n2508 (.O(FE_PHN628_n2508), 
	.I(n2508));
   DELDKHD FE_PHC627_n2895 (.O(FE_PHN627_n2895), 
	.I(n2895));
   DELDKHD FE_PHC626_n4590 (.O(FE_PHN626_n4590), 
	.I(n4590));
   DELDKHD FE_PHC625_n4599 (.O(FE_PHN625_n4599), 
	.I(n4599));
   DELDKHD FE_PHC624_n4280 (.O(FE_PHN624_n4280), 
	.I(n4280));
   DELDKHD FE_PHC623_n806 (.O(FE_PHN623_n806), 
	.I(n806));
   DELDKHD FE_PHC622_n2238 (.O(FE_PHN622_n2238), 
	.I(n2238));
   DELDKHD FE_PHC621_n3973 (.O(FE_PHN621_n3973), 
	.I(n3973));
   DELDKHD FE_PHC620_n2288 (.O(FE_PHN620_n2288), 
	.I(n2288));
   DELDKHD FE_PHC619_n2632 (.O(FE_PHN619_n2632), 
	.I(n2632));
   DELDKHD FE_PHC618_n4095 (.O(FE_PHN618_n4095), 
	.I(n4095));
   DELDKHD FE_PHC617_n1861 (.O(FE_PHN617_n1861), 
	.I(n1861));
   DELDKHD FE_PHC616_n4161 (.O(FE_PHN616_n4161), 
	.I(n4161));
   DELDKHD FE_PHC615_n3344 (.O(FE_PHN615_n3344), 
	.I(n3344));
   DELDKHD FE_PHC614_n1160 (.O(FE_PHN614_n1160), 
	.I(n1160));
   DELDKHD FE_PHC613_n2850 (.O(FE_PHN613_n2850), 
	.I(n2850));
   DELDKHD FE_PHC612_n2586 (.O(FE_PHN612_n2586), 
	.I(n2586));
   DELDKHD FE_PHC611_n1547 (.O(FE_PHN611_n1547), 
	.I(n1547));
   DELDKHD FE_PHC610_n3909 (.O(FE_PHN610_n3909), 
	.I(n3909));
   DELDKHD FE_PHC609_n4451 (.O(FE_PHN609_n4451), 
	.I(n4451));
   DELDKHD FE_PHC608_n2089 (.O(FE_PHN608_n2089), 
	.I(n2089));
   DELDKHD FE_PHC607_n3680 (.O(FE_PHN607_n3680), 
	.I(n3680));
   DELDKHD FE_PHC606_n1760 (.O(FE_PHN606_n1760), 
	.I(n1760));
   DELDKHD FE_PHC605_n1722 (.O(FE_PHN605_n1722), 
	.I(n1722));
   DELDKHD FE_PHC604_n4080 (.O(FE_PHN604_n4080), 
	.I(n4080));
   DELDKHD FE_PHC603_n1431 (.O(FE_PHN603_n1431), 
	.I(n1431));
   DELDKHD FE_PHC602_n1821 (.O(FE_PHN602_n1821), 
	.I(n1821));
   DELDKHD FE_PHC601_n602 (.O(FE_PHN601_n602), 
	.I(n602));
   DELDKHD FE_PHC600_n2265 (.O(FE_PHN600_n2265), 
	.I(n2265));
   DELDKHD FE_PHC599_n2585 (.O(FE_PHN599_n2585), 
	.I(n2585));
   DELDKHD FE_PHC598_n4466 (.O(FE_PHN598_n4466), 
	.I(n4466));
   DELDKHD FE_PHC597_n3468 (.O(FE_PHN597_n3468), 
	.I(n3468));
   DELDKHD FE_PHC596_n3663 (.O(FE_PHN596_n3663), 
	.I(n3663));
   DELDKHD FE_PHC595_n3438 (.O(FE_PHN595_n3438), 
	.I(n3438));
   DELDKHD FE_PHC594_n1834 (.O(FE_PHN594_n1834), 
	.I(n1834));
   DELDKHD FE_PHC593_n2284 (.O(FE_PHN593_n2284), 
	.I(n2284));
   DELDKHD FE_PHC592_n2553 (.O(FE_PHN592_n2553), 
	.I(n2553));
   DELDKHD FE_PHC591_n1702 (.O(FE_PHN591_n1702), 
	.I(n1702));
   DELDKHD FE_PHC590_n2229 (.O(FE_PHN590_n2229), 
	.I(n2229));
   DELDKHD FE_PHC589_n2721 (.O(FE_PHN589_n2721), 
	.I(n2721));
   DELDKHD FE_PHC588_n2859 (.O(FE_PHN588_n2859), 
	.I(n2859));
   DELDKHD FE_PHC587_n4623 (.O(FE_PHN587_n4623), 
	.I(n4623));
   DELDKHD FE_PHC586_n3509 (.O(FE_PHN586_n3509), 
	.I(n3509));
   DELDKHD FE_PHC585_n931 (.O(FE_PHN585_n931), 
	.I(n931));
   DELDKHD FE_PHC584_n3386 (.O(FE_PHN584_n3386), 
	.I(n3386));
   DELDKHD FE_PHC583_n3887 (.O(FE_PHN583_n3887), 
	.I(n3887));
   DELDKHD FE_PHC582_n1878 (.O(FE_PHN582_n1878), 
	.I(n1878));
   DELDKHD FE_PHC581_n2826 (.O(FE_PHN581_n2826), 
	.I(n2826));
   DELDKHD FE_PHC580_n1186 (.O(FE_PHN580_n1186), 
	.I(n1186));
   DELDKHD FE_PHC579_n3510 (.O(FE_PHN579_n3510), 
	.I(n3510));
   DELDKHD FE_PHC578_n3781 (.O(FE_PHN578_n3781), 
	.I(n3781));
   DELDKHD FE_PHC577_n3800 (.O(FE_PHN577_n3800), 
	.I(n3800));
   DELDKHD FE_PHC576_n4296 (.O(FE_PHN576_n4296), 
	.I(n4296));
   DELDKHD FE_PHC575_n2683 (.O(FE_PHN575_n2683), 
	.I(n2683));
   DELDKHD FE_PHC574_n740 (.O(FE_PHN574_n740), 
	.I(n740));
   DELDKHD FE_PHC573_n3246 (.O(FE_PHN573_n3246), 
	.I(n3246));
   DELDKHD FE_PHC572_n1085 (.O(FE_PHN572_n1085), 
	.I(n1085));
   DELDKHD FE_PHC571_n3560 (.O(FE_PHN571_n3560), 
	.I(n3560));
   DELDKHD FE_PHC570_n3868 (.O(FE_PHN570_n3868), 
	.I(n3868));
   DELDKHD FE_PHC569_n3537 (.O(FE_PHN569_n3537), 
	.I(n3537));
   DELDKHD FE_PHC568_n4440 (.O(FE_PHN568_n4440), 
	.I(n4440));
   DELDKHD FE_PHC567_n4604 (.O(FE_PHN567_n4604), 
	.I(n4604));
   DELDKHD FE_PHC566_n1616 (.O(FE_PHN566_n1616), 
	.I(n1616));
   DELDKHD FE_PHC565_n2583 (.O(FE_PHN565_n2583), 
	.I(n2583));
   DELDKHD FE_PHC564_n753 (.O(FE_PHN564_n753), 
	.I(n753));
   DELDKHD FE_PHC563_n2691 (.O(FE_PHN563_n2691), 
	.I(n2691));
   DELDKHD FE_PHC562_n3470 (.O(FE_PHN562_n3470), 
	.I(n3470));
   DELDKHD FE_PHC561_n3472 (.O(FE_PHN561_n3472), 
	.I(n3472));
   DELDKHD FE_PHC560_n3694 (.O(FE_PHN560_n3694), 
	.I(n3694));
   DELDKHD FE_PHC559_n1656 (.O(FE_PHN559_n1656), 
	.I(n1656));
   DELDKHD FE_PHC558_n3209 (.O(FE_PHN558_n3209), 
	.I(n3209));
   DELDKHD FE_PHC557_n4130 (.O(FE_PHN557_n4130), 
	.I(n4130));
   DELCKHD FE_PHC556_n2667 (.O(FE_PHN556_n2667), 
	.I(n2667));
   DELCKHD FE_PHC555_n4448 (.O(FE_PHN555_n4448), 
	.I(n4448));
   DELCKHD FE_PHC554_n2786 (.O(FE_PHN554_n2786), 
	.I(n2786));
   DELCKHD FE_PHC553_n3358 (.O(FE_PHN553_n3358), 
	.I(n3358));
   DELCKHD FE_PHC552_n802 (.O(FE_PHN552_n802), 
	.I(n802));
   DELCKHD FE_PHC551_n734 (.O(FE_PHN551_n734), 
	.I(n734));
   DELCKHD FE_PHC550_n3819 (.O(FE_PHN550_n3819), 
	.I(n3819));
   DELCKHD FE_PHC549_n4461 (.O(FE_PHN549_n4461), 
	.I(n4461));
   DELCKHD FE_PHC548_n3746 (.O(FE_PHN548_n3746), 
	.I(n3746));
   DELCKHD FE_PHC547_n3763 (.O(FE_PHN547_n3763), 
	.I(n3763));
   DELCKHD FE_PHC546_n793 (.O(FE_PHN546_n793), 
	.I(n793));
   DELCKHD FE_PHC545_n1790 (.O(FE_PHN545_n1790), 
	.I(n1790));
   DELCKHD FE_PHC544_n2183 (.O(FE_PHN544_n2183), 
	.I(n2183));
   DELCKHD FE_PHC543_n1690 (.O(FE_PHN543_n1690), 
	.I(n1690));
   DELCKHD FE_PHC542_n4553 (.O(FE_PHN542_n4553), 
	.I(n4553));
   DELCKHD FE_PHC541_n4044 (.O(FE_PHN541_n4044), 
	.I(n4044));
   DELCKHD FE_PHC540_n2942 (.O(FE_PHN540_n2942), 
	.I(n2942));
   DELCKHD FE_PHC539_n3881 (.O(FE_PHN539_n3881), 
	.I(n3881));
   DELCKHD FE_PHC538_n1735 (.O(FE_PHN538_n1735), 
	.I(n1735));
   DELCKHD FE_PHC537_n4622 (.O(FE_PHN537_n4622), 
	.I(n4622));
   DELCKHD FE_PHC536_n1611 (.O(FE_PHN536_n1611), 
	.I(n1611));
   DELCKHD FE_PHC535_n2839 (.O(FE_PHN535_n2839), 
	.I(n2839));
   DELCKHD FE_PHC534_n4118 (.O(FE_PHN534_n4118), 
	.I(n4118));
   DELCKHD FE_PHC533_n2744 (.O(FE_PHN533_n2744), 
	.I(n2744));
   DELCKHD FE_PHC532_n3329 (.O(FE_PHN532_n3329), 
	.I(n3329));
   DELCKHD FE_PHC531_n2354 (.O(FE_PHN531_n2354), 
	.I(n2354));
   DELCKHD FE_PHC530_n3742 (.O(FE_PHN530_n3742), 
	.I(n3742));
   DELCKHD FE_PHC529_n1957 (.O(FE_PHN529_n1957), 
	.I(n1957));
   DELCKHD FE_PHC528_n610 (.O(FE_PHN528_n610), 
	.I(n610));
   DELCKHD FE_PHC527_n1577 (.O(FE_PHN527_n1577), 
	.I(n1577));
   DELCKHD FE_PHC526_n2185 (.O(FE_PHN526_n2185), 
	.I(n2185));
   DELCKHD FE_PHC525_n2017 (.O(FE_PHN525_n2017), 
	.I(n2017));
   DELCKHD FE_PHC524_n2937 (.O(FE_PHN524_n2937), 
	.I(n2937));
   DELCKHD FE_PHC523_n1076 (.O(FE_PHN523_n1076), 
	.I(n1076));
   DELCKHD FE_PHC522_n2633 (.O(FE_PHN522_n2633), 
	.I(n2633));
   DELCKHD FE_PHC521_n3169 (.O(FE_PHN521_n3169), 
	.I(n3169));
   DELCKHD FE_PHC520_n3463 (.O(FE_PHN520_n3463), 
	.I(n3463));
   DELCKHD FE_PHC519_n1562 (.O(FE_PHN519_n1562), 
	.I(n1562));
   DELCKHD FE_PHC518_n4070 (.O(FE_PHN518_n4070), 
	.I(n4070));
   DELCKHD FE_PHC517_n3364 (.O(FE_PHN517_n3364), 
	.I(n3364));
   DELCKHD FE_PHC516_ram_29__14_ (.O(FE_PHN516_ram_29__14_), 
	.I(\ram[29][14] ));
   DELCKHD FE_PHC515_n3497 (.O(FE_PHN515_n3497), 
	.I(n3497));
   DELCKHD FE_PHC514_n3295 (.O(FE_PHN514_n3295), 
	.I(n3295));
   DELCKHD FE_PHC513_n4603 (.O(FE_PHN513_n4603), 
	.I(n4603));
   DELCKHD FE_PHC512_n736 (.O(FE_PHN512_n736), 
	.I(n736));
   DELCKHD FE_PHC511_n3838 (.O(FE_PHN511_n3838), 
	.I(n3838));
   DELCKHD FE_PHC510_n1443 (.O(FE_PHN510_n1443), 
	.I(n1443));
   DELCKHD FE_PHC509_n1055 (.O(FE_PHN509_n1055), 
	.I(n1055));
   DELCKHD FE_PHC508_n3323 (.O(FE_PHN508_n3323), 
	.I(n3323));
   DELCKHD FE_PHC507_n4441 (.O(FE_PHN507_n4441), 
	.I(n4441));
   DELCKHD FE_PHC506_n1700 (.O(FE_PHN506_n1700), 
	.I(n1700));
   DELCKHD FE_PHC505_n1816 (.O(FE_PHN505_n1816), 
	.I(n1816));
   DELCKHD FE_PHC504_n3337 (.O(FE_PHN504_n3337), 
	.I(n3337));
   DELCKHD FE_PHC503_n3676 (.O(FE_PHN503_n3676), 
	.I(n3676));
   DELCKHD FE_PHC502_n3327 (.O(FE_PHN502_n3327), 
	.I(n3327));
   DELCKHD FE_PHC501_n2456 (.O(FE_PHN501_n2456), 
	.I(n2456));
   DELCKHD FE_PHC500_n4275 (.O(FE_PHN500_n4275), 
	.I(n4275));
   DELCKHD FE_PHC499_n4609 (.O(FE_PHN499_n4609), 
	.I(n4609));
   DELCKHD FE_PHC498_n2948 (.O(FE_PHN498_n2948), 
	.I(n2948));
   DELCKHD FE_PHC497_n2915 (.O(FE_PHN497_n2915), 
	.I(n2915));
   DELCKHD FE_PHC496_n2718 (.O(FE_PHN496_n2718), 
	.I(n2718));
   DELCKHD FE_PHC495_n743 (.O(FE_PHN495_n743), 
	.I(n743));
   DELCKHD FE_PHC494_n4435 (.O(FE_PHN494_n4435), 
	.I(n4435));
   DELCKHD FE_PHC493_n4319 (.O(FE_PHN493_n4319), 
	.I(n4319));
   DELCKHD FE_PHC492_n4352 (.O(FE_PHN492_n4352), 
	.I(n4352));
   DELCKHD FE_PHC491_n1948 (.O(FE_PHN491_n1948), 
	.I(n1948));
   DELCKHD FE_PHC490_n2654 (.O(FE_PHN490_n2654), 
	.I(n2654));
   DELCKHD FE_PHC489_n3534 (.O(FE_PHN489_n3534), 
	.I(n3534));
   DELCKHD FE_PHC488_n3512 (.O(FE_PHN488_n3512), 
	.I(n3512));
   DELCKHD FE_PHC487_n3555 (.O(FE_PHN487_n3555), 
	.I(n3555));
   DELCKHD FE_PHC486_n3473 (.O(FE_PHN486_n3473), 
	.I(n3473));
   DELCKHD FE_PHC485_n4644 (.O(FE_PHN485_n4644), 
	.I(n4644));
   DELCKHD FE_PHC484_n3570 (.O(FE_PHN484_n3570), 
	.I(n3570));
   DELCKHD FE_PHC483_n3274 (.O(FE_PHN483_n3274), 
	.I(n3274));
   DELCKHD FE_PHC482_n3389 (.O(FE_PHN482_n3389), 
	.I(n3389));
   DELCKHD FE_PHC481_n4567 (.O(FE_PHN481_n4567), 
	.I(n4567));
   DELCKHD FE_PHC480_n1765 (.O(FE_PHN480_n1765), 
	.I(n1765));
   DELCKHD FE_PHC479_n2204 (.O(FE_PHN479_n2204), 
	.I(n2204));
   DELCKHD FE_PHC478_n4548 (.O(FE_PHN478_n4548), 
	.I(n4548));
   DELCKHD FE_PHC477_n2277 (.O(FE_PHN477_n2277), 
	.I(n2277));
   DELCKHD FE_PHC476_n2349 (.O(FE_PHN476_n2349), 
	.I(n2349));
   DELCKHD FE_PHC475_n2648 (.O(FE_PHN475_n2648), 
	.I(n2648));
   DELCKHD FE_PHC474_n4574 (.O(FE_PHN474_n4574), 
	.I(n4574));
   DELCKHD FE_PHC473_n2789 (.O(FE_PHN473_n2789), 
	.I(n2789));
   DELCKHD FE_PHC472_n3928 (.O(FE_PHN472_n3928), 
	.I(n3928));
   DELCKHD FE_PHC471_n4297 (.O(FE_PHN471_n4297), 
	.I(n4297));
   DELCKHD FE_PHC470_n1686 (.O(FE_PHN470_n1686), 
	.I(n1686));
   DELCKHD FE_PHC469_n4125 (.O(FE_PHN469_n4125), 
	.I(n4125));
   DELCKHD FE_PHC468_n1764 (.O(FE_PHN468_n1764), 
	.I(n1764));
   DELCKHD FE_PHC467_n2818 (.O(FE_PHN467_n2818), 
	.I(n2818));
   DELCKHD FE_PHC466_n3862 (.O(FE_PHN466_n3862), 
	.I(n3862));
   DELCKHD FE_PHC465_n769 (.O(FE_PHN465_n769), 
	.I(n769));
   DELCKHD FE_PHC464_n2254 (.O(FE_PHN464_n2254), 
	.I(n2254));
   DELCKHD FE_PHC463_n2765 (.O(FE_PHN463_n2765), 
	.I(n2765));
   DELCKHD FE_PHC462_n2348 (.O(FE_PHN462_n2348), 
	.I(n2348));
   DELCKHD FE_PHC461_n3842 (.O(FE_PHN461_n3842), 
	.I(n3842));
   DELCKHD FE_PHC460_n3912 (.O(FE_PHN460_n3912), 
	.I(n3912));
   DELCKHD FE_PHC459_n3375 (.O(FE_PHN459_n3375), 
	.I(n3375));
   DELCKHD FE_PHC458_n3877 (.O(FE_PHN458_n3877), 
	.I(n3877));
   DELCKHD FE_PHC457_n1137 (.O(FE_PHN457_n1137), 
	.I(n1137));
   DELCKHD FE_PHC456_n4129 (.O(FE_PHN456_n4129), 
	.I(n4129));
   DELCKHD FE_PHC455_n4493 (.O(FE_PHN455_n4493), 
	.I(n4493));
   DELCKHD FE_PHC454_n4282 (.O(FE_PHN454_n4282), 
	.I(n4282));
   DELCKHD FE_PHC453_n4632 (.O(FE_PHN453_n4632), 
	.I(n4632));
   DELCKHD FE_PHC452_n4589 (.O(FE_PHN452_n4589), 
	.I(n4589));
   DELCKHD FE_PHC451_n3798 (.O(FE_PHN451_n3798), 
	.I(n3798));
   DELCKHD FE_PHC450_n3362 (.O(FE_PHN450_n3362), 
	.I(n3362));
   DELCKHD FE_PHC449_n1059 (.O(FE_PHN449_n1059), 
	.I(n1059));
   DELCKHD FE_PHC448_n4565 (.O(FE_PHN448_n4565), 
	.I(n4565));
   DELCKHD FE_PHC447_n2714 (.O(FE_PHN447_n2714), 
	.I(n2714));
   DELCKHD FE_PHC446_n3579 (.O(FE_PHN446_n3579), 
	.I(n3579));
   DELCKHD FE_PHC445_n3810 (.O(FE_PHN445_n3810), 
	.I(n3810));
   DELCKHD FE_PHC444_n4602 (.O(FE_PHN444_n4602), 
	.I(n4602));
   DELCKHD FE_PHC443_n2711 (.O(FE_PHN443_n2711), 
	.I(n2711));
   DELCKHD FE_PHC442_n2205 (.O(FE_PHN442_n2205), 
	.I(n2205));
   DELCKHD FE_PHC441_n4527 (.O(FE_PHN441_n4527), 
	.I(n4527));
   DELCKHD FE_PHC440_n4503 (.O(FE_PHN440_n4503), 
	.I(n4503));
   DELCKHD FE_PHC439_n4106 (.O(FE_PHN439_n4106), 
	.I(n4106));
   DELCKHD FE_PHC438_n3633 (.O(FE_PHN438_n3633), 
	.I(n3633));
   DELCKHD FE_PHC437_n4508 (.O(FE_PHN437_n4508), 
	.I(n4508));
   DELCKHD FE_PHC436_n1406 (.O(FE_PHN436_n1406), 
	.I(n1406));
   DELCKHD FE_PHC435_n2071 (.O(FE_PHN435_n2071), 
	.I(n2071));
   DELDKHD FE_PHC434_n4471 (.O(FE_PHN434_n4471), 
	.I(n4471));
   DELDKHD FE_PHC433_n3888 (.O(FE_PHN433_n3888), 
	.I(n3888));
   DELDKHD FE_PHC432_n4512 (.O(FE_PHN432_n4512), 
	.I(n4512));
   DELDKHD FE_PHC431_n4054 (.O(FE_PHN431_n4054), 
	.I(n4054));
   DELDKHD FE_PHC430_n2236 (.O(FE_PHN430_n2236), 
	.I(n2236));
   DELDKHD FE_PHC429_n1644 (.O(FE_PHN429_n1644), 
	.I(n1644));
   DELDKHD FE_PHC428_n2365 (.O(FE_PHN428_n2365), 
	.I(n2365));
   DELDKHD FE_PHC427_n2531 (.O(FE_PHN427_n2531), 
	.I(n2531));
   DELDKHD FE_PHC426_n2637 (.O(FE_PHN426_n2637), 
	.I(n2637));
   DELDKHD FE_PHC425_n2274 (.O(FE_PHN425_n2274), 
	.I(n2274));
   DELDKHD FE_PHC424_n867 (.O(FE_PHN424_n867), 
	.I(n867));
   DELDKHD FE_PHC423_n990 (.O(FE_PHN423_n990), 
	.I(n990));
   DELDKHD FE_PHC422_n1710 (.O(FE_PHN422_n1710), 
	.I(n1710));
   DELDKHD FE_PHC421_n2356 (.O(FE_PHN421_n2356), 
	.I(n2356));
   DELDKHD FE_PHC420_n737 (.O(FE_PHN420_n737), 
	.I(n737));
   DELDKHD FE_PHC419_n3757 (.O(FE_PHN419_n3757), 
	.I(n3757));
   DELDKHD FE_PHC418_n2465 (.O(FE_PHN418_n2465), 
	.I(n2465));
   DELDKHD FE_PHC417_n1802 (.O(FE_PHN417_n1802), 
	.I(n1802));
   DELDKHD FE_PHC416_n862 (.O(FE_PHN416_n862), 
	.I(n862));
   DELDKHD FE_PHC415_n2299 (.O(FE_PHN415_n2299), 
	.I(n2299));
   DELDKHD FE_PHC414_n3156 (.O(FE_PHN414_n3156), 
	.I(n3156));
   DELDKHD FE_PHC413_n3625 (.O(FE_PHN413_n3625), 
	.I(n3625));
   DELDKHD FE_PHC412_n4566 (.O(FE_PHN412_n4566), 
	.I(n4566));
   DELDKHD FE_PHC411_n4635 (.O(FE_PHN411_n4635), 
	.I(n4635));
   DELDKHD FE_PHC410_n2032 (.O(FE_PHN410_n2032), 
	.I(n2032));
   DELDKHD FE_PHC409_n2361 (.O(FE_PHN409_n2361), 
	.I(n2361));
   DELDKHD FE_PHC408_n2435 (.O(FE_PHN408_n2435), 
	.I(n2435));
   DELDKHD FE_PHC407_n3670 (.O(FE_PHN407_n3670), 
	.I(n3670));
   DELDKHD FE_PHC406_n796 (.O(FE_PHN406_n796), 
	.I(n796));
   DELDKHD FE_PHC405_n3679 (.O(FE_PHN405_n3679), 
	.I(n3679));
   DELDKHD FE_PHC404_n1525 (.O(FE_PHN404_n1525), 
	.I(n1525));
   DELDKHD FE_PHC403_n3526 (.O(FE_PHN403_n3526), 
	.I(n3526));
   DELDKHD FE_PHC402_n1694 (.O(FE_PHN402_n1694), 
	.I(n1694));
   DELDKHD FE_PHC401_n804 (.O(FE_PHN401_n804), 
	.I(n804));
   DELDKHD FE_PHC400_n2245 (.O(FE_PHN400_n2245), 
	.I(n2245));
   DELDKHD FE_PHC399_n609 (.O(FE_PHN399_n609), 
	.I(n609));
   DELDKHD FE_PHC398_n2720 (.O(FE_PHN398_n2720), 
	.I(n2720));
   DELDKHD FE_PHC397_n1392 (.O(FE_PHN397_n1392), 
	.I(n1392));
   DELDKHD FE_PHC396_n1956 (.O(FE_PHN396_n1956), 
	.I(n1956));
   DELDKHD FE_PHC395_n2521 (.O(FE_PHN395_n2521), 
	.I(n2521));
   DELDKHD FE_PHC394_n4571 (.O(FE_PHN394_n4571), 
	.I(n4571));
   DELDKHD FE_PHC393_n1813 (.O(FE_PHN393_n1813), 
	.I(n1813));
   DELDKHD FE_PHC392_n2770 (.O(FE_PHN392_n2770), 
	.I(n2770));
   DELDKHD FE_PHC391_n2146 (.O(FE_PHN391_n2146), 
	.I(n2146));
   DELDKHD FE_PHC390_n3166 (.O(FE_PHN390_n3166), 
	.I(n3166));
   DELDKHD FE_PHC389_n1730 (.O(FE_PHN389_n1730), 
	.I(n1730));
   DELDKHD FE_PHC388_n1770 (.O(FE_PHN388_n1770), 
	.I(n1770));
   DELDKHD FE_PHC387_n4525 (.O(FE_PHN387_n4525), 
	.I(n4525));
   DELDKHD FE_PHC386_n4475 (.O(FE_PHN386_n4475), 
	.I(n4475));
   DELDKHD FE_PHC385_n2715 (.O(FE_PHN385_n2715), 
	.I(n2715));
   DELDKHD FE_PHC384_n2841 (.O(FE_PHN384_n2841), 
	.I(n2841));
   DELDKHD FE_PHC383_n3677 (.O(FE_PHN383_n3677), 
	.I(n3677));
   DELDKHD FE_PHC382_n3762 (.O(FE_PHN382_n3762), 
	.I(n3762));
   DELDKHD FE_PHC381_n3749 (.O(FE_PHN381_n3749), 
	.I(n3749));
   DELDKHD FE_PHC380_n1707 (.O(FE_PHN380_n1707), 
	.I(n1707));
   DELDKHD FE_PHC379_n3367 (.O(FE_PHN379_n3367), 
	.I(n3367));
   DELDKHD FE_PHC378_n1708 (.O(FE_PHN378_n1708), 
	.I(n1708));
   DELDKHD FE_PHC377_n1194 (.O(FE_PHN377_n1194), 
	.I(n1194));
   DELDKHD FE_PHC376_n601 (.O(FE_PHN376_n601), 
	.I(n601));
   DELDKHD FE_PHC375_n2337 (.O(FE_PHN375_n2337), 
	.I(n2337));
   DELDKHD FE_PHC374_n4246 (.O(FE_PHN374_n4246), 
	.I(n4246));
   DELDKHD FE_PHC373_n2779 (.O(FE_PHN373_n2779), 
	.I(n2779));
   DELDKHD FE_PHC372_n797 (.O(FE_PHN372_n797), 
	.I(n797));
   DELDKHD FE_PHC371_n4494 (.O(FE_PHN371_n4494), 
	.I(n4494));
   DELDKHD FE_PHC370_n3629 (.O(FE_PHN370_n3629), 
	.I(n3629));
   DELDKHD FE_PHC369_n4579 (.O(FE_PHN369_n4579), 
	.I(n4579));
   DELDKHD FE_PHC368_n4580 (.O(FE_PHN368_n4580), 
	.I(n4580));
   DELDKHD FE_PHC367_n4449 (.O(FE_PHN367_n4449), 
	.I(n4449));
   DELDKHD FE_PHC366_n4193 (.O(FE_PHN366_n4193), 
	.I(n4193));
   DELDKHD FE_PHC365_n987 (.O(FE_PHN365_n987), 
	.I(n987));
   DELDKHD FE_PHC364_n3236 (.O(FE_PHN364_n3236), 
	.I(n3236));
   DELDKHD FE_PHC363_n1509 (.O(FE_PHN363_n1509), 
	.I(n1509));
   DELDKHD FE_PHC362_n1711 (.O(FE_PHN362_n1711), 
	.I(n1711));
   DELDKHD FE_PHC361_n1065 (.O(FE_PHN361_n1065), 
	.I(n1065));
   DELDKHD FE_PHC360_n1330 (.O(FE_PHN360_n1330), 
	.I(n1330));
   DELDKHD FE_PHC359_n3531 (.O(FE_PHN359_n3531), 
	.I(n3531));
   DELDKHD FE_PHC358_n4326 (.O(FE_PHN358_n4326), 
	.I(n4326));
   DELDKHD FE_PHC357_n2473 (.O(FE_PHN357_n2473), 
	.I(n2473));
   DELDKHD FE_PHC356_n1653 (.O(FE_PHN356_n1653), 
	.I(n1653));
   DELDKHD FE_PHC355_n3354 (.O(FE_PHN355_n3354), 
	.I(n3354));
   DELDKHD FE_PHC354_n4581 (.O(FE_PHN354_n4581), 
	.I(n4581));
   DELDKHD FE_PHC353_n3608 (.O(FE_PHN353_n3608), 
	.I(n3608));
   DELDKHD FE_PHC352_n1063 (.O(FE_PHN352_n1063), 
	.I(n1063));
   DELDKHD FE_PHC351_n2647 (.O(FE_PHN351_n2647), 
	.I(n2647));
   DELDKHD FE_PHC350_n3805 (.O(FE_PHN350_n3805), 
	.I(n3805));
   DELDKHD FE_PHC349_n2294 (.O(FE_PHN349_n2294), 
	.I(n2294));
   DELDKHD FE_PHC348_n4474 (.O(FE_PHN348_n4474), 
	.I(n4474));
   DELDKHD FE_PHC347_n1792 (.O(FE_PHN347_n1792), 
	.I(n1792));
   DELDKHD FE_PHC346_n2801 (.O(FE_PHN346_n2801), 
	.I(n2801));
   DELDKHD FE_PHC345_n4257 (.O(FE_PHN345_n4257), 
	.I(n4257));
   DELDKHD FE_PHC344_n2787 (.O(FE_PHN344_n2787), 
	.I(n2787));
   DELDKHD FE_PHC343_n3165 (.O(FE_PHN343_n3165), 
	.I(n3165));
   DELDKHD FE_PHC342_n3233 (.O(FE_PHN342_n3233), 
	.I(n3233));
   DELDKHD FE_PHC341_n3743 (.O(FE_PHN341_n3743), 
	.I(n3743));
   DELDKHD FE_PHC340_n4038 (.O(FE_PHN340_n4038), 
	.I(n4038));
   DELDKHD FE_PHC339_n4613 (.O(FE_PHN339_n4613), 
	.I(n4613));
   DELDKHD FE_PHC338_n3783 (.O(FE_PHN338_n3783), 
	.I(n3783));
   DELDKHD FE_PHC337_n4318 (.O(FE_PHN337_n4318), 
	.I(n4318));
   DELDKHD FE_PHC336_n915 (.O(FE_PHN336_n915), 
	.I(n915));
   DELDKHD FE_PHC335_n1622 (.O(FE_PHN335_n1622), 
	.I(n1622));
   DELDKHD FE_PHC334_n2343 (.O(FE_PHN334_n2343), 
	.I(n2343));
   DELDKHD FE_PHC333_n3490 (.O(FE_PHN333_n3490), 
	.I(n3490));
   DELDKHD FE_PHC332_n3967 (.O(FE_PHN332_n3967), 
	.I(n3967));
   DELCKHD FE_PHC331_n3574 (.O(FE_PHN331_n3574), 
	.I(n3574));
   DELCKHD FE_PHC330_n2728 (.O(FE_PHN330_n2728), 
	.I(n2728));
   DELCKHD FE_PHC329_n3355 (.O(FE_PHN329_n3355), 
	.I(n3355));
   DELCKHD FE_PHC328_n3678 (.O(FE_PHN328_n3678), 
	.I(n3678));
   DELCKHD FE_PHC327_n3857 (.O(FE_PHN327_n3857), 
	.I(n3857));
   DELCKHD FE_PHC326_n4325 (.O(FE_PHN326_n4325), 
	.I(n4325));
   DELCKHD FE_PHC325_n3484 (.O(FE_PHN325_n3484), 
	.I(n3484));
   DELCKHD FE_PHC324_n3748 (.O(FE_PHN324_n3748), 
	.I(n3748));
   DELCKHD FE_PHC323_n3489 (.O(FE_PHN323_n3489), 
	.I(n3489));
   DELCKHD FE_PHC322_n1624 (.O(FE_PHN322_n1624), 
	.I(n1624));
   DELCKHD FE_PHC321_n2392 (.O(FE_PHN321_n2392), 
	.I(n2392));
   DELCKHD FE_PHC320_n4256 (.O(FE_PHN320_n4256), 
	.I(n4256));
   DELCKHD FE_PHC319_n3532 (.O(FE_PHN319_n3532), 
	.I(n3532));
   DELCKHD FE_PHC318_n1945 (.O(FE_PHN318_n1945), 
	.I(n1945));
   DELCKHD FE_PHC317_n4310 (.O(FE_PHN317_n4310), 
	.I(n4310));
   DELCKHD FE_PHC316_n1782 (.O(FE_PHN316_n1782), 
	.I(n1782));
   DELCKHD FE_PHC315_n3768 (.O(FE_PHN315_n3768), 
	.I(n3768));
   DELCKHD FE_PHC314_n3861 (.O(FE_PHN314_n3861), 
	.I(n3861));
   DELCKHD FE_PHC313_n4479 (.O(FE_PHN313_n4479), 
	.I(n4479));
   DELCKHD FE_PHC312_n4502 (.O(FE_PHN312_n4502), 
	.I(n4502));
   DELCKHD FE_PHC311_n1010 (.O(FE_PHN311_n1010), 
	.I(n1010));
   DELCKHD FE_PHC310_n2901 (.O(FE_PHN310_n2901), 
	.I(n2901));
   DELCKHD FE_PHC309_n4328 (.O(FE_PHN309_n4328), 
	.I(n4328));
   DELCKHD FE_PHC308_n2140 (.O(FE_PHN308_n2140), 
	.I(n2140));
   DELCKHD FE_PHC307_n2157 (.O(FE_PHN307_n2157), 
	.I(n2157));
   DELCKHD FE_PHC306_n2341 (.O(FE_PHN306_n2341), 
	.I(n2341));
   DELCKHD FE_PHC305_n3536 (.O(FE_PHN305_n3536), 
	.I(n3536));
   DELCKHD FE_PHC304_n3562 (.O(FE_PHN304_n3562), 
	.I(n3562));
   DELCKHD FE_PHC303_n2778 (.O(FE_PHN303_n2778), 
	.I(n2778));
   DELCKHD FE_PHC302_n4065 (.O(FE_PHN302_n4065), 
	.I(n4065));
   DELCKHD FE_PHC301_n3730 (.O(FE_PHN301_n3730), 
	.I(n3730));
   DELCKHD FE_PHC300_n4515 (.O(FE_PHN300_n4515), 
	.I(n4515));
   DELCKHD FE_PHC299_n2134 (.O(FE_PHN299_n2134), 
	.I(n2134));
   DELCKHD FE_PHC298_n1817 (.O(FE_PHN298_n1817), 
	.I(n1817));
   DELCKHD FE_PHC297_n2540 (.O(FE_PHN297_n2540), 
	.I(n2540));
   DELCKHD FE_PHC296_n3508 (.O(FE_PHN296_n3508), 
	.I(n3508));
   DELCKHD FE_PHC295_n4120 (.O(FE_PHN295_n4120), 
	.I(n4120));
   DELCKHD FE_PHC294_n1047 (.O(FE_PHN294_n1047), 
	.I(n1047));
   DELCKHD FE_PHC293_n2523 (.O(FE_PHN293_n2523), 
	.I(n2523));
   DELCKHD FE_PHC292_n2489 (.O(FE_PHN292_n2489), 
	.I(n2489));
   DELCKHD FE_PHC291_n4465 (.O(FE_PHN291_n4465), 
	.I(n4465));
   DELCKHD FE_PHC290_n1369 (.O(FE_PHN290_n1369), 
	.I(n1369));
   DELCKHD FE_PHC289_n3935 (.O(FE_PHN289_n3935), 
	.I(n3935));
   DELCKHD FE_PHC288_n4186 (.O(FE_PHN288_n4186), 
	.I(n4186));
   DELCKHD FE_PHC287_n4658 (.O(FE_PHN287_n4658), 
	.I(n4658));
   DELCKHD FE_PHC286_n3957 (.O(FE_PHN286_n3957), 
	.I(n3957));
   DELCKHD FE_PHC285_n2200 (.O(FE_PHN285_n2200), 
	.I(n2200));
   DELCKHD FE_PHC284_n2601 (.O(FE_PHN284_n2601), 
	.I(n2601));
   DELCKHD FE_PHC283_n4633 (.O(FE_PHN283_n4633), 
	.I(n4633));
   DELCKHD FE_PHC282_n3557 (.O(FE_PHN282_n3557), 
	.I(n3557));
   DELCKHD FE_PHC281_n4568 (.O(FE_PHN281_n4568), 
	.I(n4568));
   DELCKHD FE_PHC280_n3380 (.O(FE_PHN280_n3380), 
	.I(n3380));
   DELCKHD FE_PHC279_n2162 (.O(FE_PHN279_n2162), 
	.I(n2162));
   DELCKHD FE_PHC278_n3097 (.O(FE_PHN278_n3097), 
	.I(n3097));
   DELCKHD FE_PHC277_n1626 (.O(FE_PHN277_n1626), 
	.I(n1626));
   DELCKHD FE_PHC276_n3544 (.O(FE_PHN276_n3544), 
	.I(n3544));
   DELCKHD FE_PHC275_n1753 (.O(FE_PHN275_n1753), 
	.I(n1753));
   DELCKHD FE_PHC274_n2796 (.O(FE_PHN274_n2796), 
	.I(n2796));
   DELCKHD FE_PHC273_n4081 (.O(FE_PHN273_n4081), 
	.I(n4081));
   DELCKHD FE_PHC272_n4533 (.O(FE_PHN272_n4533), 
	.I(n4533));
   DELCKHD FE_PHC271_n2278 (.O(FE_PHN271_n2278), 
	.I(n2278));
   DELCKHD FE_PHC270_n2467 (.O(FE_PHN270_n2467), 
	.I(n2467));
   DELCKHD FE_PHC269_n2340 (.O(FE_PHN269_n2340), 
	.I(n2340));
   DELCKHD FE_PHC268_n1061 (.O(FE_PHN268_n1061), 
	.I(n1061));
   DELCKHD FE_PHC267_n1373 (.O(FE_PHN267_n1373), 
	.I(n1373));
   DELCKHD FE_PHC266_n3611 (.O(FE_PHN266_n3611), 
	.I(n3611));
   DELCKHD FE_PHC265_n3772 (.O(FE_PHN265_n3772), 
	.I(n3772));
   DELCKHD FE_PHC264_n2409 (.O(FE_PHN264_n2409), 
	.I(n2409));
   DELCKHD FE_PHC263_n4477 (.O(FE_PHN263_n4477), 
	.I(n4477));
   DELCKHD FE_PHC262_n3350 (.O(FE_PHN262_n3350), 
	.I(n3350));
   DELCKHD FE_PHC261_n2201 (.O(FE_PHN261_n2201), 
	.I(n2201));
   DELCKHD FE_PHC260_n2761 (.O(FE_PHN260_n2761), 
	.I(n2761));
   DELCKHD FE_PHC259_n1508 (.O(FE_PHN259_n1508), 
	.I(n1508));
   DELCKHD FE_PHC258_n1814 (.O(FE_PHN258_n1814), 
	.I(n1814));
   DELCKHD FE_PHC257_n3817 (.O(FE_PHN257_n3817), 
	.I(n3817));
   DELCKHD FE_PHC256_n1146 (.O(FE_PHN256_n1146), 
	.I(n1146));
   DELCKHD FE_PHC255_n1781 (.O(FE_PHN255_n1781), 
	.I(n1781));
   DELCKHD FE_PHC254_n3231 (.O(FE_PHN254_n3231), 
	.I(n3231));
   DELCKHD FE_PHC253_n3986 (.O(FE_PHN253_n3986), 
	.I(n3986));
   DELDKHD FE_PHC252_n2455 (.O(FE_PHN252_n2455), 
	.I(n2455));
   DELDKHD FE_PHC251_n1691 (.O(FE_PHN251_n1691), 
	.I(n1691));
   DELDKHD FE_PHC250_n4024 (.O(FE_PHN250_n4024), 
	.I(n4024));
   DELDKHD FE_PHC249_n2461 (.O(FE_PHN249_n2461), 
	.I(n2461));
   DELDKHD FE_PHC248_n3747 (.O(FE_PHN248_n3747), 
	.I(n3747));
   DELDKHD FE_PHC247_n2652 (.O(FE_PHN247_n2652), 
	.I(n2652));
   DELDKHD FE_PHC246_n3172 (.O(FE_PHN246_n3172), 
	.I(n3172));
   DELDKHD FE_PHC245_n763 (.O(FE_PHN245_n763), 
	.I(n763));
   DELDKHD FE_PHC244_n2588 (.O(FE_PHN244_n2588), 
	.I(n2588));
   DELDKHD FE_PHC243_n1795 (.O(FE_PHN243_n1795), 
	.I(n1795));
   DELDKHD FE_PHC242_n2174 (.O(FE_PHN242_n2174), 
	.I(n2174));
   DELDKHD FE_PHC241_n2741 (.O(FE_PHN241_n2741), 
	.I(n2741));
   DELDKHD FE_PHC240_n4247 (.O(FE_PHN240_n4247), 
	.I(n4247));
   DELDKHD FE_PHC239_n4105 (.O(FE_PHN239_n4105), 
	.I(n4105));
   DELDKHD FE_PHC238_n3572 (.O(FE_PHN238_n3572), 
	.I(n3572));
   DELDKHD FE_PHC237_n4317 (.O(FE_PHN237_n4317), 
	.I(n4317));
   DELDKHD FE_PHC236_n3863 (.O(FE_PHN236_n3863), 
	.I(n3863));
   DELDKHD FE_PHC235_n1761 (.O(FE_PHN235_n1761), 
	.I(n1761));
   DELDKHD FE_PHC234_n4191 (.O(FE_PHN234_n4191), 
	.I(n4191));
   DELDKHD FE_PHC233_n4092 (.O(FE_PHN233_n4092), 
	.I(n4092));
   DELDKHD FE_PHC232_n791 (.O(FE_PHN232_n791), 
	.I(n791));
   DELDKHD FE_PHC231_n3991 (.O(FE_PHN231_n3991), 
	.I(n3991));
   DELDKHD FE_PHC230_n3543 (.O(FE_PHN230_n3543), 
	.I(n3543));
   DELDKHD FE_PHC229_n2333 (.O(FE_PHN229_n2333), 
	.I(n2333));
   DELDKHD FE_PHC228_n3632 (.O(FE_PHN228_n3632), 
	.I(n3632));
   DELDKHD FE_PHC227_n4600 (.O(FE_PHN227_n4600), 
	.I(n4600));
   DELDKHD FE_PHC226_n1239 (.O(FE_PHN226_n1239), 
	.I(n1239));
   DELDKHD FE_PHC225_n2212 (.O(FE_PHN225_n2212), 
	.I(n2212));
   DELDKHD FE_PHC224_n3735 (.O(FE_PHN224_n3735), 
	.I(n3735));
   DELDKHD FE_PHC223_n4020 (.O(FE_PHN223_n4020), 
	.I(n4020));
   DELDKHD FE_PHC222_n2803 (.O(FE_PHN222_n2803), 
	.I(n2803));
   DELDKHD FE_PHC221_n2651 (.O(FE_PHN221_n2651), 
	.I(n2651));
   DELDKHD FE_PHC220_n4636 (.O(FE_PHN220_n4636), 
	.I(n4636));
   DELDKHD FE_PHC219_n2805 (.O(FE_PHN219_n2805), 
	.I(n2805));
   DELDKHD FE_PHC218_n3610 (.O(FE_PHN218_n3610), 
	.I(n3610));
   DELDKHD FE_PHC217_n3239 (.O(FE_PHN217_n3239), 
	.I(n3239));
   DELDKHD FE_PHC216_n2266 (.O(FE_PHN216_n2266), 
	.I(n2266));
   DELDKHD FE_PHC215_n3997 (.O(FE_PHN215_n3997), 
	.I(n3997));
   DELDKHD FE_PHC214_n3565 (.O(FE_PHN214_n3565), 
	.I(n3565));
   DELDKHD FE_PHC213_n3170 (.O(FE_PHN213_n3170), 
	.I(n3170));
   DELDKHD FE_PHC212_n4426 (.O(FE_PHN212_n4426), 
	.I(n4426));
   DELDKHD FE_PHC211_n1121 (.O(FE_PHN211_n1121), 
	.I(n1121));
   DELDKHD FE_PHC210_n4132 (.O(FE_PHN210_n4132), 
	.I(n4132));
   DELCKHD FE_PHC209_n3938 (.O(FE_PHN209_n3938), 
	.I(n3938));
   DELCKHD FE_PHC208_n3744 (.O(FE_PHN208_n3744), 
	.I(n3744));
   DELCKHD FE_PHC207_n3673 (.O(FE_PHN207_n3673), 
	.I(n3673));
   DELCKHD FE_PHC206_n1818 (.O(FE_PHN206_n1818), 
	.I(n1818));
   DELCKHD FE_PHC205_n3352 (.O(FE_PHN205_n3352), 
	.I(n3352));
   DELCKHD FE_PHC204_n1754 (.O(FE_PHN204_n1754), 
	.I(n1754));
   DELCKHD FE_PHC203_n1701 (.O(FE_PHN203_n1701), 
	.I(n1701));
   DELCKHD FE_PHC202_n2338 (.O(FE_PHN202_n2338), 
	.I(n2338));
   DELCKHD FE_PHC201_n3990 (.O(FE_PHN201_n3990), 
	.I(n3990));
   DELCKHD FE_PHC200_n4288 (.O(FE_PHN200_n4288), 
	.I(n4288));
   DELCKHD FE_PHC199_n3101 (.O(FE_PHN199_n3101), 
	.I(n3101));
   DELCKHD FE_PHC198_n2208 (.O(FE_PHN198_n2208), 
	.I(n2208));
   DELCKHD FE_PHC197_n4315 (.O(FE_PHN197_n4315), 
	.I(n4315));
   DELCKHD FE_PHC196_n3905 (.O(FE_PHN196_n3905), 
	.I(n3905));
   DELCKHD FE_PHC195_n4587 (.O(FE_PHN195_n4587), 
	.I(n4587));
   DELCKHD FE_PHC194_n2476 (.O(FE_PHN194_n2476), 
	.I(n2476));
   DELCKHD FE_PHC193_n3493 (.O(FE_PHN193_n3493), 
	.I(n3493));
   DELCKHD FE_PHC192_n735 (.O(FE_PHN192_n735), 
	.I(n735));
   DELCKHD FE_PHC191_n3682 (.O(FE_PHN191_n3682), 
	.I(n3682));
   DELCKHD FE_PHC190_n4182 (.O(FE_PHN190_n4182), 
	.I(n4182));
   DELCKHD FE_PHC189_n2712 (.O(FE_PHN189_n2712), 
	.I(n2712));
   DELCKHD FE_PHC188_n3213 (.O(FE_PHN188_n3213), 
	.I(n3213));
   DELCKHD FE_PHC187_n4084 (.O(FE_PHN187_n4084), 
	.I(n4084));
   DELCKHD FE_PHC186_n4320 (.O(FE_PHN186_n4320), 
	.I(n4320));
   DELCKHD FE_PHC185_n4376 (.O(FE_PHN185_n4376), 
	.I(n4376));
   DELCKHD FE_PHC184_n1696 (.O(FE_PHN184_n1696), 
	.I(n1696));
   DELCKHD FE_PHC183_n3491 (.O(FE_PHN183_n3491), 
	.I(n3491));
   DELCKHD FE_PHC182_n1053 (.O(FE_PHN182_n1053), 
	.I(n1053));
   DELCKHD FE_PHC181_n3292 (.O(FE_PHN181_n3292), 
	.I(n3292));
   DELCKHD FE_PHC180_n4456 (.O(FE_PHN180_n4456), 
	.I(n4456));
   DELCKHD FE_PHC179_n3754 (.O(FE_PHN179_n3754), 
	.I(n3754));
   DELCKHD FE_PHC178_n3353 (.O(FE_PHN178_n3353), 
	.I(n3353));
   DELCKHD FE_PHC177_n3300 (.O(FE_PHN177_n3300), 
	.I(n3300));
   DELCKHD FE_PHC176_n1112 (.O(FE_PHN176_n1112), 
	.I(n1112));
   DELCKHD FE_PHC175_n3167 (.O(FE_PHN175_n3167), 
	.I(n3167));
   DELCKHD FE_PHC174_n3734 (.O(FE_PHN174_n3734), 
	.I(n3734));
   DELCKHD FE_PHC173_n4004 (.O(FE_PHN173_n4004), 
	.I(n4004));
   DELCKHD FE_PHC172_n4570 (.O(FE_PHN172_n4570), 
	.I(n4570));
   DELCKHD FE_PHC171_n4190 (.O(FE_PHN171_n4190), 
	.I(n4190));
   DELCKHD FE_PHC170_n3561 (.O(FE_PHN170_n3561), 
	.I(n3561));
   DELCKHD FE_PHC169_n4582 (.O(FE_PHN169_n4582), 
	.I(n4582));
   DELCKHD FE_PHC168_n1435 (.O(FE_PHN168_n1435), 
	.I(n1435));
   DELCKHD FE_PHC167_n3580 (.O(FE_PHN167_n3580), 
	.I(n3580));
   DELCKHD FE_PHC166_n4514 (.O(FE_PHN166_n4514), 
	.I(n4514));
   DELDKHD FE_PHC165_ram_241__1_ (.O(FE_PHN165_ram_241__1_), 
	.I(\ram[241][1] ));
   DELDKHD FE_PHC164_n3164 (.O(FE_PHN164_n3164), 
	.I(n3164));
   DELDKHD FE_PHC163_n2458 (.O(FE_PHN163_n2458), 
	.I(n2458));
   DELDKHD FE_PHC162_n3234 (.O(FE_PHN162_n3234), 
	.I(n3234));
   DELDKHD FE_PHC161_n3548 (.O(FE_PHN161_n3548), 
	.I(n3548));
   DELDKHD FE_PHC160_n3618 (.O(FE_PHN160_n3618), 
	.I(n3618));
   DELDKHD FE_PHC159_n3224 (.O(FE_PHN159_n3224), 
	.I(n3224));
   DELDKHD FE_PHC158_n3563 (.O(FE_PHN158_n3563), 
	.I(n3563));
   DELDKHD FE_PHC157_n3286 (.O(FE_PHN157_n3286), 
	.I(n3286));
   DELDKHD FE_PHC156_n3499 (.O(FE_PHN156_n3499), 
	.I(n3499));
   DELDKHD FE_PHC155_n4055 (.O(FE_PHN155_n4055), 
	.I(n4055));
   DELDKHD FE_PHC154_n3365 (.O(FE_PHN154_n3365), 
	.I(n3365));
   DELDKHD FE_PHC153_n3550 (.O(FE_PHN153_n3550), 
	.I(n3550));
   DELDKHD FE_PHC152_n1049 (.O(FE_PHN152_n1049), 
	.I(n1049));
   DELDKHD FE_PHC151_n1572 (.O(FE_PHN151_n1572), 
	.I(n1572));
   DELDKHD FE_PHC150_n3564 (.O(FE_PHN150_n3564), 
	.I(n3564));
   DELDKHD FE_PHC149_n3621 (.O(FE_PHN149_n3621), 
	.I(n3621));
   DELDKHD FE_PHC148_n4522 (.O(FE_PHN148_n4522), 
	.I(n4522));
   DELDKHD FE_PHC147_n3556 (.O(FE_PHN147_n3556), 
	.I(n3556));
   DELDKHD FE_PHC146_n3609 (.O(FE_PHN146_n3609), 
	.I(n3609));
   DELDKHD FE_PHC145_n2330 (.O(FE_PHN145_n2330), 
	.I(n2330));
   DELDKHD FE_PHC144_n1634 (.O(FE_PHN144_n1634), 
	.I(n1634));
   DELDKHD FE_PHC143_n1704 (.O(FE_PHN143_n1704), 
	.I(n1704));
   DELCKHD FE_PHC142_n3864 (.O(FE_PHN142_n3864), 
	.I(n3864));
   DELCKHD FE_PHC141_n2206 (.O(FE_PHN141_n2206), 
	.I(n2206));
   DELCKHD FE_PHC140_n4313 (.O(FE_PHN140_n4313), 
	.I(n4313));
   DELCKHD FE_PHC139_n4506 (.O(FE_PHN139_n4506), 
	.I(n4506));
   DELCKHD FE_PHC138_n1713 (.O(FE_PHN138_n1713), 
	.I(n1713));
   DELCKHD FE_PHC137_n2142 (.O(FE_PHN137_n2142), 
	.I(n2142));
   DELCKHD FE_PHC136_n4573 (.O(FE_PHN136_n4573), 
	.I(n4573));
   DELCKHD FE_PHC135_n4064 (.O(FE_PHN135_n4064), 
	.I(n4064));
   DELCKHD FE_PHC134_n3606 (.O(FE_PHN134_n3606), 
	.I(n3606));
   DELCKHD FE_PHC133_n2136 (.O(FE_PHN133_n2136), 
	.I(n2136));
   DELCKHD FE_PHC132_n3106 (.O(FE_PHN132_n3106), 
	.I(n3106));
   DELCKHD FE_PHC131_n3870 (.O(FE_PHN131_n3870), 
	.I(n3870));
   DELCKHD FE_PHC130_n4068 (.O(FE_PHN130_n4068), 
	.I(n4068));
   DELCKHD FE_PHC129_n2147 (.O(FE_PHN129_n2147), 
	.I(n2147));
   DELCKHD FE_PHC128_n1695 (.O(FE_PHN128_n1695), 
	.I(n1695));
   DELCKHD FE_PHC127_n4507 (.O(FE_PHN127_n4507), 
	.I(n4507));
   DELCKHD FE_PHC126_n3866 (.O(FE_PHN126_n3866), 
	.I(n3866));
   DELCKHD FE_PHC125_n3546 (.O(FE_PHN125_n3546), 
	.I(n3546));
   DELCKHD FE_PHC124_n2273 (.O(FE_PHN124_n2273), 
	.I(n2273));
   DELCKHD FE_PHC123_n1058 (.O(FE_PHN123_n1058), 
	.I(n1058));
   DELCKHD FE_PHC122_n3226 (.O(FE_PHN122_n3226), 
	.I(n3226));
   DELCKHD FE_PHC121_n3995 (.O(FE_PHN121_n3995), 
	.I(n3995));
   DELCKHD FE_PHC120_n4509 (.O(FE_PHN120_n4509), 
	.I(n4509));
   DELDKHD FE_PHC119_n3538 (.O(FE_PHN119_n3538), 
	.I(n3538));
   DELDKHD FE_PHC118_n4446 (.O(FE_PHN118_n4446), 
	.I(n4446));
   DELDKHD FE_PHC117_n3301 (.O(FE_PHN117_n3301), 
	.I(n3301));
   DELDKHD FE_PHC116_n2207 (.O(FE_PHN116_n2207), 
	.I(n2207));
   DELDKHD FE_PHC115_n3739 (.O(FE_PHN115_n3739), 
	.I(n3739));
   DELDKHD FE_PHC114_n3807 (.O(FE_PHN114_n3807), 
	.I(n3807));
   DELDKHD FE_PHC113_n3533 (.O(FE_PHN113_n3533), 
	.I(n3533));
   DELDKHD FE_PHC112_n4577 (.O(FE_PHN112_n4577), 
	.I(n4577));
   DELDKHD FE_PHC111_n3584 (.O(FE_PHN111_n3584), 
	.I(n3584));
   DELCKHD FE_PHC110_n4504 (.O(FE_PHN110_n4504), 
	.I(n4504));
   DELCKHD FE_PHC109_n3549 (.O(FE_PHN109_n3549), 
	.I(n3549));
   DELCKHD FE_PHC108_n3568 (.O(FE_PHN108_n3568), 
	.I(n3568));
   DELCKHD FE_PHC107_n1692 (.O(FE_PHN107_n1692), 
	.I(n1692));
   DELDKHD FE_PHC106_n3619 (.O(FE_PHN106_n3619), 
	.I(n3619));
   DELDKHD FE_PHC105_n3552 (.O(FE_PHN105_n3552), 
	.I(n3552));
   DELCKHD FE_PHC104_n3545 (.O(FE_PHN104_n3545), 
	.I(n3545));
   DELCKHD FE_PHC103_n3558 (.O(FE_PHN103_n3558), 
	.I(n3558));
   DELCKHD FE_PHC102_n3554 (.O(FE_PHN102_n3554), 
	.I(n3554));
   DELCKHD FE_PHC101_n3547 (.O(FE_PHN101_n3547), 
	.I(n3547));
   DELCKHD FE_PHC100_n3542 (.O(FE_PHN100_n3542), 
	.I(n3542));
   BUFHHD FE_OFC94_mem_write (.O(FE_OFN94_mem_write), 
	.I(mem_write_en));
   BUFHHD FE_OFC93_mem_write (.O(FE_OFN93_mem_write), 
	.I(mem_write_en));
   BUFHHD FE_OFC92_mem_write (.O(FE_OFN92_mem_write), 
	.I(mem_write_en));
   BUFGHD FE_OFC91_n23 (.O(FE_OFN91_n23), 
	.I(FE_OFN89_n23));
   BUFGHD FE_OFC90_n23 (.O(FE_OFN90_n23), 
	.I(n23));
   BUFGHD FE_OFC89_n23 (.O(FE_OFN89_n23), 
	.I(n23));
   BUFGHD FE_OFC88_n22 (.O(FE_OFN88_n22), 
	.I(n22));
   BUFEHD FE_OFC87_n22 (.O(FE_OFN87_n22), 
	.I(FE_OFN86_n22));
   BUFGHD FE_OFC86_n22 (.O(FE_OFN86_n22), 
	.I(n22));
   BUFGHD FE_OFC85_n21 (.O(FE_OFN85_n21), 
	.I(n21));
   BUFEHD FE_OFC84_n21 (.O(FE_OFN84_n21), 
	.I(FE_OFN83_n21));
   BUFGHD FE_OFC83_n21 (.O(FE_OFN83_n21), 
	.I(n21));
   BUFGHD FE_OFC82_n20 (.O(FE_OFN82_n20), 
	.I(FE_OFN79_n20));
   BUFHHD FE_OFC81_n20 (.O(FE_OFN81_n20), 
	.I(FE_OFN79_n20));
   BUFEHD FE_OFC80_n20 (.O(FE_OFN80_n20), 
	.I(FE_OFN79_n20));
   BUFGHD FE_OFC79_n20 (.O(FE_OFN79_n20), 
	.I(n20));
   BUFGHD FE_OFC78_n19 (.O(FE_OFN78_n19), 
	.I(FE_OFN77_n19));
   BUFGHD FE_OFC77_n19 (.O(FE_OFN77_n19), 
	.I(FE_OFN76_n19));
   BUFGHD FE_OFC76_n19 (.O(FE_OFN76_n19), 
	.I(n19));
   BUFGHD FE_OFC75_n18 (.O(FE_OFN75_n18), 
	.I(FE_OFN74_n18));
   BUFGHD FE_OFC74_n18 (.O(FE_OFN74_n18), 
	.I(FE_OFN73_n18));
   BUFGHD FE_OFC73_n18 (.O(FE_OFN73_n18), 
	.I(n18));
   BUFGHD FE_OFC72_n17 (.O(FE_OFN72_n17), 
	.I(FE_OFN71_n17));
   BUFGHD FE_OFC71_n17 (.O(FE_OFN71_n17), 
	.I(FE_OFN70_n17));
   BUFGHD FE_OFC70_n17 (.O(FE_OFN70_n17), 
	.I(n17));
   BUFGHD FE_OFC69_n16 (.O(FE_OFN69_n16), 
	.I(FE_OFN67_n16));
   BUFGHD FE_OFC68_n16 (.O(FE_OFN68_n16), 
	.I(FE_OFN66_n16));
   BUFGHD FE_OFC67_n16 (.O(FE_OFN67_n16), 
	.I(FE_OFN66_n16));
   BUFGHD FE_OFC66_n16 (.O(FE_OFN66_n16), 
	.I(n16));
   BUFGHD FE_OFC65_n15 (.O(FE_OFN65_n15), 
	.I(FE_OFN64_n15));
   BUFGHD FE_OFC64_n15 (.O(FE_OFN64_n15), 
	.I(FE_OFN63_n15));
   BUFGHD FE_OFC63_n15 (.O(FE_OFN63_n15), 
	.I(n15));
   BUFGHD FE_OFC62_n14 (.O(FE_OFN62_n14), 
	.I(FE_OFN61_n14));
   BUFGHD FE_OFC61_n14 (.O(FE_OFN61_n14), 
	.I(n14));
   BUFEHD FE_OFC60_n14 (.O(FE_OFN60_n14), 
	.I(FE_OFN59_n14));
   BUFGHD FE_OFC59_n14 (.O(FE_OFN59_n14), 
	.I(n14));
   BUFGHD FE_OFC58_n13 (.O(FE_OFN58_n13), 
	.I(FE_OFN57_n13));
   BUFGHD FE_OFC57_n13 (.O(FE_OFN57_n13), 
	.I(FE_OFN56_n13));
   BUFGHD FE_OFC56_n13 (.O(FE_OFN56_n13), 
	.I(n13));
   BUFGHD FE_OFC55_n12 (.O(FE_OFN55_n12), 
	.I(FE_OFN53_n12));
   BUFGHD FE_OFC54_n12 (.O(FE_OFN54_n12), 
	.I(n12));
   BUFGHD FE_OFC53_n12 (.O(FE_OFN53_n12), 
	.I(n12));
   BUFGHD FE_OFC52_n11 (.O(FE_OFN52_n11), 
	.I(FE_OFN51_n11));
   BUFGHD FE_OFC51_n11 (.O(FE_OFN51_n11), 
	.I(FE_OFN50_n11));
   BUFGHD FE_OFC50_n11 (.O(FE_OFN50_n11), 
	.I(n11));
   BUFGHD FE_OFC49_n10 (.O(FE_OFN49_n10), 
	.I(FE_OFN47_n10));
   BUFGHD FE_OFC48_n10 (.O(FE_OFN48_n10), 
	.I(n10));
   BUFGHD FE_OFC47_n10 (.O(FE_OFN47_n10), 
	.I(n10));
   BUFGHD FE_OFC46_n9 (.O(FE_OFN46_n9), 
	.I(FE_OFN44_n9));
   BUFGHD FE_OFC45_n9 (.O(FE_OFN45_n9), 
	.I(n9));
   BUFGHD FE_OFC44_n9 (.O(FE_OFN44_n9), 
	.I(n9));
   BUFGHD FE_OFC43_n6 (.O(FE_OFN43_n6), 
	.I(FE_OFN41_n6));
   BUFHHD FE_OFC42_n6 (.O(FE_OFN42_n6), 
	.I(FE_OFN41_n6));
   BUFGHD FE_OFC41_n6 (.O(FE_OFN41_n6), 
	.I(n6));
   BUFGHD FE_OFC40_n6459 (.O(FE_OFN40_n6459), 
	.I(FE_OFN34_n6459));
   BUFGHD FE_OFC39_n6459 (.O(FE_OFN39_n6459), 
	.I(FE_OFN34_n6459));
   BUFHHD FE_OFC38_n6459 (.O(FE_OFN38_n6459), 
	.I(FE_OFN34_n6459));
   BUFGHD FE_OFC37_n6459 (.O(FE_OFN37_n6459), 
	.I(FE_OFN34_n6459));
   BUFHHD FE_OFC36_n6459 (.O(FE_OFN36_n6459), 
	.I(FE_OFN35_n6459));
   BUFHHD FE_OFC35_n6459 (.O(FE_OFN35_n6459), 
	.I(FE_OFN28_n6459));
   BUFHHD FE_OFC34_n6459 (.O(FE_OFN34_n6459), 
	.I(FE_OFN28_n6459));
   BUFHHD FE_OFC33_n6459 (.O(FE_OFN33_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC32_n6459 (.O(FE_OFN32_n6459), 
	.I(FE_OFN26_n6459));
   BUFHHD FE_OFC31_n6459 (.O(FE_OFN31_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC30_n6459 (.O(FE_OFN30_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC29_n6459 (.O(FE_OFN29_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC28_n6459 (.O(FE_OFN28_n6459), 
	.I(FE_OFN26_n6459));
   BUFGHD FE_OFC27_n6459 (.O(FE_OFN27_n6459), 
	.I(FE_OFN26_n6459));
   BUFHHD FE_OFC26_n6459 (.O(FE_OFN26_n6459), 
	.I(FE_OFN25_n6459));
   BUFGHD FE_OFC25_n6459 (.O(FE_OFN25_n6459), 
	.I(n6459));
   BUFHHD FE_OFC24_n6136 (.O(FE_OFN24_n6136), 
	.I(FE_OFN23_n6136));
   BUFHHD FE_OFC23_n6136 (.O(FE_OFN23_n6136), 
	.I(n6136));
   BUFHHD FE_OFC22_n6136 (.O(FE_OFN22_n6136), 
	.I(n6136));
   BUFGHD FE_OFC21_n7440 (.O(FE_OFN21_n7440), 
	.I(FE_OFN9_n7440));
   BUFHHD FE_OFC20_n7440 (.O(FE_OFN20_n7440), 
	.I(FE_OFN9_n7440));
   BUFJHD FE_OFC19_n7440 (.O(FE_OFN19_n7440), 
	.I(FE_OFN14_n7440));
   BUFHHD FE_OFC18_n7440 (.O(FE_OFN18_n7440), 
	.I(FE_OFN9_n7440));
   BUFIHD FE_OFC17_n7440 (.O(FE_OFN17_n7440), 
	.I(n7440));
   BUFIHD FE_OFC16_n7440 (.O(FE_OFN16_n7440), 
	.I(n7440));
   BUFHHD FE_OFC15_n7440 (.O(FE_OFN15_n7440), 
	.I(FE_OFN10_n7440));
   BUFHHD FE_OFC14_n7440 (.O(FE_OFN14_n7440), 
	.I(FE_OFN9_n7440));
   BUFJHD FE_OFC13_n7440 (.O(FE_OFN13_n7440), 
	.I(FE_OFN11_n7440));
   BUFHHD FE_OFC12_n7440 (.O(FE_OFN12_n7440), 
	.I(n7440));
   BUFHHD FE_OFC11_n7440 (.O(FE_OFN11_n7440), 
	.I(FE_OFN7_n7440));
   BUFJHD FE_OFC10_n7440 (.O(FE_OFN10_n7440), 
	.I(n7440));
   BUFGHD FE_OFC9_n7440 (.O(FE_OFN9_n7440), 
	.I(n7440));
   BUFJHD FE_OFC8_n7440 (.O(FE_OFN8_n7440), 
	.I(FE_OFN6_n7440));
   BUFIHD FE_OFC7_n7440 (.O(FE_OFN7_n7440), 
	.I(n7440));
   BUFIHD FE_OFC6_n7440 (.O(FE_OFN6_n7440), 
	.I(n7440));
   BUFHHD FE_OFC5_n7440 (.O(FE_OFN5_n7440), 
	.I(n7440));
   BUFGHD FE_OFC4_n7442 (.O(FE_OFN4_n7442), 
	.I(FE_OFN2_n7442));
   BUFGHD FE_OFC3_n7442 (.O(FE_OFN3_n7442), 
	.I(FE_OFN0_n7442));
   BUFJHD FE_OFC2_n7442 (.O(FE_OFN2_n7442), 
	.I(n7442));
   BUFGHD FE_OFC1_n7442 (.O(FE_OFN1_n7442), 
	.I(n7442));
   BUFGHD FE_OFC0_n7442 (.O(FE_OFN0_n7442), 
	.I(n7442));
   QDFFEHD \ram_reg[253][15]  (.Q(\ram[253][15] ), 
	.D(FE_PHN2407_n4645), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[253][14]  (.Q(\ram[253][14] ), 
	.D(FE_PHN485_n4644), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[253][13]  (.Q(\ram[253][13] ), 
	.D(FE_PHN682_n4643), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[253][12]  (.Q(\ram[253][12] ), 
	.D(FE_PHN3068_n4642), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[253][11]  (.Q(\ram[253][11] ), 
	.D(FE_PHN943_n4641), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[253][10]  (.Q(\ram[253][10] ), 
	.D(FE_PHN2006_n4640), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][9]  (.Q(\ram[253][9] ), 
	.D(FE_PHN655_n4639), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][8]  (.Q(\ram[253][8] ), 
	.D(FE_PHN783_n4638), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][7]  (.Q(\ram[253][7] ), 
	.D(FE_PHN2101_n4637), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[253][6]  (.Q(\ram[253][6] ), 
	.D(FE_PHN220_n4636), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[253][5]  (.Q(\ram[253][5] ), 
	.D(FE_PHN411_n4635), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[253][4]  (.Q(\ram[253][4] ), 
	.D(FE_PHN2779_n4634), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[253][3]  (.Q(\ram[253][3] ), 
	.D(FE_PHN283_n4633), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[253][2]  (.Q(\ram[253][2] ), 
	.D(FE_PHN453_n4632), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[253][1]  (.Q(\ram[253][1] ), 
	.D(FE_PHN2769_n4631), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[253][0]  (.Q(\ram[253][0] ), 
	.D(FE_PHN1560_n4630), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[249][15]  (.Q(\ram[249][15] ), 
	.D(FE_PHN354_n4581), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][14]  (.Q(\ram[249][14] ), 
	.D(FE_PHN368_n4580), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[249][13]  (.Q(\ram[249][13] ), 
	.D(FE_PHN369_n4579), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[249][12]  (.Q(\ram[249][12] ), 
	.D(n4578), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][11]  (.Q(\ram[249][11] ), 
	.D(FE_PHN112_n4577), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][10]  (.Q(\ram[249][10] ), 
	.D(FE_PHN665_n4576), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][9]  (.Q(\ram[249][9] ), 
	.D(FE_PHN2884_n4575), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][8]  (.Q(\ram[249][8] ), 
	.D(FE_PHN474_n4574), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[249][7]  (.Q(\ram[249][7] ), 
	.D(FE_PHN136_n4573), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][6]  (.Q(\ram[249][6] ), 
	.D(FE_PHN878_n4572), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][5]  (.Q(\ram[249][5] ), 
	.D(FE_PHN394_n4571), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][4]  (.Q(\ram[249][4] ), 
	.D(FE_PHN172_n4570), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[249][3]  (.Q(\ram[249][3] ), 
	.D(FE_PHN2545_n4569), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[249][2]  (.Q(\ram[249][2] ), 
	.D(FE_PHN281_n4568), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[249][1]  (.Q(\ram[249][1] ), 
	.D(FE_PHN481_n4567), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[249][0]  (.Q(\ram[249][0] ), 
	.D(FE_PHN412_n4566), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[245][15]  (.Q(\ram[245][15] ), 
	.D(FE_PHN662_n4517), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][14]  (.Q(\ram[245][14] ), 
	.D(FE_PHN884_n4516), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][13]  (.Q(\ram[245][13] ), 
	.D(FE_PHN300_n4515), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][12]  (.Q(\ram[245][12] ), 
	.D(FE_PHN166_n4514), 
	.CK(clk));
   QDFFEHD \ram_reg[245][11]  (.Q(\ram[245][11] ), 
	.D(FE_PHN2316_n4513), 
	.CK(clk));
   QDFFEHD \ram_reg[245][10]  (.Q(\ram[245][10] ), 
	.D(FE_PHN432_n4512), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][9]  (.Q(\ram[245][9] ), 
	.D(FE_PHN1133_n4511), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[245][8]  (.Q(\ram[245][8] ), 
	.D(FE_PHN3031_n4510), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[245][7]  (.Q(\ram[245][7] ), 
	.D(FE_PHN120_n4509), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][6]  (.Q(\ram[245][6] ), 
	.D(FE_PHN437_n4508), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][5]  (.Q(\ram[245][5] ), 
	.D(FE_PHN127_n4507), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][4]  (.Q(\ram[245][4] ), 
	.D(FE_PHN139_n4506), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][3]  (.Q(\ram[245][3] ), 
	.D(FE_PHN1218_n4505), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[245][2]  (.Q(\ram[245][2] ), 
	.D(FE_PHN110_n4504), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[245][1]  (.Q(\ram[245][1] ), 
	.D(FE_PHN440_n4503), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[245][0]  (.Q(\ram[245][0] ), 
	.D(FE_PHN312_n4502), 
	.CK(clk));
   QDFFEHD \ram_reg[241][15]  (.Q(\ram[241][15] ), 
	.D(FE_PHN1395_n4453), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[241][14]  (.Q(\ram[241][14] ), 
	.D(FE_PHN1425_n4452), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][13]  (.Q(\ram[241][13] ), 
	.D(FE_PHN609_n4451), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][12]  (.Q(\ram[241][12] ), 
	.D(FE_PHN961_n4450), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][11]  (.Q(\ram[241][11] ), 
	.D(FE_PHN367_n4449), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][10]  (.Q(\ram[241][10] ), 
	.D(FE_PHN555_n4448), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][9]  (.Q(\ram[241][9] ), 
	.D(FE_PHN1474_n4447), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][8]  (.Q(\ram[241][8] ), 
	.D(FE_PHN118_n4446), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[241][7]  (.Q(\ram[241][7] ), 
	.D(FE_PHN1088_n4445), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][6]  (.Q(\ram[241][6] ), 
	.D(FE_PHN1410_n4444), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][5]  (.Q(\ram[241][5] ), 
	.D(FE_PHN639_n4443), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][4]  (.Q(\ram[241][4] ), 
	.D(FE_PHN1757_n4442), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][3]  (.Q(\ram[241][3] ), 
	.D(FE_PHN507_n4441), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[241][2]  (.Q(\ram[241][2] ), 
	.D(FE_PHN568_n4440), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][1]  (.Q(\ram[241][1] ), 
	.D(n4439), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[241][0]  (.Q(\ram[241][0] ), 
	.D(n4438), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[237][15]  (.Q(\ram[237][15] ), 
	.D(FE_PHN4093_n4389), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][14]  (.Q(\ram[237][14] ), 
	.D(FE_PHN5468_n4388), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][13]  (.Q(\ram[237][13] ), 
	.D(FE_PHN4111_n4387), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][12]  (.Q(\ram[237][12] ), 
	.D(FE_PHN4316_n4386), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][11]  (.Q(\ram[237][11] ), 
	.D(FE_PHN4040_n4385), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][10]  (.Q(\ram[237][10] ), 
	.D(FE_PHN4039_n4384), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][9]  (.Q(\ram[237][9] ), 
	.D(FE_PHN4190_n4383), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][8]  (.Q(\ram[237][8] ), 
	.D(FE_PHN3611_n4382), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][7]  (.Q(\ram[237][7] ), 
	.D(n4381), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][6]  (.Q(\ram[237][6] ), 
	.D(FE_PHN4142_n4380), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][5]  (.Q(\ram[237][5] ), 
	.D(FE_PHN4213_n4379), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[237][4]  (.Q(\ram[237][4] ), 
	.D(FE_PHN4423_n4378), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][3]  (.Q(\ram[237][3] ), 
	.D(FE_PHN4014_n4377), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[237][2]  (.Q(\ram[237][2] ), 
	.D(FE_PHN185_n4376), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[237][1]  (.Q(\ram[237][1] ), 
	.D(FE_PHN4203_n4375), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[237][0]  (.Q(\ram[237][0] ), 
	.D(FE_PHN4328_n4374), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[233][15]  (.Q(\ram[233][15] ), 
	.D(FE_PHN326_n4325), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[233][14]  (.Q(\ram[233][14] ), 
	.D(FE_PHN4024_n4324), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[233][13]  (.Q(\ram[233][13] ), 
	.D(FE_PHN4070_n4323), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[233][12]  (.Q(\ram[233][12] ), 
	.D(FE_PHN1056_n4322), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[233][11]  (.Q(\ram[233][11] ), 
	.D(FE_PHN2148_n4321), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[233][10]  (.Q(\ram[233][10] ), 
	.D(FE_PHN186_n4320), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][9]  (.Q(\ram[233][9] ), 
	.D(FE_PHN493_n4319), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][8]  (.Q(\ram[233][8] ), 
	.D(FE_PHN337_n4318), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][7]  (.Q(\ram[233][7] ), 
	.D(FE_PHN237_n4317), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[233][6]  (.Q(\ram[233][6] ), 
	.D(FE_PHN4576_n4316), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][5]  (.Q(\ram[233][5] ), 
	.D(FE_PHN197_n4315), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[233][4]  (.Q(\ram[233][4] ), 
	.D(FE_PHN2186_n4314), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][3]  (.Q(\ram[233][3] ), 
	.D(FE_PHN140_n4313), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[233][2]  (.Q(\ram[233][2] ), 
	.D(FE_PHN2321_n4312), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[233][1]  (.Q(\ram[233][1] ), 
	.D(FE_PHN4683_n4311), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[233][0]  (.Q(\ram[233][0] ), 
	.D(FE_PHN317_n4310), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[229][15]  (.Q(\ram[229][15] ), 
	.D(FE_PHN5585_n4261), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][14]  (.Q(\ram[229][14] ), 
	.D(FE_PHN4275_n4260), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[229][13]  (.Q(\ram[229][13] ), 
	.D(FE_PHN4572_n4259), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[229][12]  (.Q(\ram[229][12] ), 
	.D(n4258), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[229][11]  (.Q(\ram[229][11] ), 
	.D(FE_PHN345_n4257), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][10]  (.Q(\ram[229][10] ), 
	.D(FE_PHN320_n4256), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][9]  (.Q(\ram[229][9] ), 
	.D(FE_PHN5222_n4255), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[229][8]  (.Q(\ram[229][8] ), 
	.D(FE_PHN4156_n4254), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][7]  (.Q(\ram[229][7] ), 
	.D(FE_PHN868_n4253), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[229][6]  (.Q(\ram[229][6] ), 
	.D(FE_PHN4631_n4252), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[229][5]  (.Q(\ram[229][5] ), 
	.D(FE_PHN5373_n4251), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[229][4]  (.Q(\ram[229][4] ), 
	.D(FE_PHN1103_n4250), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[229][3]  (.Q(\ram[229][3] ), 
	.D(n4249), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[229][2]  (.Q(\ram[229][2] ), 
	.D(FE_PHN4325_n4248), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[229][1]  (.Q(\ram[229][1] ), 
	.D(FE_PHN240_n4247), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[229][0]  (.Q(\ram[229][0] ), 
	.D(FE_PHN374_n4246), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[225][15]  (.Q(\ram[225][15] ), 
	.D(FE_PHN1052_n4197), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[225][14]  (.Q(\ram[225][14] ), 
	.D(FE_PHN4122_n4196), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][13]  (.Q(\ram[225][13] ), 
	.D(FE_PHN4012_n4195), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[225][12]  (.Q(\ram[225][12] ), 
	.D(FE_PHN4427_n4194), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][11]  (.Q(\ram[225][11] ), 
	.D(FE_PHN366_n4193), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[225][10]  (.Q(\ram[225][10] ), 
	.D(FE_PHN1762_n4192), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[225][9]  (.Q(\ram[225][9] ), 
	.D(FE_PHN234_n4191), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[225][8]  (.Q(\ram[225][8] ), 
	.D(FE_PHN171_n4190), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[225][7]  (.Q(\ram[225][7] ), 
	.D(FE_PHN1852_n4189), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[225][6]  (.Q(\ram[225][6] ), 
	.D(FE_PHN4477_n4188), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][5]  (.Q(\ram[225][5] ), 
	.D(FE_PHN3918_n4187), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[225][4]  (.Q(\ram[225][4] ), 
	.D(FE_PHN288_n4186), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[225][3]  (.Q(\ram[225][3] ), 
	.D(FE_PHN4431_n4185), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][2]  (.Q(\ram[225][2] ), 
	.D(FE_PHN1760_n4184), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[225][1]  (.Q(\ram[225][1] ), 
	.D(FE_PHN5445_n4183), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[225][0]  (.Q(\ram[225][0] ), 
	.D(FE_PHN190_n4182), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[221][15]  (.Q(\ram[221][15] ), 
	.D(FE_PHN1122_n4133), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][14]  (.Q(\ram[221][14] ), 
	.D(FE_PHN210_n4132), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][13]  (.Q(\ram[221][13] ), 
	.D(FE_PHN1923_n4131), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][12]  (.Q(\ram[221][12] ), 
	.D(FE_PHN557_n4130), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][11]  (.Q(\ram[221][11] ), 
	.D(FE_PHN456_n4129), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][10]  (.Q(\ram[221][10] ), 
	.D(FE_PHN2452_n4128), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[221][9]  (.Q(\ram[221][9] ), 
	.D(FE_PHN1258_n4127), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][8]  (.Q(\ram[221][8] ), 
	.D(FE_PHN1551_n4126), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][7]  (.Q(\ram[221][7] ), 
	.D(FE_PHN469_n4125), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[221][6]  (.Q(\ram[221][6] ), 
	.D(FE_PHN1099_n4124), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[221][5]  (.Q(\ram[221][5] ), 
	.D(FE_PHN3270_n4123), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][4]  (.Q(\ram[221][4] ), 
	.D(FE_PHN1767_n4122), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[221][3]  (.Q(\ram[221][3] ), 
	.D(FE_PHN6648_n4121), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[221][2]  (.Q(\ram[221][2] ), 
	.D(FE_PHN295_n4120), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[221][1]  (.Q(\ram[221][1] ), 
	.D(n4119), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[221][0]  (.Q(\ram[221][0] ), 
	.D(FE_PHN534_n4118), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[217][15]  (.Q(\ram[217][15] ), 
	.D(FE_PHN1677_n4069), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][14]  (.Q(\ram[217][14] ), 
	.D(FE_PHN130_n4068), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][13]  (.Q(\ram[217][13] ), 
	.D(FE_PHN1021_n4067), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][12]  (.Q(\ram[217][12] ), 
	.D(FE_PHN777_n4066), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][11]  (.Q(\ram[217][11] ), 
	.D(FE_PHN302_n4065), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[217][10]  (.Q(\ram[217][10] ), 
	.D(FE_PHN135_n4064), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][9]  (.Q(\ram[217][9] ), 
	.D(FE_PHN976_n4063), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][8]  (.Q(\ram[217][8] ), 
	.D(FE_PHN5675_n4062), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[217][7]  (.Q(\ram[217][7] ), 
	.D(FE_PHN1241_n4061), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][6]  (.Q(\ram[217][6] ), 
	.D(FE_PHN1509_n4060), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][5]  (.Q(\ram[217][5] ), 
	.D(FE_PHN1770_n4059), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[217][4]  (.Q(\ram[217][4] ), 
	.D(FE_PHN847_n4058), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[217][3]  (.Q(\ram[217][3] ), 
	.D(n4057), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[217][2]  (.Q(\ram[217][2] ), 
	.D(FE_PHN695_n4056), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[217][1]  (.Q(\ram[217][1] ), 
	.D(FE_PHN155_n4055), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[217][0]  (.Q(\ram[217][0] ), 
	.D(FE_PHN431_n4054), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[213][15]  (.Q(\ram[213][15] ), 
	.D(FE_PHN4064_n4005), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[213][14]  (.Q(\ram[213][14] ), 
	.D(FE_PHN173_n4004), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][13]  (.Q(\ram[213][13] ), 
	.D(FE_PHN4071_n4003), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[213][12]  (.Q(\ram[213][12] ), 
	.D(FE_PHN6684_n4002), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[213][11]  (.Q(\ram[213][11] ), 
	.D(FE_PHN4191_n4001), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][10]  (.Q(\ram[213][10] ), 
	.D(FE_PHN4993_n4000), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][9]  (.Q(\ram[213][9] ), 
	.D(FE_PHN4044_n3999), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[213][8]  (.Q(\ram[213][8] ), 
	.D(FE_PHN5226_n3998), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[213][7]  (.Q(\ram[213][7] ), 
	.D(FE_PHN215_n3997), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][6]  (.Q(\ram[213][6] ), 
	.D(FE_PHN5269_n3996), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][5]  (.Q(\ram[213][5] ), 
	.D(FE_PHN121_n3995), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[213][4]  (.Q(\ram[213][4] ), 
	.D(FE_PHN4384_n3994), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][3]  (.Q(\ram[213][3] ), 
	.D(FE_PHN5392_n3993), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[213][2]  (.Q(\ram[213][2] ), 
	.D(FE_PHN4378_n3992), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[213][1]  (.Q(\ram[213][1] ), 
	.D(FE_PHN231_n3991), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[213][0]  (.Q(\ram[213][0] ), 
	.D(FE_PHN201_n3990), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[209][15]  (.Q(\ram[209][15] ), 
	.D(FE_PHN708_n3941), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[209][14]  (.Q(\ram[209][14] ), 
	.D(FE_PHN4724_n3940), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[209][13]  (.Q(\ram[209][13] ), 
	.D(FE_PHN4072_n3939), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][12]  (.Q(\ram[209][12] ), 
	.D(FE_PHN209_n3938), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][11]  (.Q(\ram[209][11] ), 
	.D(FE_PHN4034_n3937), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][10]  (.Q(\ram[209][10] ), 
	.D(FE_PHN4737_n3936), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][9]  (.Q(\ram[209][9] ), 
	.D(FE_PHN289_n3935), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][8]  (.Q(\ram[209][8] ), 
	.D(FE_PHN3291_n3934), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][7]  (.Q(\ram[209][7] ), 
	.D(FE_PHN1476_n3933), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[209][6]  (.Q(\ram[209][6] ), 
	.D(FE_PHN3774_n3932), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[209][5]  (.Q(\ram[209][5] ), 
	.D(FE_PHN4025_n3931), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[209][4]  (.Q(\ram[209][4] ), 
	.D(FE_PHN4043_n3930), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[209][3]  (.Q(\ram[209][3] ), 
	.D(FE_PHN4281_n3929), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[209][2]  (.Q(\ram[209][2] ), 
	.D(FE_PHN472_n3928), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[209][1]  (.Q(\ram[209][1] ), 
	.D(FE_PHN3341_n3927), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[209][0]  (.Q(\ram[209][0] ), 
	.D(FE_PHN4017_n3926), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[205][15]  (.Q(\ram[205][15] ), 
	.D(FE_PHN458_n3877), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][14]  (.Q(\ram[205][14] ), 
	.D(FE_PHN1491_n3876), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][13]  (.Q(\ram[205][13] ), 
	.D(FE_PHN701_n3875), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[205][12]  (.Q(\ram[205][12] ), 
	.D(FE_PHN1121_n3874), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][11]  (.Q(\ram[205][11] ), 
	.D(FE_PHN1175_n3873), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][10]  (.Q(\ram[205][10] ), 
	.D(FE_PHN2126_n3872), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][9]  (.Q(\ram[205][9] ), 
	.D(FE_PHN810_n3871), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][8]  (.Q(\ram[205][8] ), 
	.D(FE_PHN131_n3870), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[205][7]  (.Q(\ram[205][7] ), 
	.D(FE_PHN1828_n3869), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][6]  (.Q(\ram[205][6] ), 
	.D(FE_PHN570_n3868), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][5]  (.Q(\ram[205][5] ), 
	.D(FE_PHN1517_n3867), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][4]  (.Q(\ram[205][4] ), 
	.D(FE_PHN126_n3866), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][3]  (.Q(\ram[205][3] ), 
	.D(FE_PHN988_n3865), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][2]  (.Q(\ram[205][2] ), 
	.D(FE_PHN142_n3864), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[205][1]  (.Q(\ram[205][1] ), 
	.D(FE_PHN236_n3863), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[205][0]  (.Q(\ram[205][0] ), 
	.D(FE_PHN466_n3862), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[201][15]  (.Q(\ram[201][15] ), 
	.D(FE_PHN1157_n3813), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][14]  (.Q(\ram[201][14] ), 
	.D(FE_PHN2294_n3812), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][13]  (.Q(\ram[201][13] ), 
	.D(FE_PHN1333_n3811), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[201][12]  (.Q(\ram[201][12] ), 
	.D(FE_PHN445_n3810), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][11]  (.Q(\ram[201][11] ), 
	.D(FE_PHN1366_n3809), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][10]  (.Q(\ram[201][10] ), 
	.D(FE_PHN1147_n3808), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][9]  (.Q(\ram[201][9] ), 
	.D(FE_PHN114_n3807), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[201][8]  (.Q(\ram[201][8] ), 
	.D(FE_PHN1237_n3806), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[201][7]  (.Q(\ram[201][7] ), 
	.D(FE_PHN350_n3805), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][6]  (.Q(\ram[201][6] ), 
	.D(FE_PHN906_n3804), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[201][5]  (.Q(\ram[201][5] ), 
	.D(n3803), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[201][4]  (.Q(\ram[201][4] ), 
	.D(FE_PHN1151_n3802), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[201][3]  (.Q(\ram[201][3] ), 
	.D(FE_PHN1415_n3801), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[201][2]  (.Q(\ram[201][2] ), 
	.D(FE_PHN577_n3800), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][1]  (.Q(\ram[201][1] ), 
	.D(FE_PHN2154_n3799), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[201][0]  (.Q(\ram[201][0] ), 
	.D(FE_PHN451_n3798), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[197][15]  (.Q(\ram[197][15] ), 
	.D(FE_PHN381_n3749), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][14]  (.Q(\ram[197][14] ), 
	.D(FE_PHN324_n3748), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][13]  (.Q(\ram[197][13] ), 
	.D(FE_PHN248_n3747), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[197][12]  (.Q(\ram[197][12] ), 
	.D(FE_PHN548_n3746), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[197][11]  (.Q(\ram[197][11] ), 
	.D(FE_PHN869_n3745), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][10]  (.Q(\ram[197][10] ), 
	.D(FE_PHN208_n3744), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][9]  (.Q(\ram[197][9] ), 
	.D(FE_PHN341_n3743), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[197][8]  (.Q(\ram[197][8] ), 
	.D(FE_PHN530_n3742), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][7]  (.Q(\ram[197][7] ), 
	.D(FE_PHN1413_n3741), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][6]  (.Q(\ram[197][6] ), 
	.D(FE_PHN1013_n3740), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][5]  (.Q(\ram[197][5] ), 
	.D(FE_PHN115_n3739), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][4]  (.Q(\ram[197][4] ), 
	.D(FE_PHN2713_n3738), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][3]  (.Q(\ram[197][3] ), 
	.D(FE_PHN909_n3737), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[197][2]  (.Q(\ram[197][2] ), 
	.D(FE_PHN2033_n3736), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[197][1]  (.Q(\ram[197][1] ), 
	.D(FE_PHN224_n3735), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[197][0]  (.Q(\ram[197][0] ), 
	.D(FE_PHN174_n3734), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[193][15]  (.Q(\ram[193][15] ), 
	.D(FE_PHN904_n3685), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][14]  (.Q(\ram[193][14] ), 
	.D(FE_PHN1464_n3684), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][13]  (.Q(\ram[193][13] ), 
	.D(FE_PHN2404_n3683), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[193][12]  (.Q(\ram[193][12] ), 
	.D(FE_PHN191_n3682), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][11]  (.Q(\ram[193][11] ), 
	.D(FE_PHN1017_n3681), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][10]  (.Q(\ram[193][10] ), 
	.D(FE_PHN607_n3680), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[193][9]  (.Q(\ram[193][9] ), 
	.D(FE_PHN405_n3679), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][8]  (.Q(\ram[193][8] ), 
	.D(FE_PHN328_n3678), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[193][7]  (.Q(\ram[193][7] ), 
	.D(FE_PHN383_n3677), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[193][6]  (.Q(\ram[193][6] ), 
	.D(FE_PHN503_n3676), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][5]  (.Q(\ram[193][5] ), 
	.D(FE_PHN838_n3675), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][4]  (.Q(\ram[193][4] ), 
	.D(FE_PHN2916_n3674), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][3]  (.Q(\ram[193][3] ), 
	.D(FE_PHN207_n3673), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[193][2]  (.Q(\ram[193][2] ), 
	.D(FE_PHN1487_n3672), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[193][1]  (.Q(\ram[193][1] ), 
	.D(FE_PHN1984_n3671), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[193][0]  (.Q(\ram[193][0] ), 
	.D(FE_PHN407_n3670), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[189][15]  (.Q(\ram[189][15] ), 
	.D(FE_PHN149_n3621), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][14]  (.Q(\ram[189][14] ), 
	.D(FE_PHN1672_n3620), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[189][13]  (.Q(\ram[189][13] ), 
	.D(FE_PHN106_n3619), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[189][12]  (.Q(\ram[189][12] ), 
	.D(FE_PHN160_n3618), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[189][11]  (.Q(\ram[189][11] ), 
	.D(FE_PHN2631_n3617), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[189][10]  (.Q(\ram[189][10] ), 
	.D(FE_PHN2917_n3616), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[189][9]  (.Q(\ram[189][9] ), 
	.D(FE_PHN1216_n3615), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[189][8]  (.Q(\ram[189][8] ), 
	.D(FE_PHN2438_n3614), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][7]  (.Q(\ram[189][7] ), 
	.D(FE_PHN1665_n3613), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][6]  (.Q(\ram[189][6] ), 
	.D(FE_PHN1782_n3612), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[189][5]  (.Q(\ram[189][5] ), 
	.D(FE_PHN266_n3611), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[189][4]  (.Q(\ram[189][4] ), 
	.D(FE_PHN218_n3610), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][3]  (.Q(\ram[189][3] ), 
	.D(FE_PHN146_n3609), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[189][2]  (.Q(\ram[189][2] ), 
	.D(FE_PHN353_n3608), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[189][1]  (.Q(\ram[189][1] ), 
	.D(FE_PHN1346_n3607), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[189][0]  (.Q(\ram[189][0] ), 
	.D(FE_PHN134_n3606), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[185][15]  (.Q(\ram[185][15] ), 
	.D(FE_PHN282_n3557), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][14]  (.Q(\ram[185][14] ), 
	.D(FE_PHN147_n3556), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][13]  (.Q(\ram[185][13] ), 
	.D(FE_PHN487_n3555), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][12]  (.Q(\ram[185][12] ), 
	.D(FE_PHN102_n3554), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[185][11]  (.Q(\ram[185][11] ), 
	.D(FE_PHN989_n3553), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][10]  (.Q(\ram[185][10] ), 
	.D(FE_PHN105_n3552), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[185][9]  (.Q(\ram[185][9] ), 
	.D(FE_PHN841_n3551), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[185][8]  (.Q(\ram[185][8] ), 
	.D(FE_PHN153_n3550), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][7]  (.Q(\ram[185][7] ), 
	.D(FE_PHN109_n3549), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][6]  (.Q(\ram[185][6] ), 
	.D(FE_PHN161_n3548), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][5]  (.Q(\ram[185][5] ), 
	.D(FE_PHN101_n3547), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][4]  (.Q(\ram[185][4] ), 
	.D(FE_PHN125_n3546), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[185][3]  (.Q(\ram[185][3] ), 
	.D(FE_PHN104_n3545), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[185][2]  (.Q(\ram[185][2] ), 
	.D(FE_PHN276_n3544), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][1]  (.Q(\ram[185][1] ), 
	.D(FE_PHN230_n3543), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[185][0]  (.Q(\ram[185][0] ), 
	.D(FE_PHN100_n3542), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[181][15]  (.Q(\ram[181][15] ), 
	.D(FE_PHN193_n3493), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[181][14]  (.Q(\ram[181][14] ), 
	.D(FE_PHN1363_n3492), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[181][13]  (.Q(\ram[181][13] ), 
	.D(FE_PHN183_n3491), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[181][12]  (.Q(\ram[181][12] ), 
	.D(FE_PHN333_n3490), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[181][11]  (.Q(\ram[181][11] ), 
	.D(FE_PHN323_n3489), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[181][10]  (.Q(\ram[181][10] ), 
	.D(FE_PHN1314_n3488), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][9]  (.Q(\ram[181][9] ), 
	.D(FE_PHN3056_n3487), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][8]  (.Q(\ram[181][8] ), 
	.D(FE_PHN860_n3486), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][7]  (.Q(\ram[181][7] ), 
	.D(FE_PHN814_n3485), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[181][6]  (.Q(\ram[181][6] ), 
	.D(FE_PHN325_n3484), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[181][5]  (.Q(\ram[181][5] ), 
	.D(FE_PHN3169_n3483), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[181][4]  (.Q(\ram[181][4] ), 
	.D(FE_PHN1504_n3482), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[181][3]  (.Q(\ram[181][3] ), 
	.D(FE_PHN3186_n3481), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[181][2]  (.Q(\ram[181][2] ), 
	.D(FE_PHN1298_n3480), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[181][1]  (.Q(\ram[181][1] ), 
	.D(FE_PHN759_n3479), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[181][0]  (.Q(\ram[181][0] ), 
	.D(FE_PHN2761_n3478), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[177][15]  (.Q(\ram[177][15] ), 
	.D(FE_PHN2687_n3429), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[177][14]  (.Q(\ram[177][14] ), 
	.D(FE_PHN1785_n3428), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][13]  (.Q(\ram[177][13] ), 
	.D(FE_PHN3217_n3427), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[177][12]  (.Q(\ram[177][12] ), 
	.D(FE_PHN2869_n3426), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[177][11]  (.Q(\ram[177][11] ), 
	.D(FE_PHN1515_n3425), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[177][10]  (.Q(\ram[177][10] ), 
	.D(FE_PHN1557_n3424), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[177][9]  (.Q(\ram[177][9] ), 
	.D(FE_PHN815_n3423), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][8]  (.Q(\ram[177][8] ), 
	.D(FE_PHN2550_n3422), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[177][7]  (.Q(\ram[177][7] ), 
	.D(FE_PHN782_n3421), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][6]  (.Q(\ram[177][6] ), 
	.D(FE_PHN1985_n3420), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[177][5]  (.Q(\ram[177][5] ), 
	.D(FE_PHN1654_n3419), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[177][4]  (.Q(\ram[177][4] ), 
	.D(FE_PHN825_n3418), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][3]  (.Q(\ram[177][3] ), 
	.D(FE_PHN2392_n3417), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[177][2]  (.Q(\ram[177][2] ), 
	.D(FE_PHN1971_n3416), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][1]  (.Q(\ram[177][1] ), 
	.D(FE_PHN1406_n3415), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[177][0]  (.Q(\ram[177][0] ), 
	.D(FE_PHN1421_n3414), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[173][15]  (.Q(\ram[173][15] ), 
	.D(FE_PHN154_n3365), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][14]  (.Q(\ram[173][14] ), 
	.D(FE_PHN517_n3364), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][13]  (.Q(\ram[173][13] ), 
	.D(FE_PHN2700_n3363), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[173][12]  (.Q(\ram[173][12] ), 
	.D(FE_PHN450_n3362), 
	.CK(clk));
   QDFFEHD \ram_reg[173][11]  (.Q(\ram[173][11] ), 
	.D(FE_PHN1706_n3361), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[173][10]  (.Q(\ram[173][10] ), 
	.D(FE_PHN894_n3360), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[173][9]  (.Q(\ram[173][9] ), 
	.D(FE_PHN1768_n3359), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][8]  (.Q(\ram[173][8] ), 
	.D(FE_PHN553_n3358), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[173][7]  (.Q(\ram[173][7] ), 
	.D(FE_PHN2094_n3357), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][6]  (.Q(\ram[173][6] ), 
	.D(FE_PHN730_n3356), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][5]  (.Q(\ram[173][5] ), 
	.D(FE_PHN329_n3355), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][4]  (.Q(\ram[173][4] ), 
	.D(FE_PHN355_n3354), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][3]  (.Q(\ram[173][3] ), 
	.D(FE_PHN178_n3353), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[173][2]  (.Q(\ram[173][2] ), 
	.D(FE_PHN205_n3352), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][1]  (.Q(\ram[173][1] ), 
	.D(FE_PHN2347_n3351), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[173][0]  (.Q(\ram[173][0] ), 
	.D(FE_PHN262_n3350), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[169][15]  (.Q(\ram[169][15] ), 
	.D(FE_PHN117_n3301), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][14]  (.Q(\ram[169][14] ), 
	.D(FE_PHN177_n3300), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][13]  (.Q(\ram[169][13] ), 
	.D(FE_PHN1176_n3299), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][12]  (.Q(\ram[169][12] ), 
	.D(FE_PHN2323_n3298), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][11]  (.Q(\ram[169][11] ), 
	.D(FE_PHN657_n3297), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][10]  (.Q(\ram[169][10] ), 
	.D(FE_PHN842_n3296), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][9]  (.Q(\ram[169][9] ), 
	.D(FE_PHN514_n3295), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][8]  (.Q(\ram[169][8] ), 
	.D(FE_PHN1594_n3294), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[169][7]  (.Q(\ram[169][7] ), 
	.D(FE_PHN1802_n3293), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][6]  (.Q(\ram[169][6] ), 
	.D(FE_PHN181_n3292), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][5]  (.Q(\ram[169][5] ), 
	.D(FE_PHN1210_n3291), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][4]  (.Q(\ram[169][4] ), 
	.D(FE_PHN1909_n3290), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][3]  (.Q(\ram[169][3] ), 
	.D(FE_PHN944_n3289), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[169][2]  (.Q(\ram[169][2] ), 
	.D(FE_PHN844_n3288), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[169][1]  (.Q(\ram[169][1] ), 
	.D(FE_PHN1657_n3287), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[169][0]  (.Q(\ram[169][0] ), 
	.D(FE_PHN157_n3286), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[165][15]  (.Q(\ram[165][15] ), 
	.D(FE_PHN2227_n3237), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[165][14]  (.Q(\ram[165][14] ), 
	.D(FE_PHN364_n3236), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[165][13]  (.Q(\ram[165][13] ), 
	.D(FE_PHN2568_n3235), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[165][12]  (.Q(\ram[165][12] ), 
	.D(FE_PHN162_n3234), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[165][11]  (.Q(\ram[165][11] ), 
	.D(FE_PHN342_n3233), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][10]  (.Q(\ram[165][10] ), 
	.D(FE_PHN1702_n3232), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][9]  (.Q(\ram[165][9] ), 
	.D(FE_PHN254_n3231), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][8]  (.Q(\ram[165][8] ), 
	.D(FE_PHN6698_n3230), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][7]  (.Q(\ram[165][7] ), 
	.D(FE_PHN1603_n3229), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][6]  (.Q(\ram[165][6] ), 
	.D(FE_PHN1108_n3228), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][5]  (.Q(\ram[165][5] ), 
	.D(FE_PHN1231_n3227), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][4]  (.Q(\ram[165][4] ), 
	.D(FE_PHN122_n3226), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[165][3]  (.Q(\ram[165][3] ), 
	.D(FE_PHN1914_n3225), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][2]  (.Q(\ram[165][2] ), 
	.D(FE_PHN159_n3224), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[165][1]  (.Q(\ram[165][1] ), 
	.D(FE_PHN4243_n3223), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[165][0]  (.Q(\ram[165][0] ), 
	.D(FE_PHN828_n3222), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[161][15]  (.Q(\ram[161][15] ), 
	.D(FE_PHN1536_n3173), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][14]  (.Q(\ram[161][14] ), 
	.D(FE_PHN246_n3172), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][13]  (.Q(\ram[161][13] ), 
	.D(FE_PHN726_n3171), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][12]  (.Q(\ram[161][12] ), 
	.D(FE_PHN213_n3170), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[161][11]  (.Q(\ram[161][11] ), 
	.D(FE_PHN521_n3169), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[161][10]  (.Q(\ram[161][10] ), 
	.D(FE_PHN805_n3168), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[161][9]  (.Q(\ram[161][9] ), 
	.D(FE_PHN175_n3167), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[161][8]  (.Q(\ram[161][8] ), 
	.D(FE_PHN390_n3166), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[161][7]  (.Q(\ram[161][7] ), 
	.D(FE_PHN343_n3165), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][6]  (.Q(\ram[161][6] ), 
	.D(FE_PHN164_n3164), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][5]  (.Q(\ram[161][5] ), 
	.D(FE_PHN1458_n3163), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[161][4]  (.Q(\ram[161][4] ), 
	.D(FE_PHN1284_n3162), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][3]  (.Q(\ram[161][3] ), 
	.D(FE_PHN1198_n3161), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][2]  (.Q(\ram[161][2] ), 
	.D(FE_PHN1806_n3160), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[161][1]  (.Q(\ram[161][1] ), 
	.D(FE_PHN925_n3159), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[161][0]  (.Q(\ram[161][0] ), 
	.D(FE_PHN2046_n3158), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[157][15]  (.Q(\ram[157][15] ), 
	.D(FE_PHN4678_n3109), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[157][14]  (.Q(\ram[157][14] ), 
	.D(FE_PHN4068_n3108), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][13]  (.Q(\ram[157][13] ), 
	.D(FE_PHN4077_n3107), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][12]  (.Q(\ram[157][12] ), 
	.D(FE_PHN132_n3106), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][11]  (.Q(\ram[157][11] ), 
	.D(FE_PHN4080_n3105), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][10]  (.Q(\ram[157][10] ), 
	.D(FE_PHN3351_n3104), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[157][9]  (.Q(\ram[157][9] ), 
	.D(FE_PHN4170_n3103), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[157][8]  (.Q(\ram[157][8] ), 
	.D(FE_PHN5475_n3102), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[157][7]  (.Q(\ram[157][7] ), 
	.D(FE_PHN199_n3101), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[157][6]  (.Q(\ram[157][6] ), 
	.D(FE_PHN5544_n3100), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[157][5]  (.Q(\ram[157][5] ), 
	.D(FE_PHN5522_n3099), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[157][4]  (.Q(\ram[157][4] ), 
	.D(FE_PHN4641_n3098), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[157][3]  (.Q(\ram[157][3] ), 
	.D(FE_PHN278_n3097), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[157][2]  (.Q(\ram[157][2] ), 
	.D(FE_PHN5482_n3096), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[157][1]  (.Q(\ram[157][1] ), 
	.D(FE_PHN4244_n3095), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[157][0]  (.Q(\ram[157][0] ), 
	.D(FE_PHN4018_n3094), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[153][15]  (.Q(\ram[153][15] ), 
	.D(FE_PHN1102_n3045), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[153][14]  (.Q(\ram[153][14] ), 
	.D(FE_PHN4656_n3044), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][13]  (.Q(\ram[153][13] ), 
	.D(FE_PHN3310_n3043), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][12]  (.Q(\ram[153][12] ), 
	.D(FE_PHN4260_n3042), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[153][11]  (.Q(\ram[153][11] ), 
	.D(n3041), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][10]  (.Q(\ram[153][10] ), 
	.D(FE_PHN3746_n3040), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[153][9]  (.Q(\ram[153][9] ), 
	.D(FE_PHN1085_n3039), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[153][8]  (.Q(\ram[153][8] ), 
	.D(FE_PHN4717_n3038), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[153][7]  (.Q(\ram[153][7] ), 
	.D(n3037), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][6]  (.Q(\ram[153][6] ), 
	.D(FE_PHN4475_n3036), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[153][5]  (.Q(\ram[153][5] ), 
	.D(FE_PHN5491_n3035), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[153][4]  (.Q(\ram[153][4] ), 
	.D(FE_PHN5713_n3034), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[153][3]  (.Q(\ram[153][3] ), 
	.D(FE_PHN4817_n3033), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][2]  (.Q(\ram[153][2] ), 
	.D(FE_PHN5497_n3032), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][1]  (.Q(\ram[153][1] ), 
	.D(FE_PHN4258_n3031), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[153][0]  (.Q(\ram[153][0] ), 
	.D(FE_PHN4294_n3030), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[149][15]  (.Q(\ram[149][15] ), 
	.D(FE_PHN4050_n2981), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][14]  (.Q(\ram[149][14] ), 
	.D(FE_PHN5275_n2980), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][13]  (.Q(\ram[149][13] ), 
	.D(FE_PHN4063_n2979), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][12]  (.Q(\ram[149][12] ), 
	.D(FE_PHN4047_n2978), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][11]  (.Q(\ram[149][11] ), 
	.D(FE_PHN4057_n2977), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[149][10]  (.Q(\ram[149][10] ), 
	.D(FE_PHN4030_n2976), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[149][9]  (.Q(\ram[149][9] ), 
	.D(FE_PHN4424_n2975), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[149][8]  (.Q(\ram[149][8] ), 
	.D(FE_PHN4728_n2974), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[149][7]  (.Q(\ram[149][7] ), 
	.D(FE_PHN4081_n2973), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][6]  (.Q(\ram[149][6] ), 
	.D(FE_PHN3445_n2972), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][5]  (.Q(\ram[149][5] ), 
	.D(FE_PHN4539_n2971), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][4]  (.Q(\ram[149][4] ), 
	.D(FE_PHN4675_n2970), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][3]  (.Q(\ram[149][3] ), 
	.D(FE_PHN4245_n2969), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][2]  (.Q(\ram[149][2] ), 
	.D(FE_PHN4284_n2968), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[149][1]  (.Q(\ram[149][1] ), 
	.D(FE_PHN4297_n2967), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[149][0]  (.Q(\ram[149][0] ), 
	.D(FE_PHN4019_n2966), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[145][15]  (.Q(\ram[145][15] ), 
	.D(FE_PHN1055_n2917), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[145][14]  (.Q(\ram[145][14] ), 
	.D(FE_PHN4666_n2916), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][13]  (.Q(\ram[145][13] ), 
	.D(FE_PHN497_n2915), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[145][12]  (.Q(\ram[145][12] ), 
	.D(FE_PHN673_n2914), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][11]  (.Q(\ram[145][11] ), 
	.D(FE_PHN1816_n2913), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[145][10]  (.Q(\ram[145][10] ), 
	.D(n2912), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[145][9]  (.Q(\ram[145][9] ), 
	.D(FE_PHN698_n2911), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][8]  (.Q(\ram[145][8] ), 
	.D(FE_PHN4747_n2910), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[145][7]  (.Q(\ram[145][7] ), 
	.D(n2909), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][6]  (.Q(\ram[145][6] ), 
	.D(FE_PHN5756_n2908), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][5]  (.Q(\ram[145][5] ), 
	.D(FE_PHN5741_n2907), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][4]  (.Q(\ram[145][4] ), 
	.D(FE_PHN3482_n2906), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][3]  (.Q(\ram[145][3] ), 
	.D(FE_PHN697_n2905), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][2]  (.Q(\ram[145][2] ), 
	.D(FE_PHN3404_n2904), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[145][1]  (.Q(\ram[145][1] ), 
	.D(n2903), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[145][0]  (.Q(\ram[145][0] ), 
	.D(n2902), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[141][15]  (.Q(\ram[141][15] ), 
	.D(FE_PHN1299_n2853), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[141][14]  (.Q(\ram[141][14] ), 
	.D(FE_PHN642_n2852), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][13]  (.Q(\ram[141][13] ), 
	.D(FE_PHN1015_n2851), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][12]  (.Q(\ram[141][12] ), 
	.D(FE_PHN613_n2850), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[141][11]  (.Q(\ram[141][11] ), 
	.D(FE_PHN892_n2849), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[141][10]  (.Q(\ram[141][10] ), 
	.D(FE_PHN940_n2848), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[141][9]  (.Q(\ram[141][9] ), 
	.D(FE_PHN1833_n2847), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][8]  (.Q(\ram[141][8] ), 
	.D(FE_PHN997_n2846), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[141][7]  (.Q(\ram[141][7] ), 
	.D(FE_PHN3015_n2845), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][6]  (.Q(\ram[141][6] ), 
	.D(FE_PHN1402_n2844), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[141][5]  (.Q(\ram[141][5] ), 
	.D(FE_PHN2079_n2843), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[141][4]  (.Q(\ram[141][4] ), 
	.D(FE_PHN2360_n2842), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][3]  (.Q(\ram[141][3] ), 
	.D(FE_PHN384_n2841), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[141][2]  (.Q(\ram[141][2] ), 
	.D(FE_PHN1502_n2840), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][1]  (.Q(\ram[141][1] ), 
	.D(FE_PHN535_n2839), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[141][0]  (.Q(\ram[141][0] ), 
	.D(FE_PHN1219_n2838), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[137][15]  (.Q(\ram[137][15] ), 
	.D(FE_PHN473_n2789), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][14]  (.Q(\ram[137][14] ), 
	.D(FE_PHN3110_n2788), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][13]  (.Q(\ram[137][13] ), 
	.D(FE_PHN344_n2787), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[137][12]  (.Q(\ram[137][12] ), 
	.D(FE_PHN554_n2786), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][11]  (.Q(\ram[137][11] ), 
	.D(FE_PHN1080_n2785), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[137][10]  (.Q(\ram[137][10] ), 
	.D(FE_PHN1404_n2784), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[137][9]  (.Q(\ram[137][9] ), 
	.D(FE_PHN747_n2783), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[137][8]  (.Q(\ram[137][8] ), 
	.D(FE_PHN2043_n2782), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[137][7]  (.Q(\ram[137][7] ), 
	.D(FE_PHN795_n2781), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][6]  (.Q(\ram[137][6] ), 
	.D(FE_PHN1519_n2780), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[137][5]  (.Q(\ram[137][5] ), 
	.D(FE_PHN373_n2779), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][4]  (.Q(\ram[137][4] ), 
	.D(FE_PHN303_n2778), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][3]  (.Q(\ram[137][3] ), 
	.D(FE_PHN1182_n2777), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][2]  (.Q(\ram[137][2] ), 
	.D(FE_PHN867_n2776), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[137][1]  (.Q(\ram[137][1] ), 
	.D(FE_PHN971_n2775), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[137][0]  (.Q(\ram[137][0] ), 
	.D(FE_PHN1471_n2774), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[133][15]  (.Q(\ram[133][15] ), 
	.D(FE_PHN1561_n2725), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][14]  (.Q(\ram[133][14] ), 
	.D(FE_PHN1180_n2724), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][13]  (.Q(\ram[133][13] ), 
	.D(FE_PHN2748_n2723), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][12]  (.Q(\ram[133][12] ), 
	.D(FE_PHN4603_n2722), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[133][11]  (.Q(\ram[133][11] ), 
	.D(FE_PHN589_n2721), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[133][10]  (.Q(\ram[133][10] ), 
	.D(FE_PHN398_n2720), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[133][9]  (.Q(\ram[133][9] ), 
	.D(n2719), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[133][8]  (.Q(\ram[133][8] ), 
	.D(FE_PHN496_n2718), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[133][7]  (.Q(\ram[133][7] ), 
	.D(FE_PHN813_n2717), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][6]  (.Q(\ram[133][6] ), 
	.D(FE_PHN2621_n2716), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][5]  (.Q(\ram[133][5] ), 
	.D(FE_PHN385_n2715), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][4]  (.Q(\ram[133][4] ), 
	.D(FE_PHN447_n2714), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[133][3]  (.Q(\ram[133][3] ), 
	.D(FE_PHN1095_n2713), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][2]  (.Q(\ram[133][2] ), 
	.D(FE_PHN189_n2712), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[133][1]  (.Q(\ram[133][1] ), 
	.D(FE_PHN443_n2711), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[133][0]  (.Q(\ram[133][0] ), 
	.D(FE_PHN634_n2710), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[129][15]  (.Q(\ram[129][15] ), 
	.D(FE_PHN2168_n2661), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][14]  (.Q(\ram[129][14] ), 
	.D(FE_PHN1640_n2660), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][13]  (.Q(\ram[129][13] ), 
	.D(FE_PHN2751_n2659), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][12]  (.Q(\ram[129][12] ), 
	.D(FE_PHN1266_n2658), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[129][11]  (.Q(\ram[129][11] ), 
	.D(FE_PHN1232_n2657), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[129][10]  (.Q(\ram[129][10] ), 
	.D(FE_PHN1479_n2656), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[129][9]  (.Q(\ram[129][9] ), 
	.D(FE_PHN651_n2655), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[129][8]  (.Q(\ram[129][8] ), 
	.D(FE_PHN490_n2654), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[129][7]  (.Q(\ram[129][7] ), 
	.D(n2653), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[129][6]  (.Q(\ram[129][6] ), 
	.D(FE_PHN247_n2652), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[129][5]  (.Q(\ram[129][5] ), 
	.D(FE_PHN221_n2651), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[129][4]  (.Q(\ram[129][4] ), 
	.D(FE_PHN1964_n2650), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[129][3]  (.Q(\ram[129][3] ), 
	.D(FE_PHN1034_n2649), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[129][2]  (.Q(\ram[129][2] ), 
	.D(FE_PHN475_n2648), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[129][1]  (.Q(\ram[129][1] ), 
	.D(FE_PHN351_n2647), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[129][0]  (.Q(\ram[129][0] ), 
	.D(FE_PHN2111_n2646), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[125][15]  (.Q(\ram[125][15] ), 
	.D(FE_PHN768_n2597), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][14]  (.Q(\ram[125][14] ), 
	.D(FE_PHN1717_n2596), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][13]  (.Q(\ram[125][13] ), 
	.D(FE_PHN1793_n2595), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][12]  (.Q(\ram[125][12] ), 
	.D(FE_PHN5721_n2594), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[125][11]  (.Q(\ram[125][11] ), 
	.D(FE_PHN1532_n2593), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[125][10]  (.Q(\ram[125][10] ), 
	.D(FE_PHN4870_n2592), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][9]  (.Q(\ram[125][9] ), 
	.D(FE_PHN1244_n2591), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[125][8]  (.Q(\ram[125][8] ), 
	.D(FE_PHN5672_n2590), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[125][7]  (.Q(\ram[125][7] ), 
	.D(FE_PHN5687_n2589), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][6]  (.Q(\ram[125][6] ), 
	.D(FE_PHN244_n2588), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][5]  (.Q(\ram[125][5] ), 
	.D(FE_PHN5748_n2587), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][4]  (.Q(\ram[125][4] ), 
	.D(FE_PHN612_n2586), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][3]  (.Q(\ram[125][3] ), 
	.D(FE_PHN599_n2585), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[125][2]  (.Q(\ram[125][2] ), 
	.D(FE_PHN1393_n2584), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[125][1]  (.Q(\ram[125][1] ), 
	.D(FE_PHN565_n2583), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[125][0]  (.Q(\ram[125][0] ), 
	.D(FE_PHN4847_n2582), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[121][15]  (.Q(\ram[121][15] ), 
	.D(FE_PHN949_n2533), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][14]  (.Q(\ram[121][14] ), 
	.D(FE_PHN646_n2532), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][13]  (.Q(\ram[121][13] ), 
	.D(FE_PHN427_n2531), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[121][12]  (.Q(\ram[121][12] ), 
	.D(FE_PHN1397_n2530), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][11]  (.Q(\ram[121][11] ), 
	.D(FE_PHN2038_n2529), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[121][10]  (.Q(\ram[121][10] ), 
	.D(FE_PHN2240_n2528), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][9]  (.Q(\ram[121][9] ), 
	.D(FE_PHN672_n2527), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][8]  (.Q(\ram[121][8] ), 
	.D(FE_PHN1027_n2526), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][7]  (.Q(\ram[121][7] ), 
	.D(FE_PHN1602_n2525), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[121][6]  (.Q(\ram[121][6] ), 
	.D(FE_PHN1172_n2524), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[121][5]  (.Q(\ram[121][5] ), 
	.D(FE_PHN293_n2523), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[121][4]  (.Q(\ram[121][4] ), 
	.D(FE_PHN2874_n2522), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[121][3]  (.Q(\ram[121][3] ), 
	.D(FE_PHN395_n2521), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[121][2]  (.Q(\ram[121][2] ), 
	.D(FE_PHN1325_n2520), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[121][1]  (.Q(\ram[121][1] ), 
	.D(FE_PHN656_n2519), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[121][0]  (.Q(\ram[121][0] ), 
	.D(FE_PHN930_n2518), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[117][15]  (.Q(\ram[117][15] ), 
	.D(FE_PHN1807_n2469), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[117][14]  (.Q(\ram[117][14] ), 
	.D(FE_PHN1563_n2468), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][13]  (.Q(\ram[117][13] ), 
	.D(FE_PHN270_n2467), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[117][12]  (.Q(\ram[117][12] ), 
	.D(FE_PHN2039_n2466), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[117][11]  (.Q(\ram[117][11] ), 
	.D(FE_PHN418_n2465), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][10]  (.Q(\ram[117][10] ), 
	.D(FE_PHN3053_n2464), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][9]  (.Q(\ram[117][9] ), 
	.D(FE_PHN650_n2463), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][8]  (.Q(\ram[117][8] ), 
	.D(FE_PHN2689_n2462), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][7]  (.Q(\ram[117][7] ), 
	.D(FE_PHN249_n2461), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][6]  (.Q(\ram[117][6] ), 
	.D(n2460), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[117][5]  (.Q(\ram[117][5] ), 
	.D(FE_PHN776_n2459), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[117][4]  (.Q(\ram[117][4] ), 
	.D(FE_PHN163_n2458), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[117][3]  (.Q(\ram[117][3] ), 
	.D(FE_PHN1213_n2457), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[117][2]  (.Q(\ram[117][2] ), 
	.D(FE_PHN501_n2456), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[117][1]  (.Q(\ram[117][1] ), 
	.D(FE_PHN252_n2455), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[117][0]  (.Q(\ram[117][0] ), 
	.D(FE_PHN946_n2454), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[113][15]  (.Q(\ram[113][15] ), 
	.D(FE_PHN4600_n2405), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[113][14]  (.Q(\ram[113][14] ), 
	.D(FE_PHN793_n2404), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[113][13]  (.Q(\ram[113][13] ), 
	.D(FE_PHN3605_n2403), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][12]  (.Q(\ram[113][12] ), 
	.D(FE_PHN6649_n2402), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[113][11]  (.Q(\ram[113][11] ), 
	.D(FE_PHN5647_n2401), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][10]  (.Q(\ram[113][10] ), 
	.D(FE_PHN3507_n2400), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][9]  (.Q(\ram[113][9] ), 
	.D(FE_PHN5035_n2399), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][8]  (.Q(\ram[113][8] ), 
	.D(FE_PHN5747_n2398), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][7]  (.Q(\ram[113][7] ), 
	.D(FE_PHN5770_n2397), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[113][6]  (.Q(\ram[113][6] ), 
	.D(FE_PHN3283_n2396), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][5]  (.Q(\ram[113][5] ), 
	.D(FE_PHN6646_n2395), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[113][4]  (.Q(\ram[113][4] ), 
	.D(FE_PHN6687_n2394), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][3]  (.Q(\ram[113][3] ), 
	.D(FE_PHN6663_n2393), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][2]  (.Q(\ram[113][2] ), 
	.D(FE_PHN321_n2392), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][1]  (.Q(\ram[113][1] ), 
	.D(FE_PHN4749_n2391), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[113][0]  (.Q(\ram[113][0] ), 
	.D(FE_PHN5752_n2390), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[109][15]  (.Q(\ram[109][15] ), 
	.D(FE_PHN306_n2341), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][14]  (.Q(\ram[109][14] ), 
	.D(FE_PHN269_n2340), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[109][13]  (.Q(\ram[109][13] ), 
	.D(FE_PHN2273_n2339), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[109][12]  (.Q(\ram[109][12] ), 
	.D(FE_PHN202_n2338), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[109][11]  (.Q(\ram[109][11] ), 
	.D(FE_PHN375_n2337), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[109][10]  (.Q(\ram[109][10] ), 
	.D(FE_PHN2425_n2336), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][9]  (.Q(\ram[109][9] ), 
	.D(FE_PHN2495_n2335), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[109][8]  (.Q(\ram[109][8] ), 
	.D(FE_PHN910_n2334), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][7]  (.Q(\ram[109][7] ), 
	.D(FE_PHN229_n2333), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[109][6]  (.Q(\ram[109][6] ), 
	.D(FE_PHN986_n2332), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][5]  (.Q(\ram[109][5] ), 
	.D(n2331), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[109][4]  (.Q(\ram[109][4] ), 
	.D(FE_PHN145_n2330), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[109][3]  (.Q(\ram[109][3] ), 
	.D(FE_PHN1950_n2329), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][2]  (.Q(\ram[109][2] ), 
	.D(FE_PHN2209_n2328), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][1]  (.Q(\ram[109][1] ), 
	.D(FE_PHN1642_n2327), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[109][0]  (.Q(\ram[109][0] ), 
	.D(FE_PHN2727_n2326), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[105][15]  (.Q(\ram[105][15] ), 
	.D(FE_PHN477_n2277), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][14]  (.Q(\ram[105][14] ), 
	.D(FE_PHN689_n2276), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][13]  (.Q(\ram[105][13] ), 
	.D(FE_PHN1610_n2275), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[105][12]  (.Q(\ram[105][12] ), 
	.D(FE_PHN425_n2274), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][11]  (.Q(\ram[105][11] ), 
	.D(FE_PHN124_n2273), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][10]  (.Q(\ram[105][10] ), 
	.D(FE_PHN1426_n2272), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[105][9]  (.Q(\ram[105][9] ), 
	.D(FE_PHN702_n2271), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][8]  (.Q(\ram[105][8] ), 
	.D(FE_PHN661_n2270), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[105][7]  (.Q(\ram[105][7] ), 
	.D(FE_PHN690_n2269), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[105][6]  (.Q(\ram[105][6] ), 
	.D(FE_PHN2107_n2268), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][5]  (.Q(\ram[105][5] ), 
	.D(FE_PHN1301_n2267), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][4]  (.Q(\ram[105][4] ), 
	.D(FE_PHN216_n2266), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[105][3]  (.Q(\ram[105][3] ), 
	.D(FE_PHN600_n2265), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[105][2]  (.Q(\ram[105][2] ), 
	.D(FE_PHN2433_n2264), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[105][1]  (.Q(\ram[105][1] ), 
	.D(FE_PHN1859_n2263), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[105][0]  (.Q(\ram[105][0] ), 
	.D(FE_PHN3613_n2262), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[101][15]  (.Q(\ram[101][15] ), 
	.D(FE_PHN1023_n2213), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[101][14]  (.Q(\ram[101][14] ), 
	.D(FE_PHN225_n2212), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][13]  (.Q(\ram[101][13] ), 
	.D(FE_PHN727_n2211), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[101][12]  (.Q(\ram[101][12] ), 
	.D(FE_PHN2790_n2210), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[101][11]  (.Q(\ram[101][11] ), 
	.D(FE_PHN2798_n2209), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[101][10]  (.Q(\ram[101][10] ), 
	.D(FE_PHN198_n2208), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][9]  (.Q(\ram[101][9] ), 
	.D(FE_PHN116_n2207), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][8]  (.Q(\ram[101][8] ), 
	.D(FE_PHN141_n2206), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][7]  (.Q(\ram[101][7] ), 
	.D(FE_PHN442_n2205), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[101][6]  (.Q(\ram[101][6] ), 
	.D(FE_PHN479_n2204), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][5]  (.Q(\ram[101][5] ), 
	.D(FE_PHN2236_n2203), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][4]  (.Q(\ram[101][4] ), 
	.D(FE_PHN2100_n2202), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[101][3]  (.Q(\ram[101][3] ), 
	.D(FE_PHN261_n2201), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[101][2]  (.Q(\ram[101][2] ), 
	.D(FE_PHN285_n2200), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[101][1]  (.Q(\ram[101][1] ), 
	.D(FE_PHN2104_n2199), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[101][0]  (.Q(\ram[101][0] ), 
	.D(FE_PHN1490_n2198), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[97][15]  (.Q(\ram[97][15] ), 
	.D(FE_PHN5679_n2149), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][14]  (.Q(\ram[97][14] ), 
	.D(FE_PHN5710_n2148), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][13]  (.Q(\ram[97][13] ), 
	.D(FE_PHN129_n2147), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[97][12]  (.Q(\ram[97][12] ), 
	.D(FE_PHN391_n2146), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[97][11]  (.Q(\ram[97][11] ), 
	.D(FE_PHN2368_n2145), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[97][10]  (.Q(\ram[97][10] ), 
	.D(FE_PHN4842_n2144), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[97][9]  (.Q(\ram[97][9] ), 
	.D(FE_PHN746_n2143), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[97][8]  (.Q(\ram[97][8] ), 
	.D(FE_PHN137_n2142), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][7]  (.Q(\ram[97][7] ), 
	.D(FE_PHN3262_n2141), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[97][6]  (.Q(\ram[97][6] ), 
	.D(FE_PHN308_n2140), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[97][5]  (.Q(\ram[97][5] ), 
	.D(FE_PHN664_n2139), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[97][4]  (.Q(\ram[97][4] ), 
	.D(FE_PHN5699_n2138), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[97][3]  (.Q(\ram[97][3] ), 
	.D(FE_PHN5653_n2137), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[97][2]  (.Q(\ram[97][2] ), 
	.D(FE_PHN133_n2136), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[97][1]  (.Q(\ram[97][1] ), 
	.D(FE_PHN6690_n2135), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[97][0]  (.Q(\ram[97][0] ), 
	.D(FE_PHN299_n2134), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[93][15]  (.Q(\ram[93][15] ), 
	.D(FE_PHN736_n2085), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][14]  (.Q(\ram[93][14] ), 
	.D(FE_PHN733_n2084), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][13]  (.Q(\ram[93][13] ), 
	.D(FE_PHN2989_n2083), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[93][12]  (.Q(\ram[93][12] ), 
	.D(FE_PHN1355_n2082), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][11]  (.Q(\ram[93][11] ), 
	.D(FE_PHN1295_n2081), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][10]  (.Q(\ram[93][10] ), 
	.D(FE_PHN2054_n2080), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[93][9]  (.Q(\ram[93][9] ), 
	.D(FE_PHN2723_n2079), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][8]  (.Q(\ram[93][8] ), 
	.D(FE_PHN2868_n2078), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[93][7]  (.Q(\ram[93][7] ), 
	.D(FE_PHN962_n2077), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][6]  (.Q(\ram[93][6] ), 
	.D(FE_PHN1980_n2076), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][5]  (.Q(\ram[93][5] ), 
	.D(FE_PHN1024_n2075), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][4]  (.Q(\ram[93][4] ), 
	.D(FE_PHN2490_n2074), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[93][3]  (.Q(\ram[93][3] ), 
	.D(n2073), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][2]  (.Q(\ram[93][2] ), 
	.D(FE_PHN1127_n2072), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[93][1]  (.Q(\ram[93][1] ), 
	.D(FE_PHN435_n2071), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[93][0]  (.Q(\ram[93][0] ), 
	.D(FE_PHN1092_n2070), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[89][15]  (.Q(\ram[89][15] ), 
	.D(FE_PHN2333_n2021), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][14]  (.Q(\ram[89][14] ), 
	.D(FE_PHN1614_n2020), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[89][13]  (.Q(\ram[89][13] ), 
	.D(FE_PHN1003_n2019), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][12]  (.Q(\ram[89][12] ), 
	.D(FE_PHN1181_n2018), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[89][11]  (.Q(\ram[89][11] ), 
	.D(FE_PHN525_n2017), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[89][10]  (.Q(\ram[89][10] ), 
	.D(FE_PHN2801_n2016), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][9]  (.Q(\ram[89][9] ), 
	.D(FE_PHN1715_n2015), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][8]  (.Q(\ram[89][8] ), 
	.D(FE_PHN1982_n2014), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][7]  (.Q(\ram[89][7] ), 
	.D(FE_PHN2122_n2013), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[89][6]  (.Q(\ram[89][6] ), 
	.D(FE_PHN3193_n2012), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][5]  (.Q(\ram[89][5] ), 
	.D(FE_PHN1489_n2011), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[89][4]  (.Q(\ram[89][4] ), 
	.D(FE_PHN1938_n2010), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][3]  (.Q(\ram[89][3] ), 
	.D(FE_PHN2231_n2009), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][2]  (.Q(\ram[89][2] ), 
	.D(FE_PHN2605_n2008), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[89][1]  (.Q(\ram[89][1] ), 
	.D(FE_PHN1632_n2007), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[89][0]  (.Q(\ram[89][0] ), 
	.D(FE_PHN1500_n2006), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[85][15]  (.Q(\ram[85][15] ), 
	.D(FE_PHN529_n1957), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][14]  (.Q(\ram[85][14] ), 
	.D(FE_PHN396_n1956), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][13]  (.Q(\ram[85][13] ), 
	.D(FE_PHN1442_n1955), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][12]  (.Q(\ram[85][12] ), 
	.D(FE_PHN1917_n1954), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][11]  (.Q(\ram[85][11] ), 
	.D(FE_PHN1194_n1953), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][10]  (.Q(\ram[85][10] ), 
	.D(n1952), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[85][9]  (.Q(\ram[85][9] ), 
	.D(FE_PHN1586_n1951), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][8]  (.Q(\ram[85][8] ), 
	.D(FE_PHN2591_n1950), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][7]  (.Q(\ram[85][7] ), 
	.D(FE_PHN1109_n1949), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[85][6]  (.Q(\ram[85][6] ), 
	.D(FE_PHN491_n1948), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[85][5]  (.Q(\ram[85][5] ), 
	.D(FE_PHN2123_n1947), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][4]  (.Q(\ram[85][4] ), 
	.D(FE_PHN2335_n1946), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][3]  (.Q(\ram[85][3] ), 
	.D(FE_PHN318_n1945), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][2]  (.Q(\ram[85][2] ), 
	.D(FE_PHN1674_n1944), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[85][1]  (.Q(\ram[85][1] ), 
	.D(FE_PHN1010_n1943), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[85][0]  (.Q(\ram[85][0] ), 
	.D(FE_PHN1688_n1942), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[81][15]  (.Q(\ram[81][15] ), 
	.D(FE_PHN1001_n1893), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][14]  (.Q(\ram[81][14] ), 
	.D(FE_PHN1407_n1892), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][13]  (.Q(\ram[81][13] ), 
	.D(n1891), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][12]  (.Q(\ram[81][12] ), 
	.D(FE_PHN916_n1890), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][11]  (.Q(\ram[81][11] ), 
	.D(FE_PHN686_n1889), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][10]  (.Q(\ram[81][10] ), 
	.D(FE_PHN1615_n1888), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[81][9]  (.Q(\ram[81][9] ), 
	.D(FE_PHN687_n1887), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[81][8]  (.Q(\ram[81][8] ), 
	.D(FE_PHN4246_n1886), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[81][7]  (.Q(\ram[81][7] ), 
	.D(FE_PHN739_n1885), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[81][6]  (.Q(\ram[81][6] ), 
	.D(FE_PHN1905_n1884), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][5]  (.Q(\ram[81][5] ), 
	.D(FE_PHN2413_n1883), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][4]  (.Q(\ram[81][4] ), 
	.D(FE_PHN807_n1882), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][3]  (.Q(\ram[81][3] ), 
	.D(FE_PHN1202_n1881), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[81][2]  (.Q(\ram[81][2] ), 
	.D(FE_PHN4370_n1880), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[81][1]  (.Q(\ram[81][1] ), 
	.D(n1879), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[81][0]  (.Q(\ram[81][0] ), 
	.D(FE_PHN582_n1878), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[77][15]  (.Q(\ram[77][15] ), 
	.D(FE_PHN3103_n1829), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][14]  (.Q(\ram[77][14] ), 
	.D(FE_PHN647_n1828), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][13]  (.Q(\ram[77][13] ), 
	.D(FE_PHN834_n1827), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][12]  (.Q(\ram[77][12] ), 
	.D(FE_PHN1664_n1826), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][11]  (.Q(\ram[77][11] ), 
	.D(FE_PHN3178_n1825), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][10]  (.Q(\ram[77][10] ), 
	.D(FE_PHN1035_n1824), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][9]  (.Q(\ram[77][9] ), 
	.D(FE_PHN2799_n1823), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][8]  (.Q(\ram[77][8] ), 
	.D(FE_PHN1567_n1822), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[77][7]  (.Q(\ram[77][7] ), 
	.D(FE_PHN602_n1821), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][6]  (.Q(\ram[77][6] ), 
	.D(FE_PHN710_n1820), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[77][5]  (.Q(\ram[77][5] ), 
	.D(FE_PHN1467_n1819), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][4]  (.Q(\ram[77][4] ), 
	.D(FE_PHN206_n1818), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][3]  (.Q(\ram[77][3] ), 
	.D(FE_PHN298_n1817), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[77][2]  (.Q(\ram[77][2] ), 
	.D(FE_PHN505_n1816), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[77][1]  (.Q(\ram[77][1] ), 
	.D(FE_PHN3214_n1815), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[77][0]  (.Q(\ram[77][0] ), 
	.D(FE_PHN258_n1814), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[73][15]  (.Q(\ram[73][15] ), 
	.D(FE_PHN480_n1765), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][14]  (.Q(\ram[73][14] ), 
	.D(FE_PHN468_n1764), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][13]  (.Q(\ram[73][13] ), 
	.D(FE_PHN1388_n1763), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[73][12]  (.Q(\ram[73][12] ), 
	.D(FE_PHN2359_n1762), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][11]  (.Q(\ram[73][11] ), 
	.D(FE_PHN235_n1761), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][10]  (.Q(\ram[73][10] ), 
	.D(FE_PHN606_n1760), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][9]  (.Q(\ram[73][9] ), 
	.D(FE_PHN2838_n1759), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][8]  (.Q(\ram[73][8] ), 
	.D(FE_PHN1242_n1758), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[73][7]  (.Q(\ram[73][7] ), 
	.D(FE_PHN3033_n1757), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][6]  (.Q(\ram[73][6] ), 
	.D(FE_PHN1989_n1756), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][5]  (.Q(\ram[73][5] ), 
	.D(FE_PHN2177_n1755), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][4]  (.Q(\ram[73][4] ), 
	.D(FE_PHN204_n1754), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[73][3]  (.Q(\ram[73][3] ), 
	.D(FE_PHN275_n1753), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[73][2]  (.Q(\ram[73][2] ), 
	.D(FE_PHN2911_n1752), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[73][1]  (.Q(\ram[73][1] ), 
	.D(FE_PHN792_n1751), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[73][0]  (.Q(\ram[73][0] ), 
	.D(FE_PHN2949_n1750), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[69][15]  (.Q(\ram[69][15] ), 
	.D(FE_PHN203_n1701), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[69][14]  (.Q(\ram[69][14] ), 
	.D(FE_PHN506_n1700), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][13]  (.Q(\ram[69][13] ), 
	.D(FE_PHN3153_n1699), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[69][12]  (.Q(\ram[69][12] ), 
	.D(FE_PHN1168_n1698), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][11]  (.Q(\ram[69][11] ), 
	.D(FE_PHN652_n1697), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][10]  (.Q(\ram[69][10] ), 
	.D(FE_PHN184_n1696), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][9]  (.Q(\ram[69][9] ), 
	.D(FE_PHN128_n1695), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][8]  (.Q(\ram[69][8] ), 
	.D(FE_PHN402_n1694), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][7]  (.Q(\ram[69][7] ), 
	.D(FE_PHN2403_n1693), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[69][6]  (.Q(\ram[69][6] ), 
	.D(FE_PHN107_n1692), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[69][5]  (.Q(\ram[69][5] ), 
	.D(FE_PHN251_n1691), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][4]  (.Q(\ram[69][4] ), 
	.D(FE_PHN543_n1690), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][3]  (.Q(\ram[69][3] ), 
	.D(FE_PHN1566_n1689), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[69][2]  (.Q(\ram[69][2] ), 
	.D(FE_PHN3208_n1688), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[69][1]  (.Q(\ram[69][1] ), 
	.D(FE_PHN2813_n1687), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[69][0]  (.Q(\ram[69][0] ), 
	.D(FE_PHN470_n1686), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[65][15]  (.Q(\ram[65][15] ), 
	.D(FE_PHN1574_n1637), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[65][14]  (.Q(\ram[65][14] ), 
	.D(FE_PHN2143_n1636), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][13]  (.Q(\ram[65][13] ), 
	.D(FE_PHN2102_n1635), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][12]  (.Q(\ram[65][12] ), 
	.D(FE_PHN144_n1634), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[65][11]  (.Q(\ram[65][11] ), 
	.D(FE_PHN1422_n1633), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][10]  (.Q(\ram[65][10] ), 
	.D(FE_PHN2210_n1632), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][9]  (.Q(\ram[65][9] ), 
	.D(FE_PHN1636_n1631), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][8]  (.Q(\ram[65][8] ), 
	.D(n1630), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][7]  (.Q(\ram[65][7] ), 
	.D(FE_PHN787_n1629), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[65][6]  (.Q(\ram[65][6] ), 
	.D(FE_PHN1018_n1628), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[65][5]  (.Q(\ram[65][5] ), 
	.D(FE_PHN929_n1627), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[65][4]  (.Q(\ram[65][4] ), 
	.D(FE_PHN277_n1626), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][3]  (.Q(\ram[65][3] ), 
	.D(FE_PHN1463_n1625), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[65][2]  (.Q(\ram[65][2] ), 
	.D(FE_PHN322_n1624), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[65][1]  (.Q(\ram[65][1] ), 
	.D(FE_PHN1520_n1623), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[65][0]  (.Q(\ram[65][0] ), 
	.D(FE_PHN335_n1622), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[61][15]  (.Q(\ram[61][15] ), 
	.D(FE_PHN2489_n1573), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][14]  (.Q(\ram[61][14] ), 
	.D(FE_PHN151_n1572), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[61][13]  (.Q(\ram[61][13] ), 
	.D(n1571), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[61][12]  (.Q(\ram[61][12] ), 
	.D(FE_PHN914_n1570), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][11]  (.Q(\ram[61][11] ), 
	.D(FE_PHN2796_n1569), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][10]  (.Q(\ram[61][10] ), 
	.D(FE_PHN2559_n1568), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][9]  (.Q(\ram[61][9] ), 
	.D(FE_PHN2096_n1567), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[61][8]  (.Q(\ram[61][8] ), 
	.D(FE_PHN1396_n1566), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][7]  (.Q(\ram[61][7] ), 
	.D(FE_PHN951_n1565), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][6]  (.Q(\ram[61][6] ), 
	.D(FE_PHN1919_n1564), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][5]  (.Q(\ram[61][5] ), 
	.D(FE_PHN1125_n1563), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][4]  (.Q(\ram[61][4] ), 
	.D(FE_PHN519_n1562), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][3]  (.Q(\ram[61][3] ), 
	.D(FE_PHN800_n1561), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[61][2]  (.Q(\ram[61][2] ), 
	.D(FE_PHN1797_n1560), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[61][1]  (.Q(\ram[61][1] ), 
	.D(FE_PHN641_n1559), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[61][0]  (.Q(\ram[61][0] ), 
	.D(FE_PHN1114_n1558), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[57][15]  (.Q(\ram[57][15] ), 
	.D(FE_PHN363_n1509), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[57][14]  (.Q(\ram[57][14] ), 
	.D(FE_PHN259_n1508), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[57][13]  (.Q(\ram[57][13] ), 
	.D(FE_PHN1011_n1507), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[57][12]  (.Q(\ram[57][12] ), 
	.D(FE_PHN984_n1506), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[57][11]  (.Q(\ram[57][11] ), 
	.D(FE_PHN1597_n1505), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][10]  (.Q(\ram[57][10] ), 
	.D(FE_PHN1647_n1504), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][9]  (.Q(\ram[57][9] ), 
	.D(FE_PHN1116_n1503), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[57][8]  (.Q(\ram[57][8] ), 
	.D(FE_PHN817_n1502), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[57][7]  (.Q(\ram[57][7] ), 
	.D(FE_PHN2756_n1501), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[57][6]  (.Q(\ram[57][6] ), 
	.D(FE_PHN1081_n1500), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][5]  (.Q(\ram[57][5] ), 
	.D(FE_PHN1653_n1499), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[57][4]  (.Q(\ram[57][4] ), 
	.D(FE_PHN2071_n1498), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[57][3]  (.Q(\ram[57][3] ), 
	.D(FE_PHN1937_n1497), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[57][2]  (.Q(\ram[57][2] ), 
	.D(FE_PHN677_n1496), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[57][1]  (.Q(\ram[57][1] ), 
	.D(FE_PHN1820_n1495), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[57][0]  (.Q(\ram[57][0] ), 
	.D(FE_PHN674_n1494), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[53][15]  (.Q(\ram[53][15] ), 
	.D(FE_PHN660_n1445), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][14]  (.Q(\ram[53][14] ), 
	.D(FE_PHN1083_n1444), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][13]  (.Q(\ram[53][13] ), 
	.D(FE_PHN510_n1443), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][12]  (.Q(\ram[53][12] ), 
	.D(FE_PHN1005_n1442), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][11]  (.Q(\ram[53][11] ), 
	.D(FE_PHN2289_n1441), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][10]  (.Q(\ram[53][10] ), 
	.D(FE_PHN809_n1440), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[53][9]  (.Q(\ram[53][9] ), 
	.D(FE_PHN931_n1439), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][8]  (.Q(\ram[53][8] ), 
	.D(FE_PHN2521_n1438), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][7]  (.Q(\ram[53][7] ), 
	.D(FE_PHN2379_n1437), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[53][6]  (.Q(\ram[53][6] ), 
	.D(FE_PHN2611_n1436), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[53][5]  (.Q(\ram[53][5] ), 
	.D(FE_PHN168_n1435), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[53][4]  (.Q(\ram[53][4] ), 
	.D(FE_PHN2461_n1434), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][3]  (.Q(\ram[53][3] ), 
	.D(FE_PHN918_n1433), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[53][2]  (.Q(\ram[53][2] ), 
	.D(FE_PHN1007_n1432), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][1]  (.Q(\ram[53][1] ), 
	.D(FE_PHN603_n1431), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[53][0]  (.Q(\ram[53][0] ), 
	.D(FE_PHN2892_n1430), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[49][15]  (.Q(\ram[49][15] ), 
	.D(FE_PHN2958_n1381), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[49][14]  (.Q(\ram[49][14] ), 
	.D(FE_PHN927_n1380), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[49][13]  (.Q(\ram[49][13] ), 
	.D(FE_PHN1236_n1379), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[49][12]  (.Q(\ram[49][12] ), 
	.D(FE_PHN1343_n1378), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][11]  (.Q(\ram[49][11] ), 
	.D(FE_PHN2009_n1377), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][10]  (.Q(\ram[49][10] ), 
	.D(FE_PHN3049_n1376), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][9]  (.Q(\ram[49][9] ), 
	.D(FE_PHN5760_n1375), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[49][8]  (.Q(\ram[49][8] ), 
	.D(FE_PHN2620_n1374), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[49][7]  (.Q(\ram[49][7] ), 
	.D(FE_PHN267_n1373), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[49][6]  (.Q(\ram[49][6] ), 
	.D(FE_PHN1892_n1372), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[49][5]  (.Q(\ram[49][5] ), 
	.D(FE_PHN1185_n1371), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][4]  (.Q(\ram[49][4] ), 
	.D(FE_PHN1146_n1370), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[49][3]  (.Q(\ram[49][3] ), 
	.D(FE_PHN290_n1369), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[49][2]  (.Q(\ram[49][2] ), 
	.D(FE_PHN1743_n1368), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[49][1]  (.Q(\ram[49][1] ), 
	.D(FE_PHN667_n1367), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[49][0]  (.Q(\ram[49][0] ), 
	.D(FE_PHN2344_n1366), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[45][15]  (.Q(\ram[45][15] ), 
	.D(FE_PHN1648_n1317), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][14]  (.Q(\ram[45][14] ), 
	.D(n1316), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][13]  (.Q(\ram[45][13] ), 
	.D(FE_PHN2258_n1315), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][12]  (.Q(\ram[45][12] ), 
	.D(FE_PHN2207_n1314), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][11]  (.Q(\ram[45][11] ), 
	.D(n1313), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][10]  (.Q(\ram[45][10] ), 
	.D(FE_PHN2059_n1312), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[45][9]  (.Q(\ram[45][9] ), 
	.D(FE_PHN2327_n1311), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][8]  (.Q(\ram[45][8] ), 
	.D(n1310), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[45][7]  (.Q(\ram[45][7] ), 
	.D(FE_PHN2888_n1309), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[45][6]  (.Q(\ram[45][6] ), 
	.D(FE_PHN1473_n1308), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][5]  (.Q(\ram[45][5] ), 
	.D(FE_PHN1529_n1307), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][4]  (.Q(\ram[45][4] ), 
	.D(FE_PHN2361_n1306), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][3]  (.Q(\ram[45][3] ), 
	.D(FE_PHN1789_n1305), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[45][2]  (.Q(\ram[45][2] ), 
	.D(FE_PHN2153_n1304), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[45][1]  (.Q(\ram[45][1] ), 
	.D(FE_PHN2301_n1303), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[45][0]  (.Q(\ram[45][0] ), 
	.D(n1302), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[41][15]  (.Q(\ram[41][15] ), 
	.D(FE_PHN1644_n1253), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][14]  (.Q(\ram[41][14] ), 
	.D(FE_PHN1691_n1252), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][13]  (.Q(\ram[41][13] ), 
	.D(FE_PHN1593_n1251), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[41][12]  (.Q(\ram[41][12] ), 
	.D(FE_PHN2185_n1250), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[41][11]  (.Q(\ram[41][11] ), 
	.D(FE_PHN654_n1249), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[41][10]  (.Q(\ram[41][10] ), 
	.D(FE_PHN1307_n1248), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][9]  (.Q(\ram[41][9] ), 
	.D(FE_PHN668_n1247), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][8]  (.Q(\ram[41][8] ), 
	.D(FE_PHN2127_n1246), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][7]  (.Q(\ram[41][7] ), 
	.D(FE_PHN1097_n1245), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[41][6]  (.Q(\ram[41][6] ), 
	.D(FE_PHN1732_n1244), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[41][5]  (.Q(\ram[41][5] ), 
	.D(FE_PHN2314_n1243), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[41][4]  (.Q(\ram[41][4] ), 
	.D(FE_PHN2526_n1242), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][3]  (.Q(\ram[41][3] ), 
	.D(FE_PHN1272_n1241), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[41][2]  (.Q(\ram[41][2] ), 
	.D(FE_PHN1277_n1240), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[41][1]  (.Q(\ram[41][1] ), 
	.D(FE_PHN226_n1239), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[41][0]  (.Q(\ram[41][0] ), 
	.D(FE_PHN1608_n1238), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[37][15]  (.Q(\ram[37][15] ), 
	.D(FE_PHN1579_n1189), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][14]  (.Q(\ram[37][14] ), 
	.D(FE_PHN875_n1188), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][13]  (.Q(\ram[37][13] ), 
	.D(FE_PHN822_n1187), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][12]  (.Q(\ram[37][12] ), 
	.D(FE_PHN580_n1186), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[37][11]  (.Q(\ram[37][11] ), 
	.D(FE_PHN1374_n1185), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[37][10]  (.Q(\ram[37][10] ), 
	.D(FE_PHN908_n1184), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[37][9]  (.Q(\ram[37][9] ), 
	.D(FE_PHN2357_n1183), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[37][8]  (.Q(\ram[37][8] ), 
	.D(FE_PHN1512_n1182), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][7]  (.Q(\ram[37][7] ), 
	.D(FE_PHN1683_n1181), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[37][6]  (.Q(\ram[37][6] ), 
	.D(FE_PHN1391_n1180), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[37][5]  (.Q(\ram[37][5] ), 
	.D(FE_PHN2080_n1179), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[37][4]  (.Q(\ram[37][4] ), 
	.D(FE_PHN5691_n1178), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[37][3]  (.Q(\ram[37][3] ), 
	.D(FE_PHN2563_n1177), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[37][2]  (.Q(\ram[37][2] ), 
	.D(FE_PHN637_n1176), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[37][1]  (.Q(\ram[37][1] ), 
	.D(FE_PHN678_n1175), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[37][0]  (.Q(\ram[37][0] ), 
	.D(FE_PHN1753_n1174), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[33][15]  (.Q(\ram[33][15] ), 
	.D(FE_PHN1444_n1125), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[33][14]  (.Q(\ram[33][14] ), 
	.D(FE_PHN985_n1124), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][13]  (.Q(\ram[33][13] ), 
	.D(FE_PHN1287_n1123), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[33][12]  (.Q(\ram[33][12] ), 
	.D(FE_PHN1815_n1122), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][11]  (.Q(\ram[33][11] ), 
	.D(FE_PHN211_n1121), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][10]  (.Q(\ram[33][10] ), 
	.D(FE_PHN2237_n1120), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[33][9]  (.Q(\ram[33][9] ), 
	.D(n1119), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[33][8]  (.Q(\ram[33][8] ), 
	.D(FE_PHN3145_n1118), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][7]  (.Q(\ram[33][7] ), 
	.D(FE_PHN2863_n1117), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[33][6]  (.Q(\ram[33][6] ), 
	.D(FE_PHN635_n1116), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][5]  (.Q(\ram[33][5] ), 
	.D(FE_PHN2406_n1115), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][4]  (.Q(\ram[33][4] ), 
	.D(FE_PHN1558_n1114), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][3]  (.Q(\ram[33][3] ), 
	.D(FE_PHN1079_n1113), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[33][2]  (.Q(\ram[33][2] ), 
	.D(FE_PHN176_n1112), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[33][1]  (.Q(\ram[33][1] ), 
	.D(FE_PHN3050_n1111), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[33][0]  (.Q(\ram[33][0] ), 
	.D(FE_PHN4586_n1110), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[29][15]  (.Q(\ram[29][15] ), 
	.D(FE_PHN268_n1061), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[29][14]  (.Q(\ram[29][14] ), 
	.D(n1060), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][13]  (.Q(\ram[29][13] ), 
	.D(FE_PHN449_n1059), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[29][12]  (.Q(\ram[29][12] ), 
	.D(FE_PHN123_n1058), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[29][11]  (.Q(\ram[29][11] ), 
	.D(FE_PHN752_n1057), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][10]  (.Q(\ram[29][10] ), 
	.D(FE_PHN4130_n1056), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[29][9]  (.Q(\ram[29][9] ), 
	.D(FE_PHN509_n1055), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][8]  (.Q(\ram[29][8] ), 
	.D(FE_PHN5683_n1054), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][7]  (.Q(\ram[29][7] ), 
	.D(FE_PHN182_n1053), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][6]  (.Q(\ram[29][6] ), 
	.D(FE_PHN717_n1052), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][5]  (.Q(\ram[29][5] ), 
	.D(FE_PHN4392_n1051), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][4]  (.Q(\ram[29][4] ), 
	.D(FE_PHN2441_n1050), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[29][3]  (.Q(\ram[29][3] ), 
	.D(FE_PHN152_n1049), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[29][2]  (.Q(\ram[29][2] ), 
	.D(FE_PHN4051_n1048), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[29][1]  (.Q(\ram[29][1] ), 
	.D(FE_PHN294_n1047), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[29][0]  (.Q(\ram[29][0] ), 
	.D(FE_PHN4750_n1046), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][15]  (.Q(\ram[25][15] ), 
	.D(FE_PHN4452_n997), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[25][14]  (.Q(\ram[25][14] ), 
	.D(FE_PHN4894_n996), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][13]  (.Q(\ram[25][13] ), 
	.D(FE_PHN1420_n995), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[25][12]  (.Q(\ram[25][12] ), 
	.D(FE_PHN5249_n994), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][11]  (.Q(\ram[25][11] ), 
	.D(FE_PHN4607_n993), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[25][10]  (.Q(\ram[25][10] ), 
	.D(FE_PHN5092_n992), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][9]  (.Q(\ram[25][9] ), 
	.D(FE_PHN4577_n991), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[25][8]  (.Q(\ram[25][8] ), 
	.D(FE_PHN423_n990), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[25][7]  (.Q(\ram[25][7] ), 
	.D(FE_PHN3560_n989), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][6]  (.Q(\ram[25][6] ), 
	.D(FE_PHN4443_n988), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[25][5]  (.Q(\ram[25][5] ), 
	.D(FE_PHN365_n987), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[25][4]  (.Q(\ram[25][4] ), 
	.D(FE_PHN4565_n986), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][3]  (.Q(\ram[25][3] ), 
	.D(FE_PHN4867_n985), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[25][2]  (.Q(\ram[25][2] ), 
	.D(FE_PHN4054_n984), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[25][1]  (.Q(\ram[25][1] ), 
	.D(FE_PHN5733_n983), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[25][0]  (.Q(\ram[25][0] ), 
	.D(FE_PHN4326_n982), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[21][15]  (.Q(\ram[21][15] ), 
	.D(FE_PHN4340_n933), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[21][14]  (.Q(\ram[21][14] ), 
	.D(FE_PHN888_n932), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][13]  (.Q(\ram[21][13] ), 
	.D(FE_PHN585_n931), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[21][12]  (.Q(\ram[21][12] ), 
	.D(FE_PHN4150_n930), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[21][11]  (.Q(\ram[21][11] ), 
	.D(FE_PHN4311_n929), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][10]  (.Q(\ram[21][10] ), 
	.D(FE_PHN4147_n928), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[21][9]  (.Q(\ram[21][9] ), 
	.D(FE_PHN4208_n927), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][8]  (.Q(\ram[21][8] ), 
	.D(FE_PHN1043_n926), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[21][7]  (.Q(\ram[21][7] ), 
	.D(FE_PHN4118_n925), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][6]  (.Q(\ram[21][6] ), 
	.D(FE_PHN2429_n924), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[21][5]  (.Q(\ram[21][5] ), 
	.D(FE_PHN1899_n923), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[21][4]  (.Q(\ram[21][4] ), 
	.D(FE_PHN4192_n922), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[21][3]  (.Q(\ram[21][3] ), 
	.D(FE_PHN5759_n921), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[21][2]  (.Q(\ram[21][2] ), 
	.D(FE_PHN5040_n920), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[21][1]  (.Q(\ram[21][1] ), 
	.D(FE_PHN4144_n919), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[21][0]  (.Q(\ram[21][0] ), 
	.D(FE_PHN5514_n918), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[17][15]  (.Q(\ram[17][15] ), 
	.D(FE_PHN3335_n869), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[17][14]  (.Q(\ram[17][14] ), 
	.D(n868), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][13]  (.Q(\ram[17][13] ), 
	.D(FE_PHN424_n867), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][12]  (.Q(\ram[17][12] ), 
	.D(FE_PHN3395_n866), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][11]  (.Q(\ram[17][11] ), 
	.D(FE_PHN4128_n865), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][10]  (.Q(\ram[17][10] ), 
	.D(FE_PHN3279_n864), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[17][9]  (.Q(\ram[17][9] ), 
	.D(FE_PHN4711_n863), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][8]  (.Q(\ram[17][8] ), 
	.D(FE_PHN416_n862), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[17][7]  (.Q(\ram[17][7] ), 
	.D(FE_PHN4444_n861), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[17][6]  (.Q(\ram[17][6] ), 
	.D(FE_PHN764_n860), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[17][5]  (.Q(\ram[17][5] ), 
	.D(FE_PHN816_n859), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[17][4]  (.Q(\ram[17][4] ), 
	.D(FE_PHN4587_n858), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[17][3]  (.Q(\ram[17][3] ), 
	.D(FE_PHN4121_n857), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][2]  (.Q(\ram[17][2] ), 
	.D(FE_PHN5422_n856), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[17][1]  (.Q(\ram[17][1] ), 
	.D(FE_PHN4083_n855), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[17][0]  (.Q(\ram[17][0] ), 
	.D(FE_PHN4697_n854), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[13][15]  (.Q(\ram[13][15] ), 
	.D(FE_PHN1230_n805), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[13][14]  (.Q(\ram[13][14] ), 
	.D(FE_PHN401_n804), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[13][13]  (.Q(\ram[13][13] ), 
	.D(FE_PHN2932_n803), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][12]  (.Q(\ram[13][12] ), 
	.D(FE_PHN552_n802), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[13][11]  (.Q(\ram[13][11] ), 
	.D(FE_PHN3158_n801), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][10]  (.Q(\ram[13][10] ), 
	.D(FE_PHN893_n800), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[13][9]  (.Q(\ram[13][9] ), 
	.D(FE_PHN2722_n799), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[13][8]  (.Q(\ram[13][8] ), 
	.D(FE_PHN1305_n798), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][7]  (.Q(\ram[13][7] ), 
	.D(FE_PHN372_n797), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[13][6]  (.Q(\ram[13][6] ), 
	.D(FE_PHN406_n796), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][5]  (.Q(\ram[13][5] ), 
	.D(FE_PHN2846_n795), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][4]  (.Q(\ram[13][4] ), 
	.D(FE_PHN2445_n794), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][3]  (.Q(\ram[13][3] ), 
	.D(FE_PHN546_n793), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[13][2]  (.Q(\ram[13][2] ), 
	.D(FE_PHN1856_n792), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[13][1]  (.Q(\ram[13][1] ), 
	.D(FE_PHN232_n791), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[13][0]  (.Q(\ram[13][0] ), 
	.D(FE_PHN1400_n790), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][15]  (.Q(\ram[9][15] ), 
	.D(FE_PHN854_n741), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][14]  (.Q(\ram[9][14] ), 
	.D(FE_PHN574_n740), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[9][13]  (.Q(\ram[9][13] ), 
	.D(FE_PHN2278_n739), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[9][12]  (.Q(\ram[9][12] ), 
	.D(FE_PHN2400_n738), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][11]  (.Q(\ram[9][11] ), 
	.D(FE_PHN420_n737), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][10]  (.Q(\ram[9][10] ), 
	.D(FE_PHN512_n736), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][9]  (.Q(\ram[9][9] ), 
	.D(FE_PHN192_n735), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][8]  (.Q(\ram[9][8] ), 
	.D(FE_PHN551_n734), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][7]  (.Q(\ram[9][7] ), 
	.D(FE_PHN718_n733), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][6]  (.Q(\ram[9][6] ), 
	.D(FE_PHN2376_n732), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][5]  (.Q(\ram[9][5] ), 
	.D(FE_PHN2654_n731), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[9][4]  (.Q(\ram[9][4] ), 
	.D(FE_PHN1414_n730), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][3]  (.Q(\ram[9][3] ), 
	.D(FE_PHN3027_n729), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[9][2]  (.Q(\ram[9][2] ), 
	.D(FE_PHN729_n728), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[9][1]  (.Q(\ram[9][1] ), 
	.D(n727), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[9][0]  (.Q(\ram[9][0] ), 
	.D(FE_PHN1803_n726), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[5][15]  (.Q(\ram[5][15] ), 
	.D(FE_PHN2262_n677), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][14]  (.Q(\ram[5][14] ), 
	.D(FE_PHN1696_n676), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][13]  (.Q(\ram[5][13] ), 
	.D(FE_PHN2212_n675), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[5][12]  (.Q(\ram[5][12] ), 
	.D(FE_PHN1737_n674), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[5][11]  (.Q(\ram[5][11] ), 
	.D(FE_PHN2346_n673), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[5][10]  (.Q(\ram[5][10] ), 
	.D(FE_PHN1113_n672), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][9]  (.Q(\ram[5][9] ), 
	.D(FE_PHN1611_n671), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[5][8]  (.Q(\ram[5][8] ), 
	.D(FE_PHN1772_n670), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][7]  (.Q(\ram[5][7] ), 
	.D(FE_PHN2088_n669), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][6]  (.Q(\ram[5][6] ), 
	.D(FE_PHN2138_n668), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[5][5]  (.Q(\ram[5][5] ), 
	.D(FE_PHN2099_n667), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[5][4]  (.Q(\ram[5][4] ), 
	.D(FE_PHN632_n666), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][3]  (.Q(\ram[5][3] ), 
	.D(FE_PHN1673_n665), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[5][2]  (.Q(\ram[5][2] ), 
	.D(FE_PHN2720_n664), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[5][1]  (.Q(\ram[5][1] ), 
	.D(FE_PHN1046_n663), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[5][0]  (.Q(\ram[5][0] ), 
	.D(FE_PHN969_n662), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[1][15]  (.Q(\ram[1][15] ), 
	.D(FE_PHN2931_n613), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[1][14]  (.Q(\ram[1][14] ), 
	.D(FE_PHN876_n612), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[1][13]  (.Q(\ram[1][13] ), 
	.D(FE_PHN1546_n611), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[1][12]  (.Q(\ram[1][12] ), 
	.D(FE_PHN528_n610), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[1][11]  (.Q(\ram[1][11] ), 
	.D(FE_PHN399_n609), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[1][10]  (.Q(\ram[1][10] ), 
	.D(FE_PHN1759_n608), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[1][9]  (.Q(\ram[1][9] ), 
	.D(FE_PHN1066_n607), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[1][8]  (.Q(\ram[1][8] ), 
	.D(FE_PHN922_n606), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[1][7]  (.Q(\ram[1][7] ), 
	.D(FE_PHN1316_n605), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[1][6]  (.Q(\ram[1][6] ), 
	.D(FE_PHN2232_n604), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[1][5]  (.Q(\ram[1][5] ), 
	.D(FE_PHN757_n603), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[1][4]  (.Q(\ram[1][4] ), 
	.D(FE_PHN601_n602), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[1][3]  (.Q(\ram[1][3] ), 
	.D(FE_PHN376_n601), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[1][2]  (.Q(\ram[1][2] ), 
	.D(FE_PHN2073_n600), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[1][1]  (.Q(\ram[1][1] ), 
	.D(FE_PHN2215_n599), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[1][0]  (.Q(\ram[1][0] ), 
	.D(FE_PHN2588_n598), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[254][15]  (.Q(\ram[254][15] ), 
	.D(FE_PHN2062_n4661), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[254][14]  (.Q(\ram[254][14] ), 
	.D(FE_PHN1590_n4660), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[254][13]  (.Q(\ram[254][13] ), 
	.D(FE_PHN722_n4659), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[254][12]  (.Q(\ram[254][12] ), 
	.D(FE_PHN287_n4658), 
	.CK(clk));
   QDFFEHD \ram_reg[254][11]  (.Q(\ram[254][11] ), 
	.D(FE_PHN1405_n4657), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][10]  (.Q(\ram[254][10] ), 
	.D(FE_PHN1267_n4656), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[254][9]  (.Q(\ram[254][9] ), 
	.D(n4655), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][8]  (.Q(\ram[254][8] ), 
	.D(FE_PHN2208_n4654), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][7]  (.Q(\ram[254][7] ), 
	.D(FE_PHN1584_n4653), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[254][6]  (.Q(\ram[254][6] ), 
	.D(FE_PHN1382_n4652), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[254][5]  (.Q(\ram[254][5] ), 
	.D(FE_PHN801_n4651), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[254][4]  (.Q(\ram[254][4] ), 
	.D(FE_PHN1870_n4650), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[254][3]  (.Q(\ram[254][3] ), 
	.D(FE_PHN2152_n4649), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[254][2]  (.Q(\ram[254][2] ), 
	.D(FE_PHN2007_n4648), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[254][1]  (.Q(\ram[254][1] ), 
	.D(FE_PHN2017_n4647), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[254][0]  (.Q(\ram[254][0] ), 
	.D(FE_PHN991_n4646), 
	.CK(clk));
   QDFFEHD \ram_reg[250][15]  (.Q(\ram[250][15] ), 
	.D(FE_PHN2307_n4597), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][14]  (.Q(\ram[250][14] ), 
	.D(FE_PHN2349_n4596), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][13]  (.Q(\ram[250][13] ), 
	.D(FE_PHN902_n4595), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[250][12]  (.Q(\ram[250][12] ), 
	.D(FE_PHN1554_n4594), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][11]  (.Q(\ram[250][11] ), 
	.D(FE_PHN1087_n4593), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][10]  (.Q(\ram[250][10] ), 
	.D(FE_PHN1569_n4592), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][9]  (.Q(\ram[250][9] ), 
	.D(FE_PHN1710_n4591), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[250][8]  (.Q(\ram[250][8] ), 
	.D(FE_PHN626_n4590), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[250][7]  (.Q(\ram[250][7] ), 
	.D(FE_PHN452_n4589), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][6]  (.Q(\ram[250][6] ), 
	.D(FE_PHN1061_n4588), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[250][5]  (.Q(\ram[250][5] ), 
	.D(FE_PHN195_n4587), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][4]  (.Q(\ram[250][4] ), 
	.D(FE_PHN1712_n4586), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[250][3]  (.Q(\ram[250][3] ), 
	.D(FE_PHN2049_n4585), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[250][2]  (.Q(\ram[250][2] ), 
	.D(FE_PHN1735_n4584), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[250][1]  (.Q(\ram[250][1] ), 
	.D(n4583), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[250][0]  (.Q(\ram[250][0] ), 
	.D(FE_PHN169_n4582), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[246][15]  (.Q(\ram[246][15] ), 
	.D(FE_PHN272_n4533), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[246][14]  (.Q(\ram[246][14] ), 
	.D(FE_PHN684_n4532), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[246][13]  (.Q(\ram[246][13] ), 
	.D(FE_PHN1276_n4531), 
	.CK(clk));
   QDFFEHD \ram_reg[246][12]  (.Q(\ram[246][12] ), 
	.D(FE_PHN1718_n4530), 
	.CK(clk));
   QDFFEHD \ram_reg[246][11]  (.Q(\ram[246][11] ), 
	.D(FE_PHN1705_n4529), 
	.CK(clk));
   QDFFEHD \ram_reg[246][10]  (.Q(\ram[246][10] ), 
	.D(FE_PHN921_n4528), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][9]  (.Q(\ram[246][9] ), 
	.D(FE_PHN441_n4527), 
	.CK(clk));
   QDFFEHD \ram_reg[246][8]  (.Q(\ram[246][8] ), 
	.D(FE_PHN1869_n4526), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][7]  (.Q(\ram[246][7] ), 
	.D(FE_PHN387_n4525), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[246][6]  (.Q(\ram[246][6] ), 
	.D(FE_PHN953_n4524), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[246][5]  (.Q(\ram[246][5] ), 
	.D(FE_PHN849_n4523), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][4]  (.Q(\ram[246][4] ), 
	.D(FE_PHN148_n4522), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[246][3]  (.Q(\ram[246][3] ), 
	.D(FE_PHN794_n4521), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[246][2]  (.Q(\ram[246][2] ), 
	.D(FE_PHN1805_n4520), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[246][1]  (.Q(\ram[246][1] ), 
	.D(FE_PHN720_n4519), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[246][0]  (.Q(\ram[246][0] ), 
	.D(FE_PHN724_n4518), 
	.CK(clk));
   QDFFEHD \ram_reg[242][15]  (.Q(\ram[242][15] ), 
	.D(FE_PHN2341_n4469), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[242][14]  (.Q(\ram[242][14] ), 
	.D(FE_PHN1689_n4468), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][13]  (.Q(\ram[242][13] ), 
	.D(FE_PHN1748_n4467), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][12]  (.Q(\ram[242][12] ), 
	.D(FE_PHN598_n4466), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][11]  (.Q(\ram[242][11] ), 
	.D(FE_PHN291_n4465), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][10]  (.Q(\ram[242][10] ), 
	.D(FE_PHN2820_n4464), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][9]  (.Q(\ram[242][9] ), 
	.D(FE_PHN1697_n4463), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][8]  (.Q(\ram[242][8] ), 
	.D(FE_PHN2904_n4462), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[242][7]  (.Q(\ram[242][7] ), 
	.D(FE_PHN549_n4461), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][6]  (.Q(\ram[242][6] ), 
	.D(FE_PHN2862_n4460), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][5]  (.Q(\ram[242][5] ), 
	.D(FE_PHN670_n4459), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][4]  (.Q(\ram[242][4] ), 
	.D(FE_PHN1389_n4458), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][3]  (.Q(\ram[242][3] ), 
	.D(FE_PHN2308_n4457), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[242][2]  (.Q(\ram[242][2] ), 
	.D(FE_PHN180_n4456), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][1]  (.Q(\ram[242][1] ), 
	.D(FE_PHN1303_n4455), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[242][0]  (.Q(\ram[242][0] ), 
	.D(FE_PHN1885_n4454), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[238][15]  (.Q(\ram[238][15] ), 
	.D(FE_PHN4055_n4405), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][14]  (.Q(\ram[238][14] ), 
	.D(FE_PHN4453_n4404), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][13]  (.Q(\ram[238][13] ), 
	.D(FE_PHN4518_n4403), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][12]  (.Q(\ram[238][12] ), 
	.D(FE_PHN4695_n4402), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][11]  (.Q(\ram[238][11] ), 
	.D(FE_PHN4567_n4401), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][10]  (.Q(\ram[238][10] ), 
	.D(FE_PHN4500_n4400), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[238][9]  (.Q(\ram[238][9] ), 
	.D(FE_PHN4021_n4399), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[238][8]  (.Q(\ram[238][8] ), 
	.D(FE_PHN3331_n4398), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][7]  (.Q(\ram[238][7] ), 
	.D(FE_PHN4386_n4397), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[238][6]  (.Q(\ram[238][6] ), 
	.D(FE_PHN4638_n4396), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[238][5]  (.Q(\ram[238][5] ), 
	.D(FE_PHN4732_n4395), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[238][4]  (.Q(\ram[238][4] ), 
	.D(FE_PHN4510_n4394), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][3]  (.Q(\ram[238][3] ), 
	.D(FE_PHN4481_n4393), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[238][2]  (.Q(\ram[238][2] ), 
	.D(FE_PHN4650_n4392), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[238][1]  (.Q(\ram[238][1] ), 
	.D(FE_PHN4484_n4391), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[238][0]  (.Q(\ram[238][0] ), 
	.D(n4390), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[234][15]  (.Q(\ram[234][15] ), 
	.D(FE_PHN2873_n4341), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[234][14]  (.Q(\ram[234][14] ), 
	.D(FE_PHN3537_n4340), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[234][13]  (.Q(\ram[234][13] ), 
	.D(FE_PHN3256_n4339), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[234][12]  (.Q(\ram[234][12] ), 
	.D(FE_PHN5118_n4338), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[234][11]  (.Q(\ram[234][11] ), 
	.D(FE_PHN855_n4337), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][10]  (.Q(\ram[234][10] ), 
	.D(FE_PHN1880_n4336), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][9]  (.Q(\ram[234][9] ), 
	.D(FE_PHN1472_n4335), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][8]  (.Q(\ram[234][8] ), 
	.D(FE_PHN4473_n4334), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][7]  (.Q(\ram[234][7] ), 
	.D(FE_PHN4352_n4333), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][6]  (.Q(\ram[234][6] ), 
	.D(FE_PHN4308_n4332), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[234][5]  (.Q(\ram[234][5] ), 
	.D(FE_PHN4188_n4331), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[234][4]  (.Q(\ram[234][4] ), 
	.D(FE_PHN2728_n4330), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[234][3]  (.Q(\ram[234][3] ), 
	.D(FE_PHN4706_n4329), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[234][2]  (.Q(\ram[234][2] ), 
	.D(FE_PHN309_n4328), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[234][1]  (.Q(\ram[234][1] ), 
	.D(FE_PHN4229_n4327), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[234][0]  (.Q(\ram[234][0] ), 
	.D(FE_PHN358_n4326), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[230][15]  (.Q(\ram[230][15] ), 
	.D(FE_PHN4568_n4277), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[230][14]  (.Q(\ram[230][14] ), 
	.D(FE_PHN4690_n4276), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[230][13]  (.Q(\ram[230][13] ), 
	.D(FE_PHN500_n4275), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[230][12]  (.Q(\ram[230][12] ), 
	.D(FE_PHN4256_n4274), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[230][11]  (.Q(\ram[230][11] ), 
	.D(FE_PHN4464_n4273), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][10]  (.Q(\ram[230][10] ), 
	.D(FE_PHN954_n4272), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][9]  (.Q(\ram[230][9] ), 
	.D(FE_PHN4387_n4271), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][8]  (.Q(\ram[230][8] ), 
	.D(FE_PHN4456_n4270), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][7]  (.Q(\ram[230][7] ), 
	.D(FE_PHN5527_n4269), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][6]  (.Q(\ram[230][6] ), 
	.D(FE_PHN4635_n4268), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[230][5]  (.Q(\ram[230][5] ), 
	.D(FE_PHN4730_n4267), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[230][4]  (.Q(\ram[230][4] ), 
	.D(FE_PHN4407_n4266), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[230][3]  (.Q(\ram[230][3] ), 
	.D(FE_PHN4740_n4265), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[230][2]  (.Q(\ram[230][2] ), 
	.D(FE_PHN1247_n4264), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[230][1]  (.Q(\ram[230][1] ), 
	.D(FE_PHN4094_n4263), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[230][0]  (.Q(\ram[230][0] ), 
	.D(FE_PHN4719_n4262), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[226][15]  (.Q(\ram[226][15] ), 
	.D(FE_PHN3644_n4213), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][14]  (.Q(\ram[226][14] ), 
	.D(FE_PHN4633_n4212), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][13]  (.Q(\ram[226][13] ), 
	.D(FE_PHN4569_n4211), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[226][12]  (.Q(\ram[226][12] ), 
	.D(FE_PHN3930_n4210), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[226][11]  (.Q(\ram[226][11] ), 
	.D(FE_PHN4700_n4209), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][10]  (.Q(\ram[226][10] ), 
	.D(FE_PHN2992_n4208), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[226][9]  (.Q(\ram[226][9] ), 
	.D(FE_PHN4726_n4207), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][8]  (.Q(\ram[226][8] ), 
	.D(FE_PHN4417_n4206), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][7]  (.Q(\ram[226][7] ), 
	.D(FE_PHN2614_n4205), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[226][6]  (.Q(\ram[226][6] ), 
	.D(FE_PHN5308_n4204), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[226][5]  (.Q(\ram[226][5] ), 
	.D(FE_PHN3249_n4203), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][4]  (.Q(\ram[226][4] ), 
	.D(FE_PHN4714_n4202), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[226][3]  (.Q(\ram[226][3] ), 
	.D(FE_PHN3383_n4201), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][2]  (.Q(\ram[226][2] ), 
	.D(FE_PHN1916_n4200), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[226][1]  (.Q(\ram[226][1] ), 
	.D(FE_PHN4485_n4199), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[226][0]  (.Q(\ram[226][0] ), 
	.D(FE_PHN846_n4198), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[222][15]  (.Q(\ram[222][15] ), 
	.D(FE_PHN2267_n4149), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[222][14]  (.Q(\ram[222][14] ), 
	.D(FE_PHN4547_n4148), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[222][13]  (.Q(\ram[222][13] ), 
	.D(FE_PHN6669_n4147), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][12]  (.Q(\ram[222][12] ), 
	.D(FE_PHN5003_n4146), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][11]  (.Q(\ram[222][11] ), 
	.D(FE_PHN1766_n4145), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[222][10]  (.Q(\ram[222][10] ), 
	.D(FE_PHN2299_n4144), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[222][9]  (.Q(\ram[222][9] ), 
	.D(FE_PHN3079_n4143), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][8]  (.Q(\ram[222][8] ), 
	.D(FE_PHN4086_n4142), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][7]  (.Q(\ram[222][7] ), 
	.D(FE_PHN2941_n4141), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[222][6]  (.Q(\ram[222][6] ), 
	.D(FE_PHN1605_n4140), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][5]  (.Q(\ram[222][5] ), 
	.D(FE_PHN6659_n4139), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][4]  (.Q(\ram[222][4] ), 
	.D(FE_PHN4109_n4138), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[222][3]  (.Q(\ram[222][3] ), 
	.D(FE_PHN4832_n4137), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][2]  (.Q(\ram[222][2] ), 
	.D(FE_PHN863_n4136), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[222][1]  (.Q(\ram[222][1] ), 
	.D(FE_PHN5763_n4135), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[222][0]  (.Q(\ram[222][0] ), 
	.D(FE_PHN3823_n4134), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[218][15]  (.Q(\ram[218][15] ), 
	.D(FE_PHN850_n4085), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][14]  (.Q(\ram[218][14] ), 
	.D(FE_PHN187_n4084), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][13]  (.Q(\ram[218][13] ), 
	.D(FE_PHN758_n4083), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][12]  (.Q(\ram[218][12] ), 
	.D(FE_PHN2125_n4082), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[218][11]  (.Q(\ram[218][11] ), 
	.D(FE_PHN273_n4081), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][10]  (.Q(\ram[218][10] ), 
	.D(FE_PHN604_n4080), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][9]  (.Q(\ram[218][9] ), 
	.D(FE_PHN2560_n4079), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[218][8]  (.Q(\ram[218][8] ), 
	.D(FE_PHN1336_n4078), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[218][7]  (.Q(\ram[218][7] ), 
	.D(FE_PHN2370_n4077), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][6]  (.Q(\ram[218][6] ), 
	.D(FE_PHN4739_n4076), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][5]  (.Q(\ram[218][5] ), 
	.D(FE_PHN2280_n4075), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[218][4]  (.Q(\ram[218][4] ), 
	.D(FE_PHN1965_n4074), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[218][3]  (.Q(\ram[218][3] ), 
	.D(FE_PHN2334_n4073), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[218][2]  (.Q(\ram[218][2] ), 
	.D(FE_PHN765_n4072), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][1]  (.Q(\ram[218][1] ), 
	.D(FE_PHN1009_n4071), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[218][0]  (.Q(\ram[218][0] ), 
	.D(FE_PHN518_n4070), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[214][15]  (.Q(\ram[214][15] ), 
	.D(FE_PHN4583_n4021), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][14]  (.Q(\ram[214][14] ), 
	.D(FE_PHN223_n4020), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][13]  (.Q(\ram[214][13] ), 
	.D(n4019), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][12]  (.Q(\ram[214][12] ), 
	.D(FE_PHN5695_n4018), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][11]  (.Q(\ram[214][11] ), 
	.D(FE_PHN4416_n4017), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][10]  (.Q(\ram[214][10] ), 
	.D(FE_PHN4615_n4016), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][9]  (.Q(\ram[214][9] ), 
	.D(FE_PHN4746_n4015), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][8]  (.Q(\ram[214][8] ), 
	.D(FE_PHN5174_n4014), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][7]  (.Q(\ram[214][7] ), 
	.D(FE_PHN4877_n4013), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][6]  (.Q(\ram[214][6] ), 
	.D(FE_PHN5732_n4012), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][5]  (.Q(\ram[214][5] ), 
	.D(FE_PHN6642_n4011), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[214][4]  (.Q(\ram[214][4] ), 
	.D(FE_PHN4255_n4010), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[214][3]  (.Q(\ram[214][3] ), 
	.D(FE_PHN4139_n4009), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][2]  (.Q(\ram[214][2] ), 
	.D(FE_PHN4133_n4008), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[214][1]  (.Q(\ram[214][1] ), 
	.D(FE_PHN4176_n4007), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[214][0]  (.Q(\ram[214][0] ), 
	.D(FE_PHN4100_n4006), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[210][15]  (.Q(\ram[210][15] ), 
	.D(FE_PHN286_n3957), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[210][14]  (.Q(\ram[210][14] ), 
	.D(FE_PHN4715_n3956), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[210][13]  (.Q(\ram[210][13] ), 
	.D(FE_PHN4327_n3955), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][12]  (.Q(\ram[210][12] ), 
	.D(FE_PHN5486_n3954), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][11]  (.Q(\ram[210][11] ), 
	.D(FE_PHN6700_n3953), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][10]  (.Q(\ram[210][10] ), 
	.D(FE_PHN4735_n3952), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][9]  (.Q(\ram[210][9] ), 
	.D(FE_PHN4738_n3951), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][8]  (.Q(\ram[210][8] ), 
	.D(FE_PHN4743_n3950), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][7]  (.Q(\ram[210][7] ), 
	.D(FE_PHN1337_n3949), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][6]  (.Q(\ram[210][6] ), 
	.D(FE_PHN4089_n3948), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][5]  (.Q(\ram[210][5] ), 
	.D(FE_PHN4991_n3947), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[210][4]  (.Q(\ram[210][4] ), 
	.D(FE_PHN4298_n3946), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[210][3]  (.Q(\ram[210][3] ), 
	.D(FE_PHN4657_n3945), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[210][2]  (.Q(\ram[210][2] ), 
	.D(FE_PHN5670_n3944), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[210][1]  (.Q(\ram[210][1] ), 
	.D(FE_PHN5413_n3943), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[210][0]  (.Q(\ram[210][0] ), 
	.D(FE_PHN4522_n3942), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[206][15]  (.Q(\ram[206][15] ), 
	.D(FE_PHN2680_n3893), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][14]  (.Q(\ram[206][14] ), 
	.D(FE_PHN2663_n3892), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[206][13]  (.Q(\ram[206][13] ), 
	.D(FE_PHN3155_n3891), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[206][12]  (.Q(\ram[206][12] ), 
	.D(FE_PHN1370_n3890), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[206][11]  (.Q(\ram[206][11] ), 
	.D(FE_PHN2221_n3889), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][10]  (.Q(\ram[206][10] ), 
	.D(FE_PHN433_n3888), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[206][9]  (.Q(\ram[206][9] ), 
	.D(FE_PHN583_n3887), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[206][8]  (.Q(\ram[206][8] ), 
	.D(FE_PHN1419_n3886), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[206][7]  (.Q(\ram[206][7] ), 
	.D(FE_PHN741_n3885), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[206][6]  (.Q(\ram[206][6] ), 
	.D(FE_PHN1935_n3884), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[206][5]  (.Q(\ram[206][5] ), 
	.D(FE_PHN965_n3883), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[206][4]  (.Q(\ram[206][4] ), 
	.D(FE_PHN658_n3882), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][3]  (.Q(\ram[206][3] ), 
	.D(FE_PHN539_n3881), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[206][2]  (.Q(\ram[206][2] ), 
	.D(FE_PHN1289_n3880), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[206][1]  (.Q(\ram[206][1] ), 
	.D(FE_PHN862_n3879), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[206][0]  (.Q(\ram[206][0] ), 
	.D(FE_PHN2576_n3878), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[202][15]  (.Q(\ram[202][15] ), 
	.D(FE_PHN903_n3829), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][14]  (.Q(\ram[202][14] ), 
	.D(FE_PHN866_n3828), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][13]  (.Q(\ram[202][13] ), 
	.D(n3827), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[202][12]  (.Q(\ram[202][12] ), 
	.D(FE_PHN2927_n3826), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][11]  (.Q(\ram[202][11] ), 
	.D(FE_PHN1652_n3825), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][10]  (.Q(\ram[202][10] ), 
	.D(FE_PHN1994_n3824), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][9]  (.Q(\ram[202][9] ), 
	.D(FE_PHN1435_n3823), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][8]  (.Q(\ram[202][8] ), 
	.D(FE_PHN952_n3822), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[202][7]  (.Q(\ram[202][7] ), 
	.D(FE_PHN1160_n3821), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][6]  (.Q(\ram[202][6] ), 
	.D(FE_PHN1143_n3820), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[202][5]  (.Q(\ram[202][5] ), 
	.D(FE_PHN550_n3819), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[202][4]  (.Q(\ram[202][4] ), 
	.D(FE_PHN2450_n3818), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][3]  (.Q(\ram[202][3] ), 
	.D(FE_PHN257_n3817), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][2]  (.Q(\ram[202][2] ), 
	.D(FE_PHN2996_n3816), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[202][1]  (.Q(\ram[202][1] ), 
	.D(FE_PHN1292_n3815), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[202][0]  (.Q(\ram[202][0] ), 
	.D(FE_PHN1050_n3814), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[198][15]  (.Q(\ram[198][15] ), 
	.D(FE_PHN2662_n3765), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][14]  (.Q(\ram[198][14] ), 
	.D(FE_PHN2036_n3764), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][13]  (.Q(\ram[198][13] ), 
	.D(FE_PHN547_n3763), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][12]  (.Q(\ram[198][12] ), 
	.D(FE_PHN382_n3762), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][11]  (.Q(\ram[198][11] ), 
	.D(FE_PHN891_n3761), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][10]  (.Q(\ram[198][10] ), 
	.D(FE_PHN852_n3760), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][9]  (.Q(\ram[198][9] ), 
	.D(FE_PHN699_n3759), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[198][8]  (.Q(\ram[198][8] ), 
	.D(FE_PHN1078_n3758), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][7]  (.Q(\ram[198][7] ), 
	.D(FE_PHN419_n3757), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][6]  (.Q(\ram[198][6] ), 
	.D(FE_PHN2512_n3756), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][5]  (.Q(\ram[198][5] ), 
	.D(FE_PHN1445_n3755), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][4]  (.Q(\ram[198][4] ), 
	.D(FE_PHN179_n3754), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[198][3]  (.Q(\ram[198][3] ), 
	.D(FE_PHN1522_n3753), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[198][2]  (.Q(\ram[198][2] ), 
	.D(FE_PHN1163_n3752), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][1]  (.Q(\ram[198][1] ), 
	.D(FE_PHN2233_n3751), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[198][0]  (.Q(\ram[198][0] ), 
	.D(FE_PHN2337_n3750), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[194][15]  (.Q(\ram[194][15] ), 
	.D(FE_PHN2274_n3701), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][14]  (.Q(\ram[194][14] ), 
	.D(FE_PHN2109_n3700), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][13]  (.Q(\ram[194][13] ), 
	.D(FE_PHN769_n3699), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[194][12]  (.Q(\ram[194][12] ), 
	.D(FE_PHN1315_n3698), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][11]  (.Q(\ram[194][11] ), 
	.D(FE_PHN3115_n3697), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][10]  (.Q(\ram[194][10] ), 
	.D(FE_PHN1514_n3696), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[194][9]  (.Q(\ram[194][9] ), 
	.D(FE_PHN1750_n3695), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][8]  (.Q(\ram[194][8] ), 
	.D(FE_PHN560_n3694), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[194][7]  (.Q(\ram[194][7] ), 
	.D(FE_PHN2503_n3693), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][6]  (.Q(\ram[194][6] ), 
	.D(FE_PHN2582_n3692), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][5]  (.Q(\ram[194][5] ), 
	.D(FE_PHN1356_n3691), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][4]  (.Q(\ram[194][4] ), 
	.D(FE_PHN1595_n3690), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][3]  (.Q(\ram[194][3] ), 
	.D(FE_PHN2569_n3689), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[194][2]  (.Q(\ram[194][2] ), 
	.D(FE_PHN3197_n3688), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[194][1]  (.Q(\ram[194][1] ), 
	.D(FE_PHN1129_n3687), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[194][0]  (.Q(\ram[194][0] ), 
	.D(FE_PHN2248_n3686), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[190][15]  (.Q(\ram[190][15] ), 
	.D(FE_PHN1926_n3637), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][14]  (.Q(\ram[190][14] ), 
	.D(FE_PHN1177_n3636), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][13]  (.Q(\ram[190][13] ), 
	.D(FE_PHN2940_n3635), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[190][12]  (.Q(\ram[190][12] ), 
	.D(FE_PHN3051_n3634), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[190][11]  (.Q(\ram[190][11] ), 
	.D(FE_PHN438_n3633), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][10]  (.Q(\ram[190][10] ), 
	.D(FE_PHN228_n3632), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][9]  (.Q(\ram[190][9] ), 
	.D(FE_PHN2834_n3631), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][8]  (.Q(\ram[190][8] ), 
	.D(FE_PHN2402_n3630), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[190][7]  (.Q(\ram[190][7] ), 
	.D(FE_PHN370_n3629), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][6]  (.Q(\ram[190][6] ), 
	.D(FE_PHN912_n3628), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[190][5]  (.Q(\ram[190][5] ), 
	.D(FE_PHN1730_n3627), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[190][4]  (.Q(\ram[190][4] ), 
	.D(FE_PHN2866_n3626), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][3]  (.Q(\ram[190][3] ), 
	.D(FE_PHN413_n3625), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[190][2]  (.Q(\ram[190][2] ), 
	.D(FE_PHN2772_n3624), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][1]  (.Q(\ram[190][1] ), 
	.D(FE_PHN1096_n3623), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[190][0]  (.Q(\ram[190][0] ), 
	.D(FE_PHN2580_n3622), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[186][15]  (.Q(\ram[186][15] ), 
	.D(FE_PHN723_n3573), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][14]  (.Q(\ram[186][14] ), 
	.D(FE_PHN238_n3572), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][13]  (.Q(\ram[186][13] ), 
	.D(FE_PHN1384_n3571), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][12]  (.Q(\ram[186][12] ), 
	.D(FE_PHN484_n3570), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[186][11]  (.Q(\ram[186][11] ), 
	.D(FE_PHN1549_n3569), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][10]  (.Q(\ram[186][10] ), 
	.D(FE_PHN108_n3568), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[186][9]  (.Q(\ram[186][9] ), 
	.D(FE_PHN2602_n3567), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[186][8]  (.Q(\ram[186][8] ), 
	.D(FE_PHN1164_n3566), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[186][7]  (.Q(\ram[186][7] ), 
	.D(FE_PHN214_n3565), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][6]  (.Q(\ram[186][6] ), 
	.D(FE_PHN150_n3564), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][5]  (.Q(\ram[186][5] ), 
	.D(FE_PHN158_n3563), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][4]  (.Q(\ram[186][4] ), 
	.D(FE_PHN304_n3562), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[186][3]  (.Q(\ram[186][3] ), 
	.D(FE_PHN170_n3561), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[186][2]  (.Q(\ram[186][2] ), 
	.D(FE_PHN571_n3560), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][1]  (.Q(\ram[186][1] ), 
	.D(FE_PHN1866_n3559), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[186][0]  (.Q(\ram[186][0] ), 
	.D(FE_PHN103_n3558), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[182][15]  (.Q(\ram[182][15] ), 
	.D(FE_PHN586_n3509), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[182][14]  (.Q(\ram[182][14] ), 
	.D(FE_PHN296_n3508), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[182][13]  (.Q(\ram[182][13] ), 
	.D(FE_PHN2447_n3507), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[182][12]  (.Q(\ram[182][12] ), 
	.D(FE_PHN2296_n3506), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[182][11]  (.Q(\ram[182][11] ), 
	.D(FE_PHN960_n3505), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[182][10]  (.Q(\ram[182][10] ), 
	.D(FE_PHN2520_n3504), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[182][9]  (.Q(\ram[182][9] ), 
	.D(FE_PHN2967_n3503), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[182][8]  (.Q(\ram[182][8] ), 
	.D(FE_PHN1895_n3502), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[182][7]  (.Q(\ram[182][7] ), 
	.D(FE_PHN643_n3501), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[182][6]  (.Q(\ram[182][6] ), 
	.D(FE_PHN2444_n3500), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[182][5]  (.Q(\ram[182][5] ), 
	.D(FE_PHN156_n3499), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[182][4]  (.Q(\ram[182][4] ), 
	.D(FE_PHN692_n3498), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[182][3]  (.Q(\ram[182][3] ), 
	.D(FE_PHN515_n3497), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[182][2]  (.Q(\ram[182][2] ), 
	.D(FE_PHN1949_n3496), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[182][1]  (.Q(\ram[182][1] ), 
	.D(FE_PHN1699_n3495), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[182][0]  (.Q(\ram[182][0] ), 
	.D(FE_PHN1604_n3494), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[178][15]  (.Q(\ram[178][15] ), 
	.D(FE_PHN2759_n3445), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][14]  (.Q(\ram[178][14] ), 
	.D(FE_PHN1830_n3444), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][13]  (.Q(\ram[178][13] ), 
	.D(FE_PHN3008_n3443), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][12]  (.Q(\ram[178][12] ), 
	.D(FE_PHN2199_n3442), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][11]  (.Q(\ram[178][11] ), 
	.D(FE_PHN957_n3441), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][10]  (.Q(\ram[178][10] ), 
	.D(FE_PHN2977_n3440), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[178][9]  (.Q(\ram[178][9] ), 
	.D(FE_PHN1728_n3439), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][8]  (.Q(\ram[178][8] ), 
	.D(FE_PHN595_n3438), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][7]  (.Q(\ram[178][7] ), 
	.D(FE_PHN2536_n3437), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][6]  (.Q(\ram[178][6] ), 
	.D(FE_PHN1831_n3436), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][5]  (.Q(\ram[178][5] ), 
	.D(FE_PHN2363_n3435), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][4]  (.Q(\ram[178][4] ), 
	.D(FE_PHN2375_n3434), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][3]  (.Q(\ram[178][3] ), 
	.D(FE_PHN2856_n3433), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[178][2]  (.Q(\ram[178][2] ), 
	.D(FE_PHN2466_n3432), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[178][1]  (.Q(\ram[178][1] ), 
	.D(FE_PHN2089_n3431), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[178][0]  (.Q(\ram[178][0] ), 
	.D(FE_PHN2742_n3430), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[174][15]  (.Q(\ram[174][15] ), 
	.D(FE_PHN1910_n3381), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][14]  (.Q(\ram[174][14] ), 
	.D(FE_PHN280_n3380), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][13]  (.Q(\ram[174][13] ), 
	.D(FE_PHN1583_n3379), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[174][12]  (.Q(\ram[174][12] ), 
	.D(FE_PHN2443_n3378), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[174][11]  (.Q(\ram[174][11] ), 
	.D(FE_PHN2775_n3377), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[174][10]  (.Q(\ram[174][10] ), 
	.D(FE_PHN2642_n3376), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[174][9]  (.Q(\ram[174][9] ), 
	.D(FE_PHN459_n3375), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][8]  (.Q(\ram[174][8] ), 
	.D(FE_PHN2352_n3374), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][7]  (.Q(\ram[174][7] ), 
	.D(FE_PHN1094_n3373), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][6]  (.Q(\ram[174][6] ), 
	.D(FE_PHN2915_n3372), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[174][5]  (.Q(\ram[174][5] ), 
	.D(FE_PHN1670_n3371), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][4]  (.Q(\ram[174][4] ), 
	.D(FE_PHN2913_n3370), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][3]  (.Q(\ram[174][3] ), 
	.D(FE_PHN1851_n3369), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[174][2]  (.Q(\ram[174][2] ), 
	.D(FE_PHN1261_n3368), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][1]  (.Q(\ram[174][1] ), 
	.D(FE_PHN379_n3367), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[174][0]  (.Q(\ram[174][0] ), 
	.D(FE_PHN770_n3366), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[170][15]  (.Q(\ram[170][15] ), 
	.D(FE_PHN1565_n3317), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][14]  (.Q(\ram[170][14] ), 
	.D(FE_PHN1708_n3316), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][13]  (.Q(\ram[170][13] ), 
	.D(FE_PHN1255_n3315), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][12]  (.Q(\ram[170][12] ), 
	.D(FE_PHN1555_n3314), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][11]  (.Q(\ram[170][11] ), 
	.D(FE_PHN644_n3313), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][10]  (.Q(\ram[170][10] ), 
	.D(FE_PHN645_n3312), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][9]  (.Q(\ram[170][9] ), 
	.D(FE_PHN942_n3311), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][8]  (.Q(\ram[170][8] ), 
	.D(FE_PHN2463_n3310), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][7]  (.Q(\ram[170][7] ), 
	.D(FE_PHN2129_n3309), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][6]  (.Q(\ram[170][6] ), 
	.D(FE_PHN2535_n3308), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][5]  (.Q(\ram[170][5] ), 
	.D(FE_PHN851_n3307), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][4]  (.Q(\ram[170][4] ), 
	.D(FE_PHN785_n3306), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[170][3]  (.Q(\ram[170][3] ), 
	.D(FE_PHN1537_n3305), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][2]  (.Q(\ram[170][2] ), 
	.D(FE_PHN1155_n3304), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[170][1]  (.Q(\ram[170][1] ), 
	.D(FE_PHN1319_n3303), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[170][0]  (.Q(\ram[170][0] ), 
	.D(FE_PHN2567_n3302), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[166][15]  (.Q(\ram[166][15] ), 
	.D(FE_PHN2047_n3253), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[166][14]  (.Q(\ram[166][14] ), 
	.D(FE_PHN2585_n3252), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][13]  (.Q(\ram[166][13] ), 
	.D(FE_PHN1592_n3251), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[166][12]  (.Q(\ram[166][12] ), 
	.D(FE_PHN2787_n3250), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][11]  (.Q(\ram[166][11] ), 
	.D(FE_PHN1704_n3249), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][10]  (.Q(\ram[166][10] ), 
	.D(FE_PHN882_n3248), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[166][9]  (.Q(\ram[166][9] ), 
	.D(FE_PHN1927_n3247), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][8]  (.Q(\ram[166][8] ), 
	.D(FE_PHN573_n3246), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][7]  (.Q(\ram[166][7] ), 
	.D(FE_PHN640_n3245), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[166][6]  (.Q(\ram[166][6] ), 
	.D(FE_PHN790_n3244), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][5]  (.Q(\ram[166][5] ), 
	.D(FE_PHN3139_n3243), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][4]  (.Q(\ram[166][4] ), 
	.D(FE_PHN2455_n3242), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[166][3]  (.Q(\ram[166][3] ), 
	.D(FE_PHN3694_n3241), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][2]  (.Q(\ram[166][2] ), 
	.D(FE_PHN1849_n3240), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[166][1]  (.Q(\ram[166][1] ), 
	.D(FE_PHN217_n3239), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[166][0]  (.Q(\ram[166][0] ), 
	.D(FE_PHN773_n3238), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][15]  (.Q(\ram[162][15] ), 
	.D(FE_PHN1228_n3189), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][14]  (.Q(\ram[162][14] ), 
	.D(FE_PHN1577_n3188), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][13]  (.Q(\ram[162][13] ), 
	.D(FE_PHN1630_n3187), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][12]  (.Q(\ram[162][12] ), 
	.D(FE_PHN2257_n3186), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][11]  (.Q(\ram[162][11] ), 
	.D(FE_PHN2538_n3185), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][10]  (.Q(\ram[162][10] ), 
	.D(FE_PHN1838_n3184), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][9]  (.Q(\ram[162][9] ), 
	.D(FE_PHN1548_n3183), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[162][8]  (.Q(\ram[162][8] ), 
	.D(FE_PHN2584_n3182), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[162][7]  (.Q(\ram[162][7] ), 
	.D(FE_PHN1904_n3181), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][6]  (.Q(\ram[162][6] ), 
	.D(FE_PHN1695_n3180), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][5]  (.Q(\ram[162][5] ), 
	.D(FE_PHN2853_n3179), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][4]  (.Q(\ram[162][4] ), 
	.D(FE_PHN1811_n3178), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][3]  (.Q(\ram[162][3] ), 
	.D(FE_PHN1900_n3177), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[162][2]  (.Q(\ram[162][2] ), 
	.D(FE_PHN859_n3176), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[162][1]  (.Q(\ram[162][1] ), 
	.D(FE_PHN2703_n3175), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[162][0]  (.Q(\ram[162][0] ), 
	.D(FE_PHN2050_n3174), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[158][15]  (.Q(\ram[158][15] ), 
	.D(FE_PHN4011_n3125), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][14]  (.Q(\ram[158][14] ), 
	.D(FE_PHN4096_n3124), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][13]  (.Q(\ram[158][13] ), 
	.D(FE_PHN4223_n3123), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][12]  (.Q(\ram[158][12] ), 
	.D(FE_PHN4360_n3122), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[158][11]  (.Q(\ram[158][11] ), 
	.D(n3121), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][10]  (.Q(\ram[158][10] ), 
	.D(FE_PHN4439_n3120), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[158][9]  (.Q(\ram[158][9] ), 
	.D(FE_PHN4541_n3119), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[158][8]  (.Q(\ram[158][8] ), 
	.D(FE_PHN4061_n3118), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[158][7]  (.Q(\ram[158][7] ), 
	.D(FE_PHN4268_n3117), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[158][6]  (.Q(\ram[158][6] ), 
	.D(FE_PHN5451_n3116), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[158][5]  (.Q(\ram[158][5] ), 
	.D(FE_PHN4141_n3115), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[158][4]  (.Q(\ram[158][4] ), 
	.D(FE_PHN4254_n3114), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[158][3]  (.Q(\ram[158][3] ), 
	.D(FE_PHN675_n3113), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[158][2]  (.Q(\ram[158][2] ), 
	.D(FE_PHN5424_n3112), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[158][1]  (.Q(\ram[158][1] ), 
	.D(FE_PHN4189_n3111), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[158][0]  (.Q(\ram[158][0] ), 
	.D(FE_PHN5460_n3110), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[154][15]  (.Q(\ram[154][15] ), 
	.D(FE_PHN706_n3061), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[154][14]  (.Q(\ram[154][14] ), 
	.D(FE_PHN5404_n3060), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[154][13]  (.Q(\ram[154][13] ), 
	.D(FE_PHN649_n3059), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[154][12]  (.Q(\ram[154][12] ), 
	.D(FE_PHN5493_n3058), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[154][11]  (.Q(\ram[154][11] ), 
	.D(FE_PHN1119_n3057), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[154][10]  (.Q(\ram[154][10] ), 
	.D(FE_PHN4162_n3056), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[154][9]  (.Q(\ram[154][9] ), 
	.D(FE_PHN4396_n3055), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[154][8]  (.Q(\ram[154][8] ), 
	.D(FE_PHN4323_n3054), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[154][7]  (.Q(\ram[154][7] ), 
	.D(FE_PHN4151_n3053), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][6]  (.Q(\ram[154][6] ), 
	.D(FE_PHN3532_n3052), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][5]  (.Q(\ram[154][5] ), 
	.D(n3051), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][4]  (.Q(\ram[154][4] ), 
	.D(FE_PHN4382_n3050), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[154][3]  (.Q(\ram[154][3] ), 
	.D(FE_PHN3419_n3049), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][2]  (.Q(\ram[154][2] ), 
	.D(FE_PHN3418_n3048), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[154][1]  (.Q(\ram[154][1] ), 
	.D(FE_PHN4875_n3047), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[154][0]  (.Q(\ram[154][0] ), 
	.D(FE_PHN4299_n3046), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[150][15]  (.Q(\ram[150][15] ), 
	.D(FE_PHN4409_n2997), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][14]  (.Q(\ram[150][14] ), 
	.D(FE_PHN4505_n2996), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][13]  (.Q(\ram[150][13] ), 
	.D(FE_PHN3880_n2995), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][12]  (.Q(\ram[150][12] ), 
	.D(FE_PHN4107_n2994), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][11]  (.Q(\ram[150][11] ), 
	.D(FE_PHN4405_n2993), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][10]  (.Q(\ram[150][10] ), 
	.D(FE_PHN3572_n2992), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[150][9]  (.Q(\ram[150][9] ), 
	.D(FE_PHN4097_n2991), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[150][8]  (.Q(\ram[150][8] ), 
	.D(FE_PHN4742_n2990), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[150][7]  (.Q(\ram[150][7] ), 
	.D(FE_PHN4579_n2989), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][6]  (.Q(\ram[150][6] ), 
	.D(FE_PHN4312_n2988), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[150][5]  (.Q(\ram[150][5] ), 
	.D(FE_PHN4630_n2987), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][4]  (.Q(\ram[150][4] ), 
	.D(FE_PHN4608_n2986), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[150][3]  (.Q(\ram[150][3] ), 
	.D(FE_PHN4259_n2985), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][2]  (.Q(\ram[150][2] ), 
	.D(FE_PHN4654_n2984), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[150][1]  (.Q(\ram[150][1] ), 
	.D(FE_PHN4612_n2983), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[150][0]  (.Q(\ram[150][0] ), 
	.D(FE_PHN4200_n2982), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[146][15]  (.Q(\ram[146][15] ), 
	.D(FE_PHN4534_n2933), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[146][14]  (.Q(\ram[146][14] ), 
	.D(FE_PHN5152_n2932), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[146][13]  (.Q(\ram[146][13] ), 
	.D(FE_PHN1233_n2931), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[146][12]  (.Q(\ram[146][12] ), 
	.D(FE_PHN4448_n2930), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[146][11]  (.Q(\ram[146][11] ), 
	.D(FE_PHN2367_n2929), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[146][10]  (.Q(\ram[146][10] ), 
	.D(FE_PHN4712_n2928), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[146][9]  (.Q(\ram[146][9] ), 
	.D(FE_PHN4617_n2927), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[146][8]  (.Q(\ram[146][8] ), 
	.D(FE_PHN3444_n2926), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[146][7]  (.Q(\ram[146][7] ), 
	.D(FE_PHN5734_n2925), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[146][6]  (.Q(\ram[146][6] ), 
	.D(FE_PHN1075_n2924), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][5]  (.Q(\ram[146][5] ), 
	.D(FE_PHN4762_n2923), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][4]  (.Q(\ram[146][4] ), 
	.D(FE_PHN4401_n2922), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[146][3]  (.Q(\ram[146][3] ), 
	.D(FE_PHN5764_n2921), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][2]  (.Q(\ram[146][2] ), 
	.D(FE_PHN4701_n2920), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[146][1]  (.Q(\ram[146][1] ), 
	.D(FE_PHN5749_n2919), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[146][0]  (.Q(\ram[146][0] ), 
	.D(FE_PHN4710_n2918), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[142][15]  (.Q(\ram[142][15] ), 
	.D(FE_PHN2960_n2869), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[142][14]  (.Q(\ram[142][14] ), 
	.D(FE_PHN3118_n2868), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[142][13]  (.Q(\ram[142][13] ), 
	.D(FE_PHN2239_n2867), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[142][12]  (.Q(\ram[142][12] ), 
	.D(FE_PHN974_n2866), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[142][11]  (.Q(\ram[142][11] ), 
	.D(FE_PHN2281_n2865), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[142][10]  (.Q(\ram[142][10] ), 
	.D(FE_PHN1591_n2864), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[142][9]  (.Q(\ram[142][9] ), 
	.D(FE_PHN2474_n2863), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[142][8]  (.Q(\ram[142][8] ), 
	.D(FE_PHN1193_n2862), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[142][7]  (.Q(\ram[142][7] ), 
	.D(FE_PHN2224_n2861), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[142][6]  (.Q(\ram[142][6] ), 
	.D(FE_PHN1613_n2860), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[142][5]  (.Q(\ram[142][5] ), 
	.D(FE_PHN588_n2859), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[142][4]  (.Q(\ram[142][4] ), 
	.D(FE_PHN1104_n2858), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[142][3]  (.Q(\ram[142][3] ), 
	.D(FE_PHN5673_n2857), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[142][2]  (.Q(\ram[142][2] ), 
	.D(FE_PHN975_n2856), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[142][1]  (.Q(\ram[142][1] ), 
	.D(FE_PHN1716_n2855), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[142][0]  (.Q(\ram[142][0] ), 
	.D(FE_PHN2189_n2854), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[138][15]  (.Q(\ram[138][15] ), 
	.D(FE_PHN219_n2805), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][14]  (.Q(\ram[138][14] ), 
	.D(FE_PHN2999_n2804), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][13]  (.Q(\ram[138][13] ), 
	.D(FE_PHN222_n2803), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[138][12]  (.Q(\ram[138][12] ), 
	.D(FE_PHN3104_n2802), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][11]  (.Q(\ram[138][11] ), 
	.D(FE_PHN346_n2801), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][10]  (.Q(\ram[138][10] ), 
	.D(FE_PHN1439_n2800), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][9]  (.Q(\ram[138][9] ), 
	.D(FE_PHN791_n2799), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[138][8]  (.Q(\ram[138][8] ), 
	.D(FE_PHN2690_n2798), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[138][7]  (.Q(\ram[138][7] ), 
	.D(FE_PHN812_n2797), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][6]  (.Q(\ram[138][6] ), 
	.D(FE_PHN274_n2796), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][5]  (.Q(\ram[138][5] ), 
	.D(FE_PHN2414_n2795), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][4]  (.Q(\ram[138][4] ), 
	.D(FE_PHN1208_n2794), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][3]  (.Q(\ram[138][3] ), 
	.D(FE_PHN2954_n2793), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][2]  (.Q(\ram[138][2] ), 
	.D(FE_PHN1252_n2792), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][1]  (.Q(\ram[138][1] ), 
	.D(FE_PHN1135_n2791), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[138][0]  (.Q(\ram[138][0] ), 
	.D(FE_PHN2692_n2790), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[134][15]  (.Q(\ram[134][15] ), 
	.D(FE_PHN241_n2741), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[134][14]  (.Q(\ram[134][14] ), 
	.D(FE_PHN5707_n2740), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[134][13]  (.Q(\ram[134][13] ), 
	.D(FE_PHN703_n2739), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[134][12]  (.Q(\ram[134][12] ), 
	.D(FE_PHN1130_n2738), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][11]  (.Q(\ram[134][11] ), 
	.D(FE_PHN1731_n2737), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[134][10]  (.Q(\ram[134][10] ), 
	.D(FE_PHN964_n2736), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][9]  (.Q(\ram[134][9] ), 
	.D(FE_PHN4447_n2735), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[134][8]  (.Q(\ram[134][8] ), 
	.D(FE_PHN2090_n2734), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[134][7]  (.Q(\ram[134][7] ), 
	.D(FE_PHN4759_n2733), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][6]  (.Q(\ram[134][6] ), 
	.D(FE_PHN4757_n2732), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][5]  (.Q(\ram[134][5] ), 
	.D(FE_PHN2072_n2731), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][4]  (.Q(\ram[134][4] ), 
	.D(FE_PHN2191_n2730), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[134][3]  (.Q(\ram[134][3] ), 
	.D(FE_PHN1827_n2729), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][2]  (.Q(\ram[134][2] ), 
	.D(FE_PHN330_n2728), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[134][1]  (.Q(\ram[134][1] ), 
	.D(FE_PHN4756_n2727), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[134][0]  (.Q(\ram[134][0] ), 
	.D(FE_PHN2498_n2726), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[130][15]  (.Q(\ram[130][15] ), 
	.D(FE_PHN1188_n2677), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][14]  (.Q(\ram[130][14] ), 
	.D(FE_PHN1924_n2676), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][13]  (.Q(\ram[130][13] ), 
	.D(FE_PHN2826_n2675), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][12]  (.Q(\ram[130][12] ), 
	.D(FE_PHN2955_n2674), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][11]  (.Q(\ram[130][11] ), 
	.D(FE_PHN676_n2673), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[130][10]  (.Q(\ram[130][10] ), 
	.D(FE_PHN2320_n2672), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[130][9]  (.Q(\ram[130][9] ), 
	.D(FE_PHN2172_n2671), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[130][8]  (.Q(\ram[130][8] ), 
	.D(FE_PHN2656_n2670), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[130][7]  (.Q(\ram[130][7] ), 
	.D(FE_PHN2542_n2669), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[130][6]  (.Q(\ram[130][6] ), 
	.D(FE_PHN1795_n2668), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[130][5]  (.Q(\ram[130][5] ), 
	.D(FE_PHN556_n2667), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[130][4]  (.Q(\ram[130][4] ), 
	.D(FE_PHN1646_n2666), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[130][3]  (.Q(\ram[130][3] ), 
	.D(FE_PHN3018_n2665), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[130][2]  (.Q(\ram[130][2] ), 
	.D(FE_PHN1662_n2664), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[130][1]  (.Q(\ram[130][1] ), 
	.D(FE_PHN2533_n2663), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[130][0]  (.Q(\ram[130][0] ), 
	.D(FE_PHN2300_n2662), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[126][15]  (.Q(\ram[126][15] ), 
	.D(FE_PHN3120_n2613), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][14]  (.Q(\ram[126][14] ), 
	.D(FE_PHN5684_n2612), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][13]  (.Q(\ram[126][13] ), 
	.D(FE_PHN5730_n2611), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][12]  (.Q(\ram[126][12] ), 
	.D(FE_PHN4930_n2610), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][11]  (.Q(\ram[126][11] ), 
	.D(FE_PHN5678_n2609), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][10]  (.Q(\ram[126][10] ), 
	.D(FE_PHN1585_n2608), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][9]  (.Q(\ram[126][9] ), 
	.D(FE_PHN2269_n2607), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[126][8]  (.Q(\ram[126][8] ), 
	.D(FE_PHN2146_n2606), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][7]  (.Q(\ram[126][7] ), 
	.D(FE_PHN4758_n2605), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[126][6]  (.Q(\ram[126][6] ), 
	.D(FE_PHN7213_n2604), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[126][5]  (.Q(\ram[126][5] ), 
	.D(FE_PHN7265_n2603), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[126][4]  (.Q(\ram[126][4] ), 
	.D(FE_PHN5722_n2602), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[126][3]  (.Q(\ram[126][3] ), 
	.D(FE_PHN284_n2601), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[126][2]  (.Q(\ram[126][2] ), 
	.D(FE_PHN4752_n2600), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][1]  (.Q(\ram[126][1] ), 
	.D(FE_PHN4426_n2599), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[126][0]  (.Q(\ram[126][0] ), 
	.D(FE_PHN7039_n2598), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[122][15]  (.Q(\ram[122][15] ), 
	.D(FE_PHN3163_n2549), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][14]  (.Q(\ram[122][14] ), 
	.D(FE_PHN1633_n2548), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][13]  (.Q(\ram[122][13] ), 
	.D(FE_PHN2058_n2547), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[122][12]  (.Q(\ram[122][12] ), 
	.D(FE_PHN2929_n2546), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][11]  (.Q(\ram[122][11] ), 
	.D(FE_PHN2738_n2545), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][10]  (.Q(\ram[122][10] ), 
	.D(FE_PHN2572_n2544), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][9]  (.Q(\ram[122][9] ), 
	.D(FE_PHN2401_n2543), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][8]  (.Q(\ram[122][8] ), 
	.D(FE_PHN2753_n2542), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][7]  (.Q(\ram[122][7] ), 
	.D(FE_PHN2315_n2541), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][6]  (.Q(\ram[122][6] ), 
	.D(FE_PHN297_n2540), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[122][5]  (.Q(\ram[122][5] ), 
	.D(FE_PHN1523_n2539), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[122][4]  (.Q(\ram[122][4] ), 
	.D(FE_PHN1348_n2538), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[122][3]  (.Q(\ram[122][3] ), 
	.D(FE_PHN1377_n2537), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[122][2]  (.Q(\ram[122][2] ), 
	.D(n2536), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[122][1]  (.Q(\ram[122][1] ), 
	.D(FE_PHN2571_n2535), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[122][0]  (.Q(\ram[122][0] ), 
	.D(FE_PHN2480_n2534), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[118][15]  (.Q(\ram[118][15] ), 
	.D(FE_PHN2230_n2485), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[118][14]  (.Q(\ram[118][14] ), 
	.D(FE_PHN881_n2484), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][13]  (.Q(\ram[118][13] ), 
	.D(FE_PHN2475_n2483), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[118][12]  (.Q(\ram[118][12] ), 
	.D(FE_PHN1942_n2482), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[118][11]  (.Q(\ram[118][11] ), 
	.D(FE_PHN1090_n2481), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[118][10]  (.Q(\ram[118][10] ), 
	.D(FE_PHN2923_n2480), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[118][9]  (.Q(\ram[118][9] ), 
	.D(FE_PHN2791_n2479), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][8]  (.Q(\ram[118][8] ), 
	.D(FE_PHN2670_n2478), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][7]  (.Q(\ram[118][7] ), 
	.D(FE_PHN1014_n2477), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][6]  (.Q(\ram[118][6] ), 
	.D(FE_PHN194_n2476), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][5]  (.Q(\ram[118][5] ), 
	.D(FE_PHN2134_n2475), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[118][4]  (.Q(\ram[118][4] ), 
	.D(FE_PHN1039_n2474), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][3]  (.Q(\ram[118][3] ), 
	.D(FE_PHN357_n2473), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][2]  (.Q(\ram[118][2] ), 
	.D(FE_PHN1138_n2472), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[118][1]  (.Q(\ram[118][1] ), 
	.D(FE_PHN2976_n2471), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[118][0]  (.Q(\ram[118][0] ), 
	.D(FE_PHN2743_n2470), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[114][15]  (.Q(\ram[114][15] ), 
	.D(FE_PHN4347_n2421), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[114][14]  (.Q(\ram[114][14] ), 
	.D(FE_PHN4655_n2420), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[114][13]  (.Q(\ram[114][13] ), 
	.D(FE_PHN4343_n2419), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[114][12]  (.Q(\ram[114][12] ), 
	.D(FE_PHN826_n2418), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][11]  (.Q(\ram[114][11] ), 
	.D(FE_PHN4801_n2417), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][10]  (.Q(\ram[114][10] ), 
	.D(FE_PHN1028_n2416), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[114][9]  (.Q(\ram[114][9] ), 
	.D(FE_PHN4205_n2415), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[114][8]  (.Q(\ram[114][8] ), 
	.D(FE_PHN5771_n2414), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][7]  (.Q(\ram[114][7] ), 
	.D(FE_PHN3497_n2413), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[114][6]  (.Q(\ram[114][6] ), 
	.D(FE_PHN5704_n2412), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[114][5]  (.Q(\ram[114][5] ), 
	.D(FE_PHN5649_n2411), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[114][4]  (.Q(\ram[114][4] ), 
	.D(FE_PHN7244_n2410), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[114][3]  (.Q(\ram[114][3] ), 
	.D(FE_PHN264_n2409), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[114][2]  (.Q(\ram[114][2] ), 
	.D(FE_PHN4209_n2408), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[114][1]  (.Q(\ram[114][1] ), 
	.D(FE_PHN5651_n2407), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[114][0]  (.Q(\ram[114][0] ), 
	.D(FE_PHN4947_n2406), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[110][15]  (.Q(\ram[110][15] ), 
	.D(FE_PHN1974_n2357), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[110][14]  (.Q(\ram[110][14] ), 
	.D(FE_PHN421_n2356), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[110][13]  (.Q(\ram[110][13] ), 
	.D(FE_PHN3199_n2355), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[110][12]  (.Q(\ram[110][12] ), 
	.D(FE_PHN531_n2354), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[110][11]  (.Q(\ram[110][11] ), 
	.D(FE_PHN1846_n2353), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[110][10]  (.Q(\ram[110][10] ), 
	.D(FE_PHN883_n2352), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[110][9]  (.Q(\ram[110][9] ), 
	.D(FE_PHN2715_n2351), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[110][8]  (.Q(\ram[110][8] ), 
	.D(FE_PHN2027_n2350), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][7]  (.Q(\ram[110][7] ), 
	.D(FE_PHN476_n2349), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[110][6]  (.Q(\ram[110][6] ), 
	.D(FE_PHN462_n2348), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][5]  (.Q(\ram[110][5] ), 
	.D(FE_PHN1911_n2347), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[110][4]  (.Q(\ram[110][4] ), 
	.D(FE_PHN1612_n2346), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][3]  (.Q(\ram[110][3] ), 
	.D(FE_PHN1686_n2345), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[110][2]  (.Q(\ram[110][2] ), 
	.D(FE_PHN2394_n2344), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][1]  (.Q(\ram[110][1] ), 
	.D(FE_PHN334_n2343), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[110][0]  (.Q(\ram[110][0] ), 
	.D(FE_PHN1253_n2342), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[106][15]  (.Q(\ram[106][15] ), 
	.D(FE_PHN2180_n2293), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][14]  (.Q(\ram[106][14] ), 
	.D(FE_PHN2077_n2292), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[106][13]  (.Q(\ram[106][13] ), 
	.D(FE_PHN2118_n2291), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[106][12]  (.Q(\ram[106][12] ), 
	.D(FE_PHN1862_n2290), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][11]  (.Q(\ram[106][11] ), 
	.D(FE_PHN1539_n2289), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[106][10]  (.Q(\ram[106][10] ), 
	.D(FE_PHN620_n2288), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[106][9]  (.Q(\ram[106][9] ), 
	.D(FE_PHN2057_n2287), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[106][8]  (.Q(\ram[106][8] ), 
	.D(FE_PHN1953_n2286), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][7]  (.Q(\ram[106][7] ), 
	.D(FE_PHN2485_n2285), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[106][6]  (.Q(\ram[106][6] ), 
	.D(FE_PHN593_n2284), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][5]  (.Q(\ram[106][5] ), 
	.D(FE_PHN1243_n2283), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[106][4]  (.Q(\ram[106][4] ), 
	.D(FE_PHN2774_n2282), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[106][3]  (.Q(\ram[106][3] ), 
	.D(FE_PHN2612_n2281), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[106][2]  (.Q(\ram[106][2] ), 
	.D(FE_PHN2515_n2280), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][1]  (.Q(\ram[106][1] ), 
	.D(FE_PHN1755_n2279), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[106][0]  (.Q(\ram[106][0] ), 
	.D(FE_PHN271_n2278), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[102][15]  (.Q(\ram[102][15] ), 
	.D(FE_PHN590_n2229), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][14]  (.Q(\ram[102][14] ), 
	.D(FE_PHN1239_n2228), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][13]  (.Q(\ram[102][13] ), 
	.D(FE_PHN3161_n2227), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[102][12]  (.Q(\ram[102][12] ), 
	.D(FE_PHN1076_n2226), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][11]  (.Q(\ram[102][11] ), 
	.D(FE_PHN1863_n2225), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[102][10]  (.Q(\ram[102][10] ), 
	.D(FE_PHN2590_n2224), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[102][9]  (.Q(\ram[102][9] ), 
	.D(FE_PHN3130_n2223), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][8]  (.Q(\ram[102][8] ), 
	.D(FE_PHN743_n2222), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][7]  (.Q(\ram[102][7] ), 
	.D(FE_PHN887_n2221), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[102][6]  (.Q(\ram[102][6] ), 
	.D(FE_PHN2618_n2220), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][5]  (.Q(\ram[102][5] ), 
	.D(FE_PHN735_n2219), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][4]  (.Q(\ram[102][4] ), 
	.D(FE_PHN1448_n2218), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][3]  (.Q(\ram[102][3] ), 
	.D(FE_PHN2988_n2217), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[102][2]  (.Q(\ram[102][2] ), 
	.D(FE_PHN2113_n2216), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[102][1]  (.Q(\ram[102][1] ), 
	.D(FE_PHN2841_n2215), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[102][0]  (.Q(\ram[102][0] ), 
	.D(FE_PHN3069_n2214), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[98][15]  (.Q(\ram[98][15] ), 
	.D(FE_PHN6682_n2165), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][14]  (.Q(\ram[98][14] ), 
	.D(FE_PHN6689_n2164), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][13]  (.Q(\ram[98][13] ), 
	.D(FE_PHN4319_n2163), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[98][12]  (.Q(\ram[98][12] ), 
	.D(FE_PHN279_n2162), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][11]  (.Q(\ram[98][11] ), 
	.D(FE_PHN5665_n2161), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[98][10]  (.Q(\ram[98][10] ), 
	.D(FE_PHN1282_n2160), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[98][9]  (.Q(\ram[98][9] ), 
	.D(FE_PHN6680_n2159), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][8]  (.Q(\ram[98][8] ), 
	.D(FE_PHN3266_n2158), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][7]  (.Q(\ram[98][7] ), 
	.D(FE_PHN307_n2157), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[98][6]  (.Q(\ram[98][6] ), 
	.D(FE_PHN5703_n2156), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][5]  (.Q(\ram[98][5] ), 
	.D(FE_PHN7232_n2155), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[98][4]  (.Q(\ram[98][4] ), 
	.D(FE_PHN6693_n2154), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[98][3]  (.Q(\ram[98][3] ), 
	.D(n2153), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[98][2]  (.Q(\ram[98][2] ), 
	.D(FE_PHN6641_n2152), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[98][1]  (.Q(\ram[98][1] ), 
	.D(FE_PHN6672_n2151), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[98][0]  (.Q(\ram[98][0] ), 
	.D(FE_PHN786_n2150), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[94][15]  (.Q(\ram[94][15] ), 
	.D(FE_PHN2694_n2101), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][14]  (.Q(\ram[94][14] ), 
	.D(FE_PHN2265_n2100), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][13]  (.Q(\ram[94][13] ), 
	.D(FE_PHN2014_n2099), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][12]  (.Q(\ram[94][12] ), 
	.D(FE_PHN3020_n2098), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][11]  (.Q(\ram[94][11] ), 
	.D(FE_PHN1723_n2097), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][10]  (.Q(\ram[94][10] ), 
	.D(FE_PHN2103_n2096), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][9]  (.Q(\ram[94][9] ), 
	.D(FE_PHN1659_n2095), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][8]  (.Q(\ram[94][8] ), 
	.D(FE_PHN928_n2094), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[94][7]  (.Q(\ram[94][7] ), 
	.D(FE_PHN2865_n2093), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][6]  (.Q(\ram[94][6] ), 
	.D(FE_PHN1542_n2092), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][5]  (.Q(\ram[94][5] ), 
	.D(FE_PHN2228_n2091), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[94][4]  (.Q(\ram[94][4] ), 
	.D(FE_PHN2338_n2090), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][3]  (.Q(\ram[94][3] ), 
	.D(FE_PHN608_n2089), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][2]  (.Q(\ram[94][2] ), 
	.D(FE_PHN1687_n2088), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[94][1]  (.Q(\ram[94][1] ), 
	.D(FE_PHN2373_n2087), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[94][0]  (.Q(\ram[94][0] ), 
	.D(FE_PHN2922_n2086), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[90][15]  (.Q(\ram[90][15] ), 
	.D(FE_PHN2745_n2037), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][14]  (.Q(\ram[90][14] ), 
	.D(FE_PHN2985_n2036), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[90][13]  (.Q(\ram[90][13] ), 
	.D(FE_PHN2619_n2035), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][12]  (.Q(\ram[90][12] ), 
	.D(FE_PHN1745_n2034), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[90][11]  (.Q(\ram[90][11] ), 
	.D(FE_PHN2040_n2033), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[90][10]  (.Q(\ram[90][10] ), 
	.D(FE_PHN410_n2032), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][9]  (.Q(\ram[90][9] ), 
	.D(FE_PHN3012_n2031), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][8]  (.Q(\ram[90][8] ), 
	.D(FE_PHN2973_n2030), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][7]  (.Q(\ram[90][7] ), 
	.D(FE_PHN2354_n2029), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][6]  (.Q(\ram[90][6] ), 
	.D(FE_PHN1784_n2028), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][5]  (.Q(\ram[90][5] ), 
	.D(FE_PHN1053_n2027), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[90][4]  (.Q(\ram[90][4] ), 
	.D(FE_PHN1729_n2026), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][3]  (.Q(\ram[90][3] ), 
	.D(FE_PHN1552_n2025), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[90][2]  (.Q(\ram[90][2] ), 
	.D(FE_PHN2540_n2024), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][1]  (.Q(\ram[90][1] ), 
	.D(FE_PHN2699_n2023), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[90][0]  (.Q(\ram[90][0] ), 
	.D(FE_PHN2409_n2022), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[86][15]  (.Q(\ram[86][15] ), 
	.D(FE_PHN2132_n1973), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][14]  (.Q(\ram[86][14] ), 
	.D(FE_PHN2399_n1972), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][13]  (.Q(\ram[86][13] ), 
	.D(FE_PHN1740_n1971), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][12]  (.Q(\ram[86][12] ), 
	.D(FE_PHN2369_n1970), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[86][11]  (.Q(\ram[86][11] ), 
	.D(FE_PHN3002_n1969), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][10]  (.Q(\ram[86][10] ), 
	.D(FE_PHN2218_n1968), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[86][9]  (.Q(\ram[86][9] ), 
	.D(FE_PHN2020_n1967), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][8]  (.Q(\ram[86][8] ), 
	.D(FE_PHN2002_n1966), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[86][7]  (.Q(\ram[86][7] ), 
	.D(FE_PHN1485_n1965), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][6]  (.Q(\ram[86][6] ), 
	.D(FE_PHN2583_n1964), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][5]  (.Q(\ram[86][5] ), 
	.D(FE_PHN2963_n1963), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][4]  (.Q(\ram[86][4] ), 
	.D(FE_PHN3201_n1962), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][3]  (.Q(\ram[86][3] ), 
	.D(FE_PHN2806_n1961), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][2]  (.Q(\ram[86][2] ), 
	.D(FE_PHN1788_n1960), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[86][1]  (.Q(\ram[86][1] ), 
	.D(FE_PHN2682_n1959), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[86][0]  (.Q(\ram[86][0] ), 
	.D(FE_PHN2500_n1958), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[82][15]  (.Q(\ram[82][15] ), 
	.D(FE_PHN1680_n1909), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][14]  (.Q(\ram[82][14] ), 
	.D(FE_PHN5762_n1908), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][13]  (.Q(\ram[82][13] ), 
	.D(FE_PHN1347_n1907), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][12]  (.Q(\ram[82][12] ), 
	.D(FE_PHN4400_n1906), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][11]  (.Q(\ram[82][11] ), 
	.D(FE_PHN4193_n1905), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[82][10]  (.Q(\ram[82][10] ), 
	.D(FE_PHN3716_n1904), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[82][9]  (.Q(\ram[82][9] ), 
	.D(FE_PHN1235_n1903), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[82][8]  (.Q(\ram[82][8] ), 
	.D(FE_PHN4290_n1902), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][7]  (.Q(\ram[82][7] ), 
	.D(FE_PHN3142_n1901), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[82][6]  (.Q(\ram[82][6] ), 
	.D(FE_PHN1378_n1900), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][5]  (.Q(\ram[82][5] ), 
	.D(FE_PHN4356_n1899), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][4]  (.Q(\ram[82][4] ), 
	.D(FE_PHN2423_n1898), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[82][3]  (.Q(\ram[82][3] ), 
	.D(FE_PHN2972_n1897), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[82][2]  (.Q(\ram[82][2] ), 
	.D(FE_PHN4288_n1896), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[82][1]  (.Q(\ram[82][1] ), 
	.D(FE_PHN1508_n1895), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[82][0]  (.Q(\ram[82][0] ), 
	.D(FE_PHN2499_n1894), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[78][15]  (.Q(\ram[78][15] ), 
	.D(FE_PHN926_n1845), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][14]  (.Q(\ram[78][14] ), 
	.D(FE_PHN1477_n1844), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[78][13]  (.Q(\ram[78][13] ), 
	.D(FE_PHN1025_n1843), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][12]  (.Q(\ram[78][12] ), 
	.D(FE_PHN1780_n1842), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][11]  (.Q(\ram[78][11] ), 
	.D(FE_PHN905_n1841), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][10]  (.Q(\ram[78][10] ), 
	.D(FE_PHN1162_n1840), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][9]  (.Q(\ram[78][9] ), 
	.D(FE_PHN1955_n1839), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[78][8]  (.Q(\ram[78][8] ), 
	.D(n1838), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[78][7]  (.Q(\ram[78][7] ), 
	.D(FE_PHN1416_n1837), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[78][6]  (.Q(\ram[78][6] ), 
	.D(FE_PHN1796_n1836), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][5]  (.Q(\ram[78][5] ), 
	.D(FE_PHN1521_n1835), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][4]  (.Q(\ram[78][4] ), 
	.D(FE_PHN594_n1834), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[78][3]  (.Q(\ram[78][3] ), 
	.D(FE_PHN1387_n1833), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[78][2]  (.Q(\ram[78][2] ), 
	.D(FE_PHN995_n1832), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[78][1]  (.Q(\ram[78][1] ), 
	.D(FE_PHN691_n1831), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[78][0]  (.Q(\ram[78][0] ), 
	.D(FE_PHN1484_n1830), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[74][15]  (.Q(\ram[74][15] ), 
	.D(FE_PHN255_n1781), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][14]  (.Q(\ram[74][14] ), 
	.D(FE_PHN3188_n1780), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][13]  (.Q(\ram[74][13] ), 
	.D(FE_PHN2910_n1779), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[74][12]  (.Q(\ram[74][12] ), 
	.D(FE_PHN2395_n1778), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][11]  (.Q(\ram[74][11] ), 
	.D(FE_PHN865_n1777), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][10]  (.Q(\ram[74][10] ), 
	.D(FE_PHN2482_n1776), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][9]  (.Q(\ram[74][9] ), 
	.D(FE_PHN2128_n1775), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[74][8]  (.Q(\ram[74][8] ), 
	.D(FE_PHN2677_n1774), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[74][7]  (.Q(\ram[74][7] ), 
	.D(FE_PHN3228_n1773), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][6]  (.Q(\ram[74][6] ), 
	.D(FE_PHN3154_n1772), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][5]  (.Q(\ram[74][5] ), 
	.D(FE_PHN681_n1771), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][4]  (.Q(\ram[74][4] ), 
	.D(FE_PHN388_n1770), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[74][3]  (.Q(\ram[74][3] ), 
	.D(FE_PHN1313_n1769), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[74][2]  (.Q(\ram[74][2] ), 
	.D(FE_PHN2060_n1768), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[74][1]  (.Q(\ram[74][1] ), 
	.D(FE_PHN2609_n1767), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[74][0]  (.Q(\ram[74][0] ), 
	.D(FE_PHN2012_n1766), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[70][15]  (.Q(\ram[70][15] ), 
	.D(FE_PHN1668_n1717), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][14]  (.Q(\ram[70][14] ), 
	.D(FE_PHN728_n1716), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][13]  (.Q(\ram[70][13] ), 
	.D(FE_PHN895_n1715), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][12]  (.Q(\ram[70][12] ), 
	.D(FE_PHN3117_n1714), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][11]  (.Q(\ram[70][11] ), 
	.D(FE_PHN138_n1713), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][10]  (.Q(\ram[70][10] ), 
	.D(FE_PHN2162_n1712), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][9]  (.Q(\ram[70][9] ), 
	.D(FE_PHN362_n1711), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[70][8]  (.Q(\ram[70][8] ), 
	.D(FE_PHN422_n1710), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][7]  (.Q(\ram[70][7] ), 
	.D(FE_PHN1538_n1709), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][6]  (.Q(\ram[70][6] ), 
	.D(FE_PHN378_n1708), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][5]  (.Q(\ram[70][5] ), 
	.D(FE_PHN380_n1707), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][4]  (.Q(\ram[70][4] ), 
	.D(FE_PHN2201_n1706), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[70][3]  (.Q(\ram[70][3] ), 
	.D(FE_PHN2991_n1705), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[70][2]  (.Q(\ram[70][2] ), 
	.D(FE_PHN143_n1704), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[70][1]  (.Q(\ram[70][1] ), 
	.D(FE_PHN719_n1703), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[70][0]  (.Q(\ram[70][0] ), 
	.D(FE_PHN591_n1702), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[66][15]  (.Q(\ram[66][15] ), 
	.D(FE_PHN356_n1653), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][14]  (.Q(\ram[66][14] ), 
	.D(FE_PHN3077_n1652), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][13]  (.Q(\ram[66][13] ), 
	.D(FE_PHN1251_n1651), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[66][12]  (.Q(\ram[66][12] ), 
	.D(FE_PHN802_n1650), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[66][11]  (.Q(\ram[66][11] ), 
	.D(FE_PHN1839_n1649), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][10]  (.Q(\ram[66][10] ), 
	.D(FE_PHN1979_n1648), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[66][9]  (.Q(\ram[66][9] ), 
	.D(FE_PHN683_n1647), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[66][8]  (.Q(\ram[66][8] ), 
	.D(FE_PHN2069_n1646), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][7]  (.Q(\ram[66][7] ), 
	.D(FE_PHN968_n1645), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][6]  (.Q(\ram[66][6] ), 
	.D(FE_PHN429_n1644), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][5]  (.Q(\ram[66][5] ), 
	.D(FE_PHN1304_n1643), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][4]  (.Q(\ram[66][4] ), 
	.D(FE_PHN2981_n1642), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][3]  (.Q(\ram[66][3] ), 
	.D(FE_PHN1882_n1641), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][2]  (.Q(\ram[66][2] ), 
	.D(FE_PHN653_n1640), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[66][1]  (.Q(\ram[66][1] ), 
	.D(FE_PHN2158_n1639), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[66][0]  (.Q(\ram[66][0] ), 
	.D(FE_PHN2261_n1638), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[62][15]  (.Q(\ram[62][15] ), 
	.D(FE_PHN2486_n1589), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][14]  (.Q(\ram[62][14] ), 
	.D(FE_PHN1142_n1588), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][13]  (.Q(\ram[62][13] ), 
	.D(FE_PHN2350_n1587), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][12]  (.Q(\ram[62][12] ), 
	.D(FE_PHN1990_n1586), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[62][11]  (.Q(\ram[62][11] ), 
	.D(FE_PHN2181_n1585), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][10]  (.Q(\ram[62][10] ), 
	.D(FE_PHN2685_n1584), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][9]  (.Q(\ram[62][9] ), 
	.D(FE_PHN2110_n1583), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[62][8]  (.Q(\ram[62][8] ), 
	.D(FE_PHN1925_n1582), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][7]  (.Q(\ram[62][7] ), 
	.D(FE_PHN1137_n1581), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[62][6]  (.Q(\ram[62][6] ), 
	.D(FE_PHN2752_n1580), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][5]  (.Q(\ram[62][5] ), 
	.D(FE_PHN3017_n1579), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][4]  (.Q(\ram[62][4] ), 
	.D(FE_PHN2733_n1578), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[62][3]  (.Q(\ram[62][3] ), 
	.D(FE_PHN527_n1577), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[62][2]  (.Q(\ram[62][2] ), 
	.D(FE_PHN2693_n1576), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[62][1]  (.Q(\ram[62][1] ), 
	.D(FE_PHN1408_n1575), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[62][0]  (.Q(\ram[62][0] ), 
	.D(FE_PHN3045_n1574), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[58][15]  (.Q(\ram[58][15] ), 
	.D(FE_PHN404_n1525), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[58][14]  (.Q(\ram[58][14] ), 
	.D(FE_PHN808_n1524), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[58][13]  (.Q(\ram[58][13] ), 
	.D(FE_PHN923_n1523), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[58][12]  (.Q(\ram[58][12] ), 
	.D(FE_PHN1070_n1522), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][11]  (.Q(\ram[58][11] ), 
	.D(FE_PHN1637_n1521), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][10]  (.Q(\ram[58][10] ), 
	.D(FE_PHN2283_n1520), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[58][9]  (.Q(\ram[58][9] ), 
	.D(FE_PHN2666_n1519), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][8]  (.Q(\ram[58][8] ), 
	.D(FE_PHN2691_n1518), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[58][7]  (.Q(\ram[58][7] ), 
	.D(FE_PHN2249_n1517), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][6]  (.Q(\ram[58][6] ), 
	.D(FE_PHN1853_n1516), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][5]  (.Q(\ram[58][5] ), 
	.D(FE_PHN1357_n1515), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[58][4]  (.Q(\ram[58][4] ), 
	.D(FE_PHN2161_n1514), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][3]  (.Q(\ram[58][3] ), 
	.D(FE_PHN2522_n1513), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[58][2]  (.Q(\ram[58][2] ), 
	.D(FE_PHN2295_n1512), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][1]  (.Q(\ram[58][1] ), 
	.D(FE_PHN3191_n1511), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[58][0]  (.Q(\ram[58][0] ), 
	.D(FE_PHN1352_n1510), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[54][15]  (.Q(\ram[54][15] ), 
	.D(FE_PHN3076_n1461), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][14]  (.Q(\ram[54][14] ), 
	.D(FE_PHN2586_n1460), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[54][13]  (.Q(\ram[54][13] ), 
	.D(FE_PHN1724_n1459), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[54][12]  (.Q(\ram[54][12] ), 
	.D(FE_PHN2594_n1458), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][11]  (.Q(\ram[54][11] ), 
	.D(FE_PHN2843_n1457), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][10]  (.Q(\ram[54][10] ), 
	.D(FE_PHN2637_n1456), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][9]  (.Q(\ram[54][9] ), 
	.D(FE_PHN2928_n1455), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][8]  (.Q(\ram[54][8] ), 
	.D(FE_PHN2953_n1454), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][7]  (.Q(\ram[54][7] ), 
	.D(FE_PHN2372_n1453), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][6]  (.Q(\ram[54][6] ), 
	.D(FE_PHN3113_n1452), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][5]  (.Q(\ram[54][5] ), 
	.D(FE_PHN3005_n1451), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][4]  (.Q(\ram[54][4] ), 
	.D(FE_PHN956_n1450), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][3]  (.Q(\ram[54][3] ), 
	.D(FE_PHN3159_n1449), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[54][2]  (.Q(\ram[54][2] ), 
	.D(FE_PHN2997_n1448), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][1]  (.Q(\ram[54][1] ), 
	.D(FE_PHN2773_n1447), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[54][0]  (.Q(\ram[54][0] ), 
	.D(FE_PHN938_n1446), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[50][15]  (.Q(\ram[50][15] ), 
	.D(FE_PHN2190_n1397), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[50][14]  (.Q(\ram[50][14] ), 
	.D(FE_PHN1983_n1396), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[50][13]  (.Q(\ram[50][13] ), 
	.D(FE_PHN2882_n1395), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[50][12]  (.Q(\ram[50][12] ), 
	.D(FE_PHN1270_n1394), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][11]  (.Q(\ram[50][11] ), 
	.D(FE_PHN1966_n1393), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][10]  (.Q(\ram[50][10] ), 
	.D(FE_PHN397_n1392), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][9]  (.Q(\ram[50][9] ), 
	.D(FE_PHN2114_n1391), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[50][8]  (.Q(\ram[50][8] ), 
	.D(FE_PHN1713_n1390), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[50][7]  (.Q(\ram[50][7] ), 
	.D(FE_PHN2517_n1389), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[50][6]  (.Q(\ram[50][6] ), 
	.D(FE_PHN1878_n1388), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[50][5]  (.Q(\ram[50][5] ), 
	.D(FE_PHN1117_n1387), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][4]  (.Q(\ram[50][4] ), 
	.D(FE_PHN1101_n1386), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[50][3]  (.Q(\ram[50][3] ), 
	.D(FE_PHN1196_n1385), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[50][2]  (.Q(\ram[50][2] ), 
	.D(FE_PHN1019_n1384), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[50][1]  (.Q(\ram[50][1] ), 
	.D(FE_PHN2508_n1383), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[50][0]  (.Q(\ram[50][0] ), 
	.D(FE_PHN3182_n1382), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[46][15]  (.Q(\ram[46][15] ), 
	.D(FE_PHN1850_n1333), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[46][14]  (.Q(\ram[46][14] ), 
	.D(FE_PHN1461_n1332), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][13]  (.Q(\ram[46][13] ), 
	.D(FE_PHN2763_n1331), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[46][12]  (.Q(\ram[46][12] ), 
	.D(FE_PHN360_n1330), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[46][11]  (.Q(\ram[46][11] ), 
	.D(FE_PHN967_n1329), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][10]  (.Q(\ram[46][10] ), 
	.D(FE_PHN3194_n1328), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[46][9]  (.Q(\ram[46][9] ), 
	.D(FE_PHN1401_n1327), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[46][8]  (.Q(\ram[46][8] ), 
	.D(FE_PHN2345_n1326), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[46][7]  (.Q(\ram[46][7] ), 
	.D(FE_PHN2950_n1325), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[46][6]  (.Q(\ram[46][6] ), 
	.D(FE_PHN3198_n1324), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][5]  (.Q(\ram[46][5] ), 
	.D(FE_PHN2164_n1323), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][4]  (.Q(\ram[46][4] ), 
	.D(FE_PHN2491_n1322), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][3]  (.Q(\ram[46][3] ), 
	.D(FE_PHN1792_n1321), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[46][2]  (.Q(\ram[46][2] ), 
	.D(n1320), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][1]  (.Q(\ram[46][1] ), 
	.D(FE_PHN2004_n1319), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[46][0]  (.Q(\ram[46][0] ), 
	.D(FE_PHN2342_n1318), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[42][15]  (.Q(\ram[42][15] ), 
	.D(FE_PHN3138_n1269), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[42][14]  (.Q(\ram[42][14] ), 
	.D(FE_PHN2765_n1268), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][13]  (.Q(\ram[42][13] ), 
	.D(FE_PHN2418_n1267), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][12]  (.Q(\ram[42][12] ), 
	.D(FE_PHN2905_n1266), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[42][11]  (.Q(\ram[42][11] ), 
	.D(FE_PHN2139_n1265), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][10]  (.Q(\ram[42][10] ), 
	.D(FE_PHN2786_n1264), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[42][9]  (.Q(\ram[42][9] ), 
	.D(FE_PHN2610_n1263), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[42][8]  (.Q(\ram[42][8] ), 
	.D(FE_PHN2250_n1262), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][7]  (.Q(\ram[42][7] ), 
	.D(FE_PHN1932_n1261), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[42][6]  (.Q(\ram[42][6] ), 
	.D(FE_PHN1071_n1260), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][5]  (.Q(\ram[42][5] ), 
	.D(FE_PHN3032_n1259), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][4]  (.Q(\ram[42][4] ), 
	.D(FE_PHN1894_n1258), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][3]  (.Q(\ram[42][3] ), 
	.D(FE_PHN2388_n1257), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[42][2]  (.Q(\ram[42][2] ), 
	.D(FE_PHN2336_n1256), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[42][1]  (.Q(\ram[42][1] ), 
	.D(FE_PHN803_n1255), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[42][0]  (.Q(\ram[42][0] ), 
	.D(FE_PHN3148_n1254), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[38][15]  (.Q(\ram[38][15] ), 
	.D(FE_PHN2900_n1205), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][14]  (.Q(\ram[38][14] ), 
	.D(FE_PHN1578_n1204), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][13]  (.Q(\ram[38][13] ), 
	.D(FE_PHN3129_n1203), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][12]  (.Q(\ram[38][12] ), 
	.D(FE_PHN1365_n1202), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[38][11]  (.Q(\ram[38][11] ), 
	.D(FE_PHN2256_n1201), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[38][10]  (.Q(\ram[38][10] ), 
	.D(FE_PHN2718_n1200), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[38][9]  (.Q(\ram[38][9] ), 
	.D(FE_PHN2157_n1199), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][8]  (.Q(\ram[38][8] ), 
	.D(FE_PHN2509_n1198), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[38][7]  (.Q(\ram[38][7] ), 
	.D(FE_PHN3223_n1197), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[38][6]  (.Q(\ram[38][6] ), 
	.D(FE_PHN1148_n1196), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[38][5]  (.Q(\ram[38][5] ), 
	.D(FE_PHN2431_n1195), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[38][4]  (.Q(\ram[38][4] ), 
	.D(FE_PHN377_n1194), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[38][3]  (.Q(\ram[38][3] ), 
	.D(FE_PHN2165_n1193), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[38][2]  (.Q(\ram[38][2] ), 
	.D(FE_PHN1207_n1192), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[38][1]  (.Q(\ram[38][1] ), 
	.D(FE_PHN857_n1191), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[38][0]  (.Q(\ram[38][0] ), 
	.D(FE_PHN5676_n1190), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[34][15]  (.Q(\ram[34][15] ), 
	.D(FE_PHN1948_n1141), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][14]  (.Q(\ram[34][14] ), 
	.D(FE_PHN1254_n1140), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][13]  (.Q(\ram[34][13] ), 
	.D(FE_PHN1879_n1139), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][12]  (.Q(\ram[34][12] ), 
	.D(FE_PHN1424_n1138), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[34][11]  (.Q(\ram[34][11] ), 
	.D(FE_PHN457_n1137), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][10]  (.Q(\ram[34][10] ), 
	.D(FE_PHN1959_n1136), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[34][9]  (.Q(\ram[34][9] ), 
	.D(FE_PHN2589_n1135), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][8]  (.Q(\ram[34][8] ), 
	.D(FE_PHN3060_n1134), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[34][7]  (.Q(\ram[34][7] ), 
	.D(FE_PHN2889_n1133), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[34][6]  (.Q(\ram[34][6] ), 
	.D(FE_PHN3215_n1132), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][5]  (.Q(\ram[34][5] ), 
	.D(FE_PHN1601_n1131), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][4]  (.Q(\ram[34][4] ), 
	.D(FE_PHN1084_n1130), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[34][3]  (.Q(\ram[34][3] ), 
	.D(FE_PHN1650_n1129), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[34][2]  (.Q(\ram[34][2] ), 
	.D(FE_PHN870_n1128), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[34][1]  (.Q(\ram[34][1] ), 
	.D(FE_PHN2729_n1127), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[34][0]  (.Q(\ram[34][0] ), 
	.D(FE_PHN959_n1126), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[30][15]  (.Q(\ram[30][15] ), 
	.D(FE_PHN4212_n1077), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[30][14]  (.Q(\ram[30][14] ), 
	.D(FE_PHN523_n1076), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][13]  (.Q(\ram[30][13] ), 
	.D(FE_PHN1308_n1075), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[30][12]  (.Q(\ram[30][12] ), 
	.D(FE_PHN4397_n1074), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[30][11]  (.Q(\ram[30][11] ), 
	.D(FE_PHN1332_n1073), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][10]  (.Q(\ram[30][10] ), 
	.D(FE_PHN4230_n1072), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[30][9]  (.Q(\ram[30][9] ), 
	.D(FE_PHN1469_n1071), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][8]  (.Q(\ram[30][8] ), 
	.D(FE_PHN2496_n1070), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][7]  (.Q(\ram[30][7] ), 
	.D(FE_PHN4289_n1069), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][6]  (.Q(\ram[30][6] ), 
	.D(FE_PHN3685_n1068), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][5]  (.Q(\ram[30][5] ), 
	.D(FE_PHN1418_n1067), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][4]  (.Q(\ram[30][4] ), 
	.D(FE_PHN4705_n1066), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[30][3]  (.Q(\ram[30][3] ), 
	.D(FE_PHN361_n1065), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[30][2]  (.Q(\ram[30][2] ), 
	.D(FE_PHN4282_n1064), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[30][1]  (.Q(\ram[30][1] ), 
	.D(FE_PHN352_n1063), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[30][0]  (.Q(\ram[30][0] ), 
	.D(FE_PHN3330_n1062), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[26][15]  (.Q(\ram[26][15] ), 
	.D(FE_PHN3269_n1013), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][14]  (.Q(\ram[26][14] ), 
	.D(FE_PHN5750_n1012), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][13]  (.Q(\ram[26][13] ), 
	.D(FE_PHN1834_n1011), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][12]  (.Q(\ram[26][12] ), 
	.D(FE_PHN311_n1010), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][11]  (.Q(\ram[26][11] ), 
	.D(FE_PHN5094_n1009), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][10]  (.Q(\ram[26][10] ), 
	.D(FE_PHN4131_n1008), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][9]  (.Q(\ram[26][9] ), 
	.D(FE_PHN4891_n1007), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][8]  (.Q(\ram[26][8] ), 
	.D(FE_PHN3875_n1006), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][7]  (.Q(\ram[26][7] ), 
	.D(FE_PHN5441_n1005), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][6]  (.Q(\ram[26][6] ), 
	.D(FE_PHN832_n1004), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][5]  (.Q(\ram[26][5] ), 
	.D(FE_PHN5746_n1003), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][4]  (.Q(\ram[26][4] ), 
	.D(FE_PHN4394_n1002), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[26][3]  (.Q(\ram[26][3] ), 
	.D(FE_PHN4882_n1001), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[26][2]  (.Q(\ram[26][2] ), 
	.D(FE_PHN4455_n1000), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[26][1]  (.Q(\ram[26][1] ), 
	.D(FE_PHN4517_n999), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[26][0]  (.Q(\ram[26][0] ), 
	.D(FE_PHN3569_n998), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[22][15]  (.Q(\ram[22][15] ), 
	.D(FE_PHN4354_n949), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][14]  (.Q(\ram[22][14] ), 
	.D(FE_PHN4581_n948), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][13]  (.Q(\ram[22][13] ), 
	.D(FE_PHN4242_n947), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[22][12]  (.Q(\ram[22][12] ), 
	.D(FE_PHN5095_n946), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[22][11]  (.Q(\ram[22][11] ), 
	.D(FE_PHN4228_n945), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][10]  (.Q(\ram[22][10] ), 
	.D(FE_PHN4474_n944), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[22][9]  (.Q(\ram[22][9] ), 
	.D(FE_PHN4168_n943), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][8]  (.Q(\ram[22][8] ), 
	.D(FE_PHN933_n942), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][7]  (.Q(\ram[22][7] ), 
	.D(FE_PHN4470_n941), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][6]  (.Q(\ram[22][6] ), 
	.D(FE_PHN2313_n940), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[22][5]  (.Q(\ram[22][5] ), 
	.D(FE_PHN2531_n939), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[22][4]  (.Q(\ram[22][4] ), 
	.D(FE_PHN3535_n938), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][3]  (.Q(\ram[22][3] ), 
	.D(FE_PHN2719_n937), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[22][2]  (.Q(\ram[22][2] ), 
	.D(FE_PHN5186_n936), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[22][1]  (.Q(\ram[22][1] ), 
	.D(FE_PHN4611_n935), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[22][0]  (.Q(\ram[22][0] ), 
	.D(FE_PHN5537_n934), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[18][15]  (.Q(\ram[18][15] ), 
	.D(FE_PHN4393_n885), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[18][14]  (.Q(\ram[18][14] ), 
	.D(FE_PHN4165_n884), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][13]  (.Q(\ram[18][13] ), 
	.D(FE_PHN1874_n883), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[18][12]  (.Q(\ram[18][12] ), 
	.D(FE_PHN4575_n882), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][11]  (.Q(\ram[18][11] ), 
	.D(FE_PHN4457_n881), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[18][10]  (.Q(\ram[18][10] ), 
	.D(FE_PHN4688_n880), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][9]  (.Q(\ram[18][9] ), 
	.D(FE_PHN3305_n879), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[18][8]  (.Q(\ram[18][8] ), 
	.D(FE_PHN4592_n878), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][7]  (.Q(\ram[18][7] ), 
	.D(FE_PHN4601_n877), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[18][6]  (.Q(\ram[18][6] ), 
	.D(FE_PHN5293_n876), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][5]  (.Q(\ram[18][5] ), 
	.D(FE_PHN839_n875), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[18][4]  (.Q(\ram[18][4] ), 
	.D(FE_PHN4673_n874), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][3]  (.Q(\ram[18][3] ), 
	.D(FE_PHN4734_n873), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[18][2]  (.Q(\ram[18][2] ), 
	.D(FE_PHN4249_n872), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[18][1]  (.Q(\ram[18][1] ), 
	.D(FE_PHN5570_n871), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[18][0]  (.Q(\ram[18][0] ), 
	.D(FE_PHN4504_n870), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[14][15]  (.Q(\ram[14][15] ), 
	.D(FE_PHN1681_n821), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][14]  (.Q(\ram[14][14] ), 
	.D(FE_PHN696_n820), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][13]  (.Q(\ram[14][13] ), 
	.D(FE_PHN2750_n819), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][12]  (.Q(\ram[14][12] ), 
	.D(FE_PHN877_n818), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[14][11]  (.Q(\ram[14][11] ), 
	.D(FE_PHN1881_n817), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[14][10]  (.Q(\ram[14][10] ), 
	.D(FE_PHN1506_n816), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[14][9]  (.Q(\ram[14][9] ), 
	.D(FE_PHN2024_n815), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[14][8]  (.Q(\ram[14][8] ), 
	.D(FE_PHN2730_n814), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][7]  (.Q(\ram[14][7] ), 
	.D(FE_PHN934_n813), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][6]  (.Q(\ram[14][6] ), 
	.D(FE_PHN3152_n812), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][5]  (.Q(\ram[14][5] ), 
	.D(FE_PHN3066_n811), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[14][4]  (.Q(\ram[14][4] ), 
	.D(FE_PHN1264_n810), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][3]  (.Q(\ram[14][3] ), 
	.D(FE_PHN3225_n809), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[14][2]  (.Q(\ram[14][2] ), 
	.D(FE_PHN1907_n808), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[14][1]  (.Q(\ram[14][1] ), 
	.D(FE_PHN1801_n807), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[14][0]  (.Q(\ram[14][0] ), 
	.D(FE_PHN623_n806), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[10][15]  (.Q(\ram[10][15] ), 
	.D(FE_PHN1709_n757), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][14]  (.Q(\ram[10][14] ), 
	.D(FE_PHN2633_n756), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[10][13]  (.Q(\ram[10][13] ), 
	.D(FE_PHN2815_n755), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[10][12]  (.Q(\ram[10][12] ), 
	.D(FE_PHN2845_n754), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[10][11]  (.Q(\ram[10][11] ), 
	.D(FE_PHN564_n753), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[10][10]  (.Q(\ram[10][10] ), 
	.D(FE_PHN2229_n752), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][9]  (.Q(\ram[10][9] ), 
	.D(FE_PHN804_n751), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[10][8]  (.Q(\ram[10][8] ), 
	.D(FE_PHN745_n750), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][7]  (.Q(\ram[10][7] ), 
	.D(FE_PHN3189_n749), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][6]  (.Q(\ram[10][6] ), 
	.D(FE_PHN1598_n748), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][5]  (.Q(\ram[10][5] ), 
	.D(FE_PHN2225_n747), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[10][4]  (.Q(\ram[10][4] ), 
	.D(FE_PHN2962_n746), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[10][3]  (.Q(\ram[10][3] ), 
	.D(FE_PHN2149_n745), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[10][2]  (.Q(\ram[10][2] ), 
	.D(FE_PHN2260_n744), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[10][1]  (.Q(\ram[10][1] ), 
	.D(FE_PHN495_n743), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[10][0]  (.Q(\ram[10][0] ), 
	.D(FE_PHN2615_n742), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[6][15]  (.Q(\ram[6][15] ), 
	.D(FE_PHN1693_n693), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][14]  (.Q(\ram[6][14] ), 
	.D(FE_PHN2453_n692), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][13]  (.Q(\ram[6][13] ), 
	.D(FE_PHN2914_n691), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[6][12]  (.Q(\ram[6][12] ), 
	.D(FE_PHN1804_n690), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[6][11]  (.Q(\ram[6][11] ), 
	.D(FE_PHN1059_n689), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[6][10]  (.Q(\ram[6][10] ), 
	.D(FE_PHN3135_n688), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][9]  (.Q(\ram[6][9] ), 
	.D(FE_PHN2564_n687), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[6][8]  (.Q(\ram[6][8] ), 
	.D(FE_PHN2214_n686), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][7]  (.Q(\ram[6][7] ), 
	.D(FE_PHN2312_n685), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][6]  (.Q(\ram[6][6] ), 
	.D(FE_PHN2860_n684), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[6][5]  (.Q(\ram[6][5] ), 
	.D(FE_PHN1223_n683), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[6][4]  (.Q(\ram[6][4] ), 
	.D(FE_PHN1922_n682), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][3]  (.Q(\ram[6][3] ), 
	.D(FE_PHN2724_n681), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[6][2]  (.Q(\ram[6][2] ), 
	.D(FE_PHN2078_n680), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[6][1]  (.Q(\ram[6][1] ), 
	.D(FE_PHN1317_n679), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[6][0]  (.Q(\ram[6][0] ), 
	.D(FE_PHN1639_n678), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[2][15]  (.Q(\ram[2][15] ), 
	.D(FE_PHN2811_n629), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[2][14]  (.Q(\ram[2][14] ), 
	.D(FE_PHN2112_n628), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][13]  (.Q(\ram[2][13] ), 
	.D(FE_PHN2511_n627), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[2][12]  (.Q(\ram[2][12] ), 
	.D(FE_PHN1498_n626), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][11]  (.Q(\ram[2][11] ), 
	.D(FE_PHN3218_n625), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[2][10]  (.Q(\ram[2][10] ), 
	.D(FE_PHN1398_n624), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[2][9]  (.Q(\ram[2][9] ), 
	.D(FE_PHN2829_n623), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[2][8]  (.Q(\ram[2][8] ), 
	.D(FE_PHN2596_n622), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[2][7]  (.Q(\ram[2][7] ), 
	.D(FE_PHN2048_n621), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[2][6]  (.Q(\ram[2][6] ), 
	.D(FE_PHN3061_n620), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[2][5]  (.Q(\ram[2][5] ), 
	.D(FE_PHN775_n619), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[2][4]  (.Q(\ram[2][4] ), 
	.D(FE_PHN1051_n618), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][3]  (.Q(\ram[2][3] ), 
	.D(FE_PHN1008_n617), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[2][2]  (.Q(\ram[2][2] ), 
	.D(FE_PHN3011_n616), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][1]  (.Q(\ram[2][1] ), 
	.D(FE_PHN1045_n615), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[2][0]  (.Q(\ram[2][0] ), 
	.D(FE_PHN1455_n614), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[252][15]  (.Q(\ram[252][15] ), 
	.D(FE_PHN2355_n4629), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[252][14]  (.Q(\ram[252][14] ), 
	.D(FE_PHN2018_n4628), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[252][13]  (.Q(\ram[252][13] ), 
	.D(FE_PHN1281_n4627), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][12]  (.Q(\ram[252][12] ), 
	.D(FE_PHN1323_n4626), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[252][11]  (.Q(\ram[252][11] ), 
	.D(FE_PHN900_n4625), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[252][10]  (.Q(\ram[252][10] ), 
	.D(FE_PHN947_n4624), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][9]  (.Q(\ram[252][9] ), 
	.D(FE_PHN587_n4623), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][8]  (.Q(\ram[252][8] ), 
	.D(FE_PHN537_n4622), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[252][7]  (.Q(\ram[252][7] ), 
	.D(FE_PHN2216_n4621), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[252][6]  (.Q(\ram[252][6] ), 
	.D(FE_PHN2317_n4620), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[252][5]  (.Q(\ram[252][5] ), 
	.D(FE_PHN1840_n4619), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[252][4]  (.Q(\ram[252][4] ), 
	.D(FE_PHN633_n4618), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[252][3]  (.Q(\ram[252][3] ), 
	.D(FE_PHN1184_n4617), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[252][2]  (.Q(\ram[252][2] ), 
	.D(FE_PHN999_n4616), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[252][1]  (.Q(\ram[252][1] ), 
	.D(FE_PHN2432_n4615), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[252][0]  (.Q(\ram[252][0] ), 
	.D(FE_PHN2411_n4614), 
	.CK(clk));
   QDFFEHD \ram_reg[248][15]  (.Q(\ram[248][15] ), 
	.D(FE_PHN448_n4565), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][14]  (.Q(\ram[248][14] ), 
	.D(FE_PHN1761_n4564), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][13]  (.Q(\ram[248][13] ), 
	.D(FE_PHN1694_n4563), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][12]  (.Q(\ram[248][12] ), 
	.D(FE_PHN2021_n4562), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[248][11]  (.Q(\ram[248][11] ), 
	.D(FE_PHN2544_n4561), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][10]  (.Q(\ram[248][10] ), 
	.D(FE_PHN2558_n4560), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][9]  (.Q(\ram[248][9] ), 
	.D(FE_PHN1915_n4559), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][8]  (.Q(\ram[248][8] ), 
	.D(FE_PHN2042_n4558), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[248][7]  (.Q(\ram[248][7] ), 
	.D(FE_PHN3124_n4557), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][6]  (.Q(\ram[248][6] ), 
	.D(FE_PHN1278_n4556), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][5]  (.Q(\ram[248][5] ), 
	.D(FE_PHN784_n4555), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[248][4]  (.Q(\ram[248][4] ), 
	.D(FE_PHN771_n4554), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[248][3]  (.Q(\ram[248][3] ), 
	.D(FE_PHN542_n4553), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[248][2]  (.Q(\ram[248][2] ), 
	.D(FE_PHN1334_n4552), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[248][1]  (.Q(\ram[248][1] ), 
	.D(FE_PHN1865_n4551), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[248][0]  (.Q(\ram[248][0] ), 
	.D(FE_PHN1209_n4550), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][15]  (.Q(\ram[244][15] ), 
	.D(FE_PHN721_n4501), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][14]  (.Q(\ram[244][14] ), 
	.D(FE_PHN1456_n4500), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[244][13]  (.Q(\ram[244][13] ), 
	.D(FE_PHN1036_n4499), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][12]  (.Q(\ram[244][12] ), 
	.D(FE_PHN889_n4498), 
	.CK(clk));
   QDFFEHD \ram_reg[244][11]  (.Q(\ram[244][11] ), 
	.D(FE_PHN2946_n4497), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][10]  (.Q(\ram[244][10] ), 
	.D(n4496), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][9]  (.Q(\ram[244][9] ), 
	.D(FE_PHN700_n4495), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[244][8]  (.Q(\ram[244][8] ), 
	.D(FE_PHN371_n4494), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[244][7]  (.Q(\ram[244][7] ), 
	.D(FE_PHN455_n4493), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[244][6]  (.Q(\ram[244][6] ), 
	.D(FE_PHN1627_n4492), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][5]  (.Q(\ram[244][5] ), 
	.D(FE_PHN1809_n4491), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][4]  (.Q(\ram[244][4] ), 
	.D(FE_PHN1896_n4490), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][3]  (.Q(\ram[244][3] ), 
	.D(FE_PHN1958_n4489), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[244][2]  (.Q(\ram[244][2] ), 
	.D(FE_PHN1434_n4488), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[244][1]  (.Q(\ram[244][1] ), 
	.D(FE_PHN1634_n4487), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[244][0]  (.Q(\ram[244][0] ), 
	.D(FE_PHN996_n4486), 
	.CK(clk));
   QDFFEHD \ram_reg[240][15]  (.Q(\ram[240][15] ), 
	.D(FE_PHN2464_n4437), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[240][14]  (.Q(\ram[240][14] ), 
	.D(FE_PHN685_n4436), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][13]  (.Q(\ram[240][13] ), 
	.D(FE_PHN494_n4435), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][12]  (.Q(\ram[240][12] ), 
	.D(FE_PHN679_n4434), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[240][11]  (.Q(\ram[240][11] ), 
	.D(FE_PHN1375_n4433), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[240][10]  (.Q(\ram[240][10] ), 
	.D(FE_PHN1353_n4432), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][9]  (.Q(\ram[240][9] ), 
	.D(FE_PHN1376_n4431), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[240][8]  (.Q(\ram[240][8] ), 
	.D(FE_PHN2839_n4430), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][7]  (.Q(\ram[240][7] ), 
	.D(FE_PHN1029_n4429), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[240][6]  (.Q(\ram[240][6] ), 
	.D(FE_PHN2695_n4428), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][5]  (.Q(\ram[240][5] ), 
	.D(FE_PHN1057_n4427), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[240][4]  (.Q(\ram[240][4] ), 
	.D(FE_PHN212_n4426), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][3]  (.Q(\ram[240][3] ), 
	.D(FE_PHN766_n4425), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][2]  (.Q(\ram[240][2] ), 
	.D(FE_PHN789_n4424), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][1]  (.Q(\ram[240][1] ), 
	.D(FE_PHN2623_n4423), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[240][0]  (.Q(\ram[240][0] ), 
	.D(FE_PHN890_n4422), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[236][15]  (.Q(\ram[236][15] ), 
	.D(FE_PHN4499_n4373), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][14]  (.Q(\ram[236][14] ), 
	.D(FE_PHN4048_n4372), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[236][13]  (.Q(\ram[236][13] ), 
	.D(FE_PHN4099_n4371), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][12]  (.Q(\ram[236][12] ), 
	.D(FE_PHN4410_n4370), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[236][11]  (.Q(\ram[236][11] ), 
	.D(FE_PHN5177_n4369), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[236][10]  (.Q(\ram[236][10] ), 
	.D(FE_PHN4640_n4368), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[236][9]  (.Q(\ram[236][9] ), 
	.D(FE_PHN4091_n4367), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[236][8]  (.Q(\ram[236][8] ), 
	.D(FE_PHN4733_n4366), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[236][7]  (.Q(\ram[236][7] ), 
	.D(FE_PHN6666_n4365), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[236][6]  (.Q(\ram[236][6] ), 
	.D(FE_PHN4660_n4364), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[236][5]  (.Q(\ram[236][5] ), 
	.D(FE_PHN4226_n4363), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][4]  (.Q(\ram[236][4] ), 
	.D(FE_PHN4277_n4362), 
	.CK(clk_m__L3_N50));
   QDFFEHD \ram_reg[236][3]  (.Q(\ram[236][3] ), 
	.D(FE_PHN4278_n4361), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[236][2]  (.Q(\ram[236][2] ), 
	.D(FE_PHN3427_n4360), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[236][1]  (.Q(\ram[236][1] ), 
	.D(FE_PHN4074_n4359), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[236][0]  (.Q(\ram[236][0] ), 
	.D(FE_PHN4377_n4358), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[232][15]  (.Q(\ram[232][15] ), 
	.D(FE_PHN2366_n4309), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[232][14]  (.Q(\ram[232][14] ), 
	.D(FE_PHN4492_n4308), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[232][13]  (.Q(\ram[232][13] ), 
	.D(FE_PHN4264_n4307), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[232][12]  (.Q(\ram[232][12] ), 
	.D(FE_PHN1390_n4306), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][11]  (.Q(\ram[232][11] ), 
	.D(FE_PHN2793_n4305), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[232][10]  (.Q(\ram[232][10] ), 
	.D(FE_PHN3000_n4304), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][9]  (.Q(\ram[232][9] ), 
	.D(FE_PHN1929_n4303), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][8]  (.Q(\ram[232][8] ), 
	.D(FE_PHN740_n4302), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][7]  (.Q(\ram[232][7] ), 
	.D(FE_PHN2263_n4301), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][6]  (.Q(\ram[232][6] ), 
	.D(FE_PHN5144_n4300), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[232][5]  (.Q(\ram[232][5] ), 
	.D(FE_PHN4661_n4299), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[232][4]  (.Q(\ram[232][4] ), 
	.D(FE_PHN1988_n4298), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[232][3]  (.Q(\ram[232][3] ), 
	.D(FE_PHN471_n4297), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[232][2]  (.Q(\ram[232][2] ), 
	.D(FE_PHN576_n4296), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[232][1]  (.Q(\ram[232][1] ), 
	.D(FE_PHN4119_n4295), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[232][0]  (.Q(\ram[232][0] ), 
	.D(FE_PHN4516_n4294), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[228][15]  (.Q(\ram[228][15] ), 
	.D(FE_PHN5535_n4245), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[228][14]  (.Q(\ram[228][14] ), 
	.D(FE_PHN4301_n4244), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[228][13]  (.Q(\ram[228][13] ), 
	.D(FE_PHN4561_n4243), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[228][12]  (.Q(\ram[228][12] ), 
	.D(FE_PHN4402_n4242), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[228][11]  (.Q(\ram[228][11] ), 
	.D(FE_PHN4619_n4241), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][10]  (.Q(\ram[228][10] ), 
	.D(FE_PHN4703_n4240), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][9]  (.Q(\ram[228][9] ), 
	.D(FE_PHN5484_n4239), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][8]  (.Q(\ram[228][8] ), 
	.D(FE_PHN4116_n4238), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[228][7]  (.Q(\ram[228][7] ), 
	.D(FE_PHN1783_n4237), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[228][6]  (.Q(\ram[228][6] ), 
	.D(FE_PHN4736_n4236), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[228][5]  (.Q(\ram[228][5] ), 
	.D(FE_PHN4721_n4235), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[228][4]  (.Q(\ram[228][4] ), 
	.D(FE_PHN1679_n4234), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[228][3]  (.Q(\ram[228][3] ), 
	.D(FE_PHN4718_n4233), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[228][2]  (.Q(\ram[228][2] ), 
	.D(FE_PHN4597_n4232), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[228][1]  (.Q(\ram[228][1] ), 
	.D(FE_PHN4589_n4231), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[228][0]  (.Q(\ram[228][0] ), 
	.D(FE_PHN5517_n4230), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][15]  (.Q(\ram[224][15] ), 
	.D(FE_PHN4573_n4181), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][14]  (.Q(\ram[224][14] ), 
	.D(FE_PHN3299_n4180), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][13]  (.Q(\ram[224][13] ), 
	.D(FE_PHN3541_n4179), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][12]  (.Q(\ram[224][12] ), 
	.D(FE_PHN4685_n4178), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][11]  (.Q(\ram[224][11] ), 
	.D(FE_PHN1214_n4177), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][10]  (.Q(\ram[224][10] ), 
	.D(FE_PHN2800_n4176), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[224][9]  (.Q(\ram[224][9] ), 
	.D(FE_PHN4753_n4175), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][8]  (.Q(\ram[224][8] ), 
	.D(FE_PHN3415_n4174), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][7]  (.Q(\ram[224][7] ), 
	.D(FE_PHN3121_n4173), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[224][6]  (.Q(\ram[224][6] ), 
	.D(FE_PHN4618_n4172), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[224][5]  (.Q(\ram[224][5] ), 
	.D(FE_PHN4716_n4171), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[224][4]  (.Q(\ram[224][4] ), 
	.D(FE_PHN4751_n4170), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][3]  (.Q(\ram[224][3] ), 
	.D(FE_PHN4570_n4169), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[224][2]  (.Q(\ram[224][2] ), 
	.D(FE_PHN3948_n4168), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[224][1]  (.Q(\ram[224][1] ), 
	.D(FE_PHN4263_n4167), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[224][0]  (.Q(\ram[224][0] ), 
	.D(FE_PHN4433_n4166), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[220][15]  (.Q(\ram[220][15] ), 
	.D(FE_PHN2055_n4117), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][14]  (.Q(\ram[220][14] ), 
	.D(FE_PHN4526_n4116), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][13]  (.Q(\ram[220][13] ), 
	.D(FE_PHN1961_n4115), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][12]  (.Q(\ram[220][12] ), 
	.D(FE_PHN5668_n4114), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][11]  (.Q(\ram[220][11] ), 
	.D(FE_PHN742_n4113), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][10]  (.Q(\ram[220][10] ), 
	.D(FE_PHN1020_n4112), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][9]  (.Q(\ram[220][9] ), 
	.D(FE_PHN4166_n4111), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][8]  (.Q(\ram[220][8] ), 
	.D(FE_PHN4222_n4110), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][7]  (.Q(\ram[220][7] ), 
	.D(FE_PHN2990_n4109), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][6]  (.Q(\ram[220][6] ), 
	.D(FE_PHN1368_n4108), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[220][5]  (.Q(\ram[220][5] ), 
	.D(FE_PHN5656_n4107), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[220][4]  (.Q(\ram[220][4] ), 
	.D(FE_PHN439_n4106), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][3]  (.Q(\ram[220][3] ), 
	.D(FE_PHN239_n4105), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[220][2]  (.Q(\ram[220][2] ), 
	.D(FE_PHN2978_n4104), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[220][1]  (.Q(\ram[220][1] ), 
	.D(FE_PHN3713_n4103), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[220][0]  (.Q(\ram[220][0] ), 
	.D(FE_PHN6678_n4102), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[216][15]  (.Q(\ram[216][15] ), 
	.D(FE_PHN977_n4053), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][14]  (.Q(\ram[216][14] ), 
	.D(FE_PHN1749_n4052), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][13]  (.Q(\ram[216][13] ), 
	.D(FE_PHN1350_n4051), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][12]  (.Q(\ram[216][12] ), 
	.D(FE_PHN2570_n4050), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][11]  (.Q(\ram[216][11] ), 
	.D(FE_PHN4623_n4049), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[216][10]  (.Q(\ram[216][10] ), 
	.D(FE_PHN1049_n4048), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][9]  (.Q(\ram[216][9] ), 
	.D(FE_PHN2674_n4047), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[216][8]  (.Q(\ram[216][8] ), 
	.D(FE_PHN4677_n4046), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][7]  (.Q(\ram[216][7] ), 
	.D(FE_PHN1779_n4045), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][6]  (.Q(\ram[216][6] ), 
	.D(FE_PHN541_n4044), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[216][5]  (.Q(\ram[216][5] ), 
	.D(FE_PHN3086_n4043), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[216][4]  (.Q(\ram[216][4] ), 
	.D(FE_PHN2213_n4042), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[216][3]  (.Q(\ram[216][3] ), 
	.D(FE_PHN1719_n4041), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][2]  (.Q(\ram[216][2] ), 
	.D(FE_PHN1044_n4040), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][1]  (.Q(\ram[216][1] ), 
	.D(FE_PHN1651_n4039), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[216][0]  (.Q(\ram[216][0] ), 
	.D(FE_PHN340_n4038), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[212][15]  (.Q(\ram[212][15] ), 
	.D(FE_PHN4546_n3989), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[212][14]  (.Q(\ram[212][14] ), 
	.D(FE_PHN4322_n3988), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][13]  (.Q(\ram[212][13] ), 
	.D(FE_PHN5214_n3987), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][12]  (.Q(\ram[212][12] ), 
	.D(FE_PHN253_n3986), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][11]  (.Q(\ram[212][11] ), 
	.D(FE_PHN4434_n3985), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][10]  (.Q(\ram[212][10] ), 
	.D(FE_PHN4320_n3984), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][9]  (.Q(\ram[212][9] ), 
	.D(FE_PHN4292_n3983), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][8]  (.Q(\ram[212][8] ), 
	.D(FE_PHN4137_n3982), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][7]  (.Q(\ram[212][7] ), 
	.D(FE_PHN5709_n3981), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][6]  (.Q(\ram[212][6] ), 
	.D(FE_PHN4674_n3980), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][5]  (.Q(\ram[212][5] ), 
	.D(FE_PHN4146_n3979), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[212][4]  (.Q(\ram[212][4] ), 
	.D(FE_PHN4169_n3978), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[212][3]  (.Q(\ram[212][3] ), 
	.D(FE_PHN4310_n3977), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][2]  (.Q(\ram[212][2] ), 
	.D(FE_PHN4662_n3976), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[212][1]  (.Q(\ram[212][1] ), 
	.D(FE_PHN5163_n3975), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[212][0]  (.Q(\ram[212][0] ), 
	.D(FE_PHN4383_n3974), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[208][15]  (.Q(\ram[208][15] ), 
	.D(FE_PHN824_n3925), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[208][14]  (.Q(\ram[208][14] ), 
	.D(FE_PHN4669_n3924), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[208][13]  (.Q(\ram[208][13] ), 
	.D(FE_PHN6651_n3923), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][12]  (.Q(\ram[208][12] ), 
	.D(FE_PHN5499_n3922), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][11]  (.Q(\ram[208][11] ), 
	.D(FE_PHN4367_n3921), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[208][10]  (.Q(\ram[208][10] ), 
	.D(FE_PHN4748_n3920), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[208][9]  (.Q(\ram[208][9] ), 
	.D(FE_PHN5182_n3919), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][8]  (.Q(\ram[208][8] ), 
	.D(FE_PHN3681_n3918), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][7]  (.Q(\ram[208][7] ), 
	.D(FE_PHN4741_n3917), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[208][6]  (.Q(\ram[208][6] ), 
	.D(FE_PHN4691_n3916), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][5]  (.Q(\ram[208][5] ), 
	.D(FE_PHN3403_n3915), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[208][4]  (.Q(\ram[208][4] ), 
	.D(FE_PHN5474_n3914), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[208][3]  (.Q(\ram[208][3] ), 
	.D(FE_PHN4502_n3913), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[208][2]  (.Q(\ram[208][2] ), 
	.D(FE_PHN460_n3912), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[208][1]  (.Q(\ram[208][1] ), 
	.D(FE_PHN4240_n3911), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[208][0]  (.Q(\ram[208][0] ), 
	.D(FE_PHN4430_n3910), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[204][15]  (.Q(\ram[204][15] ), 
	.D(FE_PHN314_n3861), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][14]  (.Q(\ram[204][14] ), 
	.D(FE_PHN2795_n3860), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][13]  (.Q(\ram[204][13] ), 
	.D(FE_PHN1174_n3859), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[204][12]  (.Q(\ram[204][12] ), 
	.D(FE_PHN2309_n3858), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][11]  (.Q(\ram[204][11] ), 
	.D(FE_PHN327_n3857), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][10]  (.Q(\ram[204][10] ), 
	.D(FE_PHN2601_n3856), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][9]  (.Q(\ram[204][9] ), 
	.D(FE_PHN2397_n3855), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][8]  (.Q(\ram[204][8] ), 
	.D(FE_PHN3092_n3854), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][7]  (.Q(\ram[204][7] ), 
	.D(FE_PHN737_n3853), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][6]  (.Q(\ram[204][6] ), 
	.D(FE_PHN1936_n3852), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[204][5]  (.Q(\ram[204][5] ), 
	.D(FE_PHN1179_n3851), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][4]  (.Q(\ram[204][4] ), 
	.D(FE_PHN1844_n3850), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][3]  (.Q(\ram[204][3] ), 
	.D(FE_PHN2328_n3849), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][2]  (.Q(\ram[204][2] ), 
	.D(FE_PHN3206_n3848), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[204][1]  (.Q(\ram[204][1] ), 
	.D(FE_PHN1751_n3847), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[204][0]  (.Q(\ram[204][0] ), 
	.D(FE_PHN3192_n3846), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[200][15]  (.Q(\ram[200][15] ), 
	.D(FE_PHN3134_n3797), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[200][14]  (.Q(\ram[200][14] ), 
	.D(FE_PHN778_n3796), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][13]  (.Q(\ram[200][13] ), 
	.D(FE_PHN2529_n3795), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][12]  (.Q(\ram[200][12] ), 
	.D(FE_PHN993_n3794), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[200][11]  (.Q(\ram[200][11] ), 
	.D(FE_PHN1628_n3793), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][10]  (.Q(\ram[200][10] ), 
	.D(FE_PHN2646_n3792), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[200][9]  (.Q(\ram[200][9] ), 
	.D(FE_PHN2543_n3791), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][8]  (.Q(\ram[200][8] ), 
	.D(FE_PHN1963_n3790), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][7]  (.Q(\ram[200][7] ), 
	.D(FE_PHN1541_n3789), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][6]  (.Q(\ram[200][6] ), 
	.D(FE_PHN1294_n3788), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][5]  (.Q(\ram[200][5] ), 
	.D(FE_PHN1813_n3787), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][4]  (.Q(\ram[200][4] ), 
	.D(FE_PHN2933_n3786), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][3]  (.Q(\ram[200][3] ), 
	.D(FE_PHN1660_n3785), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][2]  (.Q(\ram[200][2] ), 
	.D(FE_PHN3119_n3784), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[200][1]  (.Q(\ram[200][1] ), 
	.D(FE_PHN338_n3783), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[200][0]  (.Q(\ram[200][0] ), 
	.D(FE_PHN2616_n3782), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[196][15]  (.Q(\ram[196][15] ), 
	.D(FE_PHN709_n3733), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[196][14]  (.Q(\ram[196][14] ), 
	.D(FE_PHN1483_n3732), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][13]  (.Q(\ram[196][13] ), 
	.D(FE_PHN2285_n3731), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[196][12]  (.Q(\ram[196][12] ), 
	.D(FE_PHN301_n3730), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[196][11]  (.Q(\ram[196][11] ), 
	.D(FE_PHN2053_n3729), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][10]  (.Q(\ram[196][10] ), 
	.D(FE_PHN1167_n3728), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][9]  (.Q(\ram[196][9] ), 
	.D(FE_PHN2182_n3727), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[196][8]  (.Q(\ram[196][8] ), 
	.D(FE_PHN987_n3726), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][7]  (.Q(\ram[196][7] ), 
	.D(FE_PHN1285_n3725), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][6]  (.Q(\ram[196][6] ), 
	.D(FE_PHN811_n3724), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][5]  (.Q(\ram[196][5] ), 
	.D(FE_PHN2362_n3723), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][4]  (.Q(\ram[196][4] ), 
	.D(FE_PHN2467_n3722), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][3]  (.Q(\ram[196][3] ), 
	.D(FE_PHN1062_n3721), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[196][2]  (.Q(\ram[196][2] ), 
	.D(FE_PHN853_n3720), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[196][1]  (.Q(\ram[196][1] ), 
	.D(FE_PHN1930_n3719), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[196][0]  (.Q(\ram[196][0] ), 
	.D(FE_PHN1773_n3718), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[192][15]  (.Q(\ram[192][15] ), 
	.D(FE_PHN2818_n3669), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][14]  (.Q(\ram[192][14] ), 
	.D(FE_PHN2749_n3668), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][13]  (.Q(\ram[192][13] ), 
	.D(FE_PHN1877_n3667), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][12]  (.Q(\ram[192][12] ), 
	.D(FE_PHN1734_n3666), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][11]  (.Q(\ram[192][11] ), 
	.D(FE_PHN2747_n3665), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][10]  (.Q(\ram[192][10] ), 
	.D(FE_PHN2184_n3664), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][9]  (.Q(\ram[192][9] ), 
	.D(FE_PHN596_n3663), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][8]  (.Q(\ram[192][8] ), 
	.D(FE_PHN1790_n3662), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][7]  (.Q(\ram[192][7] ), 
	.D(FE_PHN1857_n3661), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][6]  (.Q(\ram[192][6] ), 
	.D(FE_PHN1629_n3660), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][5]  (.Q(\ram[192][5] ), 
	.D(FE_PHN2310_n3659), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][4]  (.Q(\ram[192][4] ), 
	.D(FE_PHN1478_n3658), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][3]  (.Q(\ram[192][3] ), 
	.D(FE_PHN2630_n3657), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[192][2]  (.Q(\ram[192][2] ), 
	.D(FE_PHN2387_n3656), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[192][1]  (.Q(\ram[192][1] ), 
	.D(FE_PHN2085_n3655), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[192][0]  (.Q(\ram[192][0] ), 
	.D(FE_PHN2513_n3654), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[188][15]  (.Q(\ram[188][15] ), 
	.D(FE_PHN1858_n3605), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][14]  (.Q(\ram[188][14] ), 
	.D(FE_PHN1067_n3604), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][13]  (.Q(\ram[188][13] ), 
	.D(FE_PHN2502_n3603), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][12]  (.Q(\ram[188][12] ), 
	.D(FE_PHN2163_n3602), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][11]  (.Q(\ram[188][11] ), 
	.D(FE_PHN1884_n3601), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[188][10]  (.Q(\ram[188][10] ), 
	.D(FE_PHN1635_n3600), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][9]  (.Q(\ram[188][9] ), 
	.D(FE_PHN2206_n3599), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[188][8]  (.Q(\ram[188][8] ), 
	.D(FE_PHN2912_n3598), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][7]  (.Q(\ram[188][7] ), 
	.D(FE_PHN2194_n3597), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][6]  (.Q(\ram[188][6] ), 
	.D(FE_PHN1525_n3596), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][5]  (.Q(\ram[188][5] ), 
	.D(FE_PHN1110_n3595), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][4]  (.Q(\ram[188][4] ), 
	.D(FE_PHN2081_n3594), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][3]  (.Q(\ram[188][3] ), 
	.D(FE_PHN1798_n3593), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[188][2]  (.Q(\ram[188][2] ), 
	.D(FE_PHN3205_n3592), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[188][1]  (.Q(\ram[188][1] ), 
	.D(FE_PHN638_n3591), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[188][0]  (.Q(\ram[188][0] ), 
	.D(FE_PHN2022_n3590), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][15]  (.Q(\ram[184][15] ), 
	.D(FE_PHN3183_n3541), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][14]  (.Q(\ram[184][14] ), 
	.D(FE_PHN2939_n3540), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][13]  (.Q(\ram[184][13] ), 
	.D(FE_PHN1534_n3539), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[184][12]  (.Q(\ram[184][12] ), 
	.D(FE_PHN119_n3538), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[184][11]  (.Q(\ram[184][11] ), 
	.D(FE_PHN569_n3537), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][10]  (.Q(\ram[184][10] ), 
	.D(FE_PHN305_n3536), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][9]  (.Q(\ram[184][9] ), 
	.D(FE_PHN3108_n3535), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][8]  (.Q(\ram[184][8] ), 
	.D(FE_PHN489_n3534), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][7]  (.Q(\ram[184][7] ), 
	.D(FE_PHN113_n3533), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[184][6]  (.Q(\ram[184][6] ), 
	.D(FE_PHN319_n3532), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[184][5]  (.Q(\ram[184][5] ), 
	.D(FE_PHN359_n3531), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[184][4]  (.Q(\ram[184][4] ), 
	.D(FE_PHN919_n3530), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[184][3]  (.Q(\ram[184][3] ), 
	.D(FE_PHN1403_n3529), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[184][2]  (.Q(\ram[184][2] ), 
	.D(FE_PHN821_n3528), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][1]  (.Q(\ram[184][1] ), 
	.D(FE_PHN1818_n3527), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[184][0]  (.Q(\ram[184][0] ), 
	.D(FE_PHN403_n3526), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[180][15]  (.Q(\ram[180][15] ), 
	.D(FE_PHN2063_n3477), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[180][14]  (.Q(\ram[180][14] ), 
	.D(FE_PHN2318_n3476), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[180][13]  (.Q(\ram[180][13] ), 
	.D(FE_PHN2827_n3475), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[180][12]  (.Q(\ram[180][12] ), 
	.D(FE_PHN2142_n3474), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][11]  (.Q(\ram[180][11] ), 
	.D(FE_PHN486_n3473), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[180][10]  (.Q(\ram[180][10] ), 
	.D(FE_PHN561_n3472), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][9]  (.Q(\ram[180][9] ), 
	.D(FE_PHN3168_n3471), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][8]  (.Q(\ram[180][8] ), 
	.D(FE_PHN562_n3470), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][7]  (.Q(\ram[180][7] ), 
	.D(FE_PHN3203_n3469), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][6]  (.Q(\ram[180][6] ), 
	.D(FE_PHN597_n3468), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][5]  (.Q(\ram[180][5] ), 
	.D(FE_PHN3095_n3467), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][4]  (.Q(\ram[180][4] ), 
	.D(FE_PHN3003_n3466), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][3]  (.Q(\ram[180][3] ), 
	.D(FE_PHN762_n3465), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[180][2]  (.Q(\ram[180][2] ), 
	.D(FE_PHN1306_n3464), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[180][1]  (.Q(\ram[180][1] ), 
	.D(FE_PHN520_n3463), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[180][0]  (.Q(\ram[180][0] ), 
	.D(FE_PHN3030_n3462), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[176][15]  (.Q(\ram[176][15] ), 
	.D(FE_PHN2275_n3413), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[176][14]  (.Q(\ram[176][14] ), 
	.D(FE_PHN1787_n3412), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][13]  (.Q(\ram[176][13] ), 
	.D(FE_PHN1153_n3411), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[176][12]  (.Q(\ram[176][12] ), 
	.D(FE_PHN2065_n3410), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[176][11]  (.Q(\ram[176][11] ), 
	.D(FE_PHN2734_n3409), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[176][10]  (.Q(\ram[176][10] ), 
	.D(FE_PHN2487_n3408), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[176][9]  (.Q(\ram[176][9] ), 
	.D(FE_PHN1845_n3407), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][8]  (.Q(\ram[176][8] ), 
	.D(FE_PHN1211_n3406), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[176][7]  (.Q(\ram[176][7] ), 
	.D(FE_PHN2211_n3405), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][6]  (.Q(\ram[176][6] ), 
	.D(FE_PHN864_n3404), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][5]  (.Q(\ram[176][5] ), 
	.D(FE_PHN1038_n3403), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][4]  (.Q(\ram[176][4] ), 
	.D(FE_PHN2457_n3402), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][3]  (.Q(\ram[176][3] ), 
	.D(FE_PHN2627_n3401), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][2]  (.Q(\ram[176][2] ), 
	.D(FE_PHN2293_n3400), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[176][1]  (.Q(\ram[176][1] ), 
	.D(FE_PHN1488_n3399), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[176][0]  (.Q(\ram[176][0] ), 
	.D(FE_PHN1187_n3398), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[172][15]  (.Q(\ram[172][15] ), 
	.D(FE_PHN755_n3349), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[172][14]  (.Q(\ram[172][14] ), 
	.D(FE_PHN1089_n3348), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][13]  (.Q(\ram[172][13] ), 
	.D(FE_PHN1450_n3347), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[172][12]  (.Q(\ram[172][12] ), 
	.D(FE_PHN1132_n3346), 
	.CK(clk));
   QDFFEHD \ram_reg[172][11]  (.Q(\ram[172][11] ), 
	.D(FE_PHN2166_n3345), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[172][10]  (.Q(\ram[172][10] ), 
	.D(FE_PHN615_n3344), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[172][9]  (.Q(\ram[172][9] ), 
	.D(FE_PHN2894_n3343), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][8]  (.Q(\ram[172][8] ), 
	.D(FE_PHN1367_n3342), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[172][7]  (.Q(\ram[172][7] ), 
	.D(FE_PHN2390_n3341), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[172][6]  (.Q(\ram[172][6] ), 
	.D(FE_PHN1159_n3340), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][5]  (.Q(\ram[172][5] ), 
	.D(FE_PHN1040_n3339), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[172][4]  (.Q(\ram[172][4] ), 
	.D(FE_PHN2587_n3338), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[172][3]  (.Q(\ram[172][3] ), 
	.D(FE_PHN504_n3337), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[172][2]  (.Q(\ram[172][2] ), 
	.D(FE_PHN1475_n3336), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[172][1]  (.Q(\ram[172][1] ), 
	.D(FE_PHN1622_n3335), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[172][0]  (.Q(\ram[172][0] ), 
	.D(FE_PHN1449_n3334), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][15]  (.Q(\ram[168][15] ), 
	.D(FE_PHN2822_n3285), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][14]  (.Q(\ram[168][14] ), 
	.D(FE_PHN3207_n3284), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][13]  (.Q(\ram[168][13] ), 
	.D(FE_PHN1342_n3283), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][12]  (.Q(\ram[168][12] ), 
	.D(FE_PHN1497_n3282), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][11]  (.Q(\ram[168][11] ), 
	.D(FE_PHN1738_n3281), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[168][10]  (.Q(\ram[168][10] ), 
	.D(FE_PHN3167_n3280), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[168][9]  (.Q(\ram[168][9] ), 
	.D(FE_PHN1098_n3279), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][8]  (.Q(\ram[168][8] ), 
	.D(FE_PHN1825_n3278), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[168][7]  (.Q(\ram[168][7] ), 
	.D(FE_PHN738_n3277), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[168][6]  (.Q(\ram[168][6] ), 
	.D(FE_PHN1513_n3276), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][5]  (.Q(\ram[168][5] ), 
	.D(FE_PHN2921_n3275), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[168][4]  (.Q(\ram[168][4] ), 
	.D(FE_PHN483_n3274), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[168][3]  (.Q(\ram[168][3] ), 
	.D(FE_PHN1004_n3273), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[168][2]  (.Q(\ram[168][2] ), 
	.D(FE_PHN2762_n3272), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[168][1]  (.Q(\ram[168][1] ), 
	.D(FE_PHN836_n3271), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[168][0]  (.Q(\ram[168][0] ), 
	.D(FE_PHN1777_n3270), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[164][15]  (.Q(\ram[164][15] ), 
	.D(FE_PHN1960_n3221), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[164][14]  (.Q(\ram[164][14] ), 
	.D(FE_PHN3122_n3220), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][13]  (.Q(\ram[164][13] ), 
	.D(FE_PHN5217_n3219), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[164][12]  (.Q(\ram[164][12] ), 
	.D(FE_PHN1423_n3218), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][11]  (.Q(\ram[164][11] ), 
	.D(FE_PHN5083_n3217), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[164][10]  (.Q(\ram[164][10] ), 
	.D(FE_PHN1700_n3216), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[164][9]  (.Q(\ram[164][9] ), 
	.D(FE_PHN1259_n3215), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][8]  (.Q(\ram[164][8] ), 
	.D(FE_PHN1136_n3214), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][7]  (.Q(\ram[164][7] ), 
	.D(FE_PHN188_n3213), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[164][6]  (.Q(\ram[164][6] ), 
	.D(FE_PHN4519_n3212), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][5]  (.Q(\ram[164][5] ), 
	.D(FE_PHN1901_n3211), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][4]  (.Q(\ram[164][4] ), 
	.D(FE_PHN4708_n3210), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[164][3]  (.Q(\ram[164][3] ), 
	.D(FE_PHN558_n3209), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][2]  (.Q(\ram[164][2] ), 
	.D(FE_PHN1575_n3208), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[164][1]  (.Q(\ram[164][1] ), 
	.D(FE_PHN4535_n3207), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[164][0]  (.Q(\ram[164][0] ), 
	.D(FE_PHN1742_n3206), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][15]  (.Q(\ram[160][15] ), 
	.D(FE_PHN2562_n3157), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][14]  (.Q(\ram[160][14] ), 
	.D(FE_PHN414_n3156), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][13]  (.Q(\ram[160][13] ), 
	.D(FE_PHN1047_n3155), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][12]  (.Q(\ram[160][12] ), 
	.D(FE_PHN1279_n3154), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][11]  (.Q(\ram[160][11] ), 
	.D(FE_PHN2541_n3153), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][10]  (.Q(\ram[160][10] ), 
	.D(FE_PHN3213_n3152), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][9]  (.Q(\ram[160][9] ), 
	.D(FE_PHN2537_n3151), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[160][8]  (.Q(\ram[160][8] ), 
	.D(FE_PHN5688_n3150), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[160][7]  (.Q(\ram[160][7] ), 
	.D(FE_PHN2440_n3149), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][6]  (.Q(\ram[160][6] ), 
	.D(FE_PHN2356_n3148), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][5]  (.Q(\ram[160][5] ), 
	.D(FE_PHN1446_n3147), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[160][4]  (.Q(\ram[160][4] ), 
	.D(FE_PHN1774_n3146), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[160][3]  (.Q(\ram[160][3] ), 
	.D(FE_PHN1300_n3145), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][2]  (.Q(\ram[160][2] ), 
	.D(FE_PHN2446_n3144), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[160][1]  (.Q(\ram[160][1] ), 
	.D(FE_PHN3116_n3143), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[160][0]  (.Q(\ram[160][0] ), 
	.D(FE_PHN2832_n3142), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[156][15]  (.Q(\ram[156][15] ), 
	.D(FE_PHN4351_n3093), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][14]  (.Q(\ram[156][14] ), 
	.D(FE_PHN4079_n3092), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][13]  (.Q(\ram[156][13] ), 
	.D(FE_PHN5573_n3091), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][12]  (.Q(\ram[156][12] ), 
	.D(FE_PHN4332_n3090), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][11]  (.Q(\ram[156][11] ), 
	.D(FE_PHN4206_n3089), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[156][10]  (.Q(\ram[156][10] ), 
	.D(FE_PHN4532_n3088), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[156][9]  (.Q(\ram[156][9] ), 
	.D(FE_PHN4287_n3087), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[156][8]  (.Q(\ram[156][8] ), 
	.D(FE_PHN4659_n3086), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[156][7]  (.Q(\ram[156][7] ), 
	.D(FE_PHN4318_n3085), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[156][6]  (.Q(\ram[156][6] ), 
	.D(FE_PHN5503_n3084), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[156][5]  (.Q(\ram[156][5] ), 
	.D(FE_PHN4252_n3083), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[156][4]  (.Q(\ram[156][4] ), 
	.D(FE_PHN4584_n3082), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[156][3]  (.Q(\ram[156][3] ), 
	.D(FE_PHN4120_n3081), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[156][2]  (.Q(\ram[156][2] ), 
	.D(FE_PHN4379_n3080), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[156][1]  (.Q(\ram[156][1] ), 
	.D(FE_PHN3889_n3079), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[156][0]  (.Q(\ram[156][0] ), 
	.D(FE_PHN5473_n3078), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[152][15]  (.Q(\ram[152][15] ), 
	.D(FE_PHN5237_n3029), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[152][14]  (.Q(\ram[152][14] ), 
	.D(FE_PHN3759_n3028), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[152][13]  (.Q(\ram[152][13] ), 
	.D(FE_PHN4187_n3027), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[152][12]  (.Q(\ram[152][12] ), 
	.D(FE_PHN4173_n3026), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[152][11]  (.Q(\ram[152][11] ), 
	.D(FE_PHN5314_n3025), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[152][10]  (.Q(\ram[152][10] ), 
	.D(FE_PHN3612_n3024), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[152][9]  (.Q(\ram[152][9] ), 
	.D(FE_PHN5289_n3023), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[152][8]  (.Q(\ram[152][8] ), 
	.D(FE_PHN4049_n3022), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[152][7]  (.Q(\ram[152][7] ), 
	.D(FE_PHN4937_n3021), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][6]  (.Q(\ram[152][6] ), 
	.D(FE_PHN4639_n3020), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[152][5]  (.Q(\ram[152][5] ), 
	.D(FE_PHN4127_n3019), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[152][4]  (.Q(\ram[152][4] ), 
	.D(FE_PHN4524_n3018), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[152][3]  (.Q(\ram[152][3] ), 
	.D(FE_PHN4944_n3017), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][2]  (.Q(\ram[152][2] ), 
	.D(FE_PHN4469_n3016), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][1]  (.Q(\ram[152][1] ), 
	.D(FE_PHN4598_n3015), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[152][0]  (.Q(\ram[152][0] ), 
	.D(FE_PHN4372_n3014), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[148][15]  (.Q(\ram[148][15] ), 
	.D(FE_PHN4645_n2965), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][14]  (.Q(\ram[148][14] ), 
	.D(FE_PHN3490_n2964), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][13]  (.Q(\ram[148][13] ), 
	.D(FE_PHN4648_n2963), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][12]  (.Q(\ram[148][12] ), 
	.D(FE_PHN4970_n2962), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][11]  (.Q(\ram[148][11] ), 
	.D(FE_PHN4102_n2961), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[148][10]  (.Q(\ram[148][10] ), 
	.D(FE_PHN4395_n2960), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[148][9]  (.Q(\ram[148][9] ), 
	.D(FE_PHN4408_n2959), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[148][8]  (.Q(\ram[148][8] ), 
	.D(FE_PHN4215_n2958), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[148][7]  (.Q(\ram[148][7] ), 
	.D(FE_PHN4720_n2957), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[148][6]  (.Q(\ram[148][6] ), 
	.D(FE_PHN4084_n2956), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[148][5]  (.Q(\ram[148][5] ), 
	.D(FE_PHN4090_n2955), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[148][4]  (.Q(\ram[148][4] ), 
	.D(FE_PHN4523_n2954), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[148][3]  (.Q(\ram[148][3] ), 
	.D(FE_PHN4265_n2953), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[148][2]  (.Q(\ram[148][2] ), 
	.D(FE_PHN4211_n2952), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[148][1]  (.Q(\ram[148][1] ), 
	.D(FE_PHN4497_n2951), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[148][0]  (.Q(\ram[148][0] ), 
	.D(FE_PHN4644_n2950), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[144][15]  (.Q(\ram[144][15] ), 
	.D(FE_PHN310_n2901), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[144][14]  (.Q(\ram[144][14] ), 
	.D(FE_PHN4269_n2900), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][13]  (.Q(\ram[144][13] ), 
	.D(FE_PHN840_n2899), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[144][12]  (.Q(\ram[144][12] ), 
	.D(FE_PHN4529_n2898), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[144][11]  (.Q(\ram[144][11] ), 
	.D(FE_PHN5253_n2897), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][10]  (.Q(\ram[144][10] ), 
	.D(FE_PHN5506_n2896), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[144][9]  (.Q(\ram[144][9] ), 
	.D(FE_PHN627_n2895), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][8]  (.Q(\ram[144][8] ), 
	.D(n2894), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[144][7]  (.Q(\ram[144][7] ), 
	.D(FE_PHN5744_n2893), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][6]  (.Q(\ram[144][6] ), 
	.D(FE_PHN6664_n2892), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][5]  (.Q(\ram[144][5] ), 
	.D(FE_PHN4596_n2891), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][4]  (.Q(\ram[144][4] ), 
	.D(FE_PHN4888_n2890), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][3]  (.Q(\ram[144][3] ), 
	.D(FE_PHN4864_n2889), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[144][2]  (.Q(\ram[144][2] ), 
	.D(FE_PHN4693_n2888), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[144][1]  (.Q(\ram[144][1] ), 
	.D(FE_PHN4804_n2887), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[144][0]  (.Q(\ram[144][0] ), 
	.D(FE_PHN4709_n2886), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[140][15]  (.Q(\ram[140][15] ), 
	.D(FE_PHN1265_n2837), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][14]  (.Q(\ram[140][14] ), 
	.D(FE_PHN979_n2836), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][13]  (.Q(\ram[140][13] ), 
	.D(FE_PHN818_n2835), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][12]  (.Q(\ram[140][12] ), 
	.D(FE_PHN1676_n2834), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[140][11]  (.Q(\ram[140][11] ), 
	.D(FE_PHN1158_n2833), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[140][10]  (.Q(\ram[140][10] ), 
	.D(FE_PHN2008_n2832), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[140][9]  (.Q(\ram[140][9] ), 
	.D(FE_PHN1189_n2831), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[140][8]  (.Q(\ram[140][8] ), 
	.D(FE_PHN1891_n2830), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[140][7]  (.Q(\ram[140][7] ), 
	.D(FE_PHN2374_n2829), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[140][6]  (.Q(\ram[140][6] ), 
	.D(FE_PHN1711_n2828), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[140][5]  (.Q(\ram[140][5] ), 
	.D(FE_PHN1810_n2827), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[140][4]  (.Q(\ram[140][4] ), 
	.D(FE_PHN581_n2826), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[140][3]  (.Q(\ram[140][3] ), 
	.D(FE_PHN1161_n2825), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[140][2]  (.Q(\ram[140][2] ), 
	.D(FE_PHN2287_n2824), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[140][1]  (.Q(\ram[140][1] ), 
	.D(FE_PHN1245_n2823), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[140][0]  (.Q(\ram[140][0] ), 
	.D(FE_PHN1412_n2822), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[136][15]  (.Q(\ram[136][15] ), 
	.D(FE_PHN3112_n2773), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][14]  (.Q(\ram[136][14] ), 
	.D(FE_PHN1855_n2772), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][13]  (.Q(\ram[136][13] ), 
	.D(FE_PHN2460_n2771), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[136][12]  (.Q(\ram[136][12] ), 
	.D(FE_PHN392_n2770), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][11]  (.Q(\ram[136][11] ), 
	.D(FE_PHN2789_n2769), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][10]  (.Q(\ram[136][10] ), 
	.D(FE_PHN2030_n2768), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[136][9]  (.Q(\ram[136][9] ), 
	.D(FE_PHN1429_n2767), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][8]  (.Q(\ram[136][8] ), 
	.D(FE_PHN2817_n2766), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[136][7]  (.Q(\ram[136][7] ), 
	.D(FE_PHN463_n2765), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[136][6]  (.Q(\ram[136][6] ), 
	.D(FE_PHN1752_n2764), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[136][5]  (.Q(\ram[136][5] ), 
	.D(FE_PHN1224_n2763), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[136][4]  (.Q(\ram[136][4] ), 
	.D(FE_PHN1559_n2762), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[136][3]  (.Q(\ram[136][3] ), 
	.D(FE_PHN260_n2761), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[136][2]  (.Q(\ram[136][2] ), 
	.D(FE_PHN2706_n2760), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[136][1]  (.Q(\ram[136][1] ), 
	.D(FE_PHN2675_n2759), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[136][0]  (.Q(\ram[136][0] ), 
	.D(FE_PHN2701_n2758), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[132][15]  (.Q(\ram[132][15] ), 
	.D(FE_PHN1898_n2709), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[132][14]  (.Q(\ram[132][14] ), 
	.D(FE_PHN2606_n2708), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[132][13]  (.Q(\ram[132][13] ), 
	.D(FE_PHN2160_n2707), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[132][12]  (.Q(\ram[132][12] ), 
	.D(FE_PHN2458_n2706), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[132][11]  (.Q(\ram[132][11] ), 
	.D(FE_PHN1447_n2705), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[132][10]  (.Q(\ram[132][10] ), 
	.D(FE_PHN1111_n2704), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[132][9]  (.Q(\ram[132][9] ), 
	.D(FE_PHN3496_n2703), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[132][8]  (.Q(\ram[132][8] ), 
	.D(n2702), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[132][7]  (.Q(\ram[132][7] ), 
	.D(FE_PHN5661_n2701), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[132][6]  (.Q(\ram[132][6] ), 
	.D(FE_PHN3128_n2700), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[132][5]  (.Q(\ram[132][5] ), 
	.D(FE_PHN1220_n2699), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[132][4]  (.Q(\ram[132][4] ), 
	.D(FE_PHN1908_n2698), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[132][3]  (.Q(\ram[132][3] ), 
	.D(FE_PHN5761_n2697), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[132][2]  (.Q(\ram[132][2] ), 
	.D(FE_PHN6565_n2696), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[132][1]  (.Q(\ram[132][1] ), 
	.D(FE_PHN5708_n2695), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[132][0]  (.Q(\ram[132][0] ), 
	.D(FE_PHN2169_n2694), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[128][15]  (.Q(\ram[128][15] ), 
	.D(FE_PHN1951_n2645), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][14]  (.Q(\ram[128][14] ), 
	.D(FE_PHN1197_n2644), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][13]  (.Q(\ram[128][13] ), 
	.D(FE_PHN1344_n2643), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][12]  (.Q(\ram[128][12] ), 
	.D(FE_PHN2641_n2642), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[128][11]  (.Q(\ram[128][11] ), 
	.D(FE_PHN1234_n2641), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[128][10]  (.Q(\ram[128][10] ), 
	.D(FE_PHN1655_n2640), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[128][9]  (.Q(\ram[128][9] ), 
	.D(FE_PHN2297_n2639), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[128][8]  (.Q(\ram[128][8] ), 
	.D(FE_PHN920_n2638), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[128][7]  (.Q(\ram[128][7] ), 
	.D(FE_PHN426_n2637), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[128][6]  (.Q(\ram[128][6] ), 
	.D(FE_PHN3099_n2636), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][5]  (.Q(\ram[128][5] ), 
	.D(FE_PHN1641_n2635), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][4]  (.Q(\ram[128][4] ), 
	.D(FE_PHN1468_n2634), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][3]  (.Q(\ram[128][3] ), 
	.D(FE_PHN522_n2633), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][2]  (.Q(\ram[128][2] ), 
	.D(FE_PHN619_n2632), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[128][1]  (.Q(\ram[128][1] ), 
	.D(FE_PHN2476_n2631), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[128][0]  (.Q(\ram[128][0] ), 
	.D(FE_PHN2952_n2630), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[124][15]  (.Q(\ram[124][15] ), 
	.D(FE_PHN2702_n2581), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[124][14]  (.Q(\ram[124][14] ), 
	.D(FE_PHN4671_n2580), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[124][13]  (.Q(\ram[124][13] ), 
	.D(FE_PHN1192_n2579), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[124][12]  (.Q(\ram[124][12] ), 
	.D(FE_PHN6652_n2578), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[124][11]  (.Q(\ram[124][11] ), 
	.D(FE_PHN4953_n2577), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[124][10]  (.Q(\ram[124][10] ), 
	.D(FE_PHN5715_n2576), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[124][9]  (.Q(\ram[124][9] ), 
	.D(FE_PHN2850_n2575), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[124][8]  (.Q(\ram[124][8] ), 
	.D(FE_PHN4582_n2574), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[124][7]  (.Q(\ram[124][7] ), 
	.D(FE_PHN2506_n2573), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[124][6]  (.Q(\ram[124][6] ), 
	.D(FE_PHN5702_n2572), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][5]  (.Q(\ram[124][5] ), 
	.D(FE_PHN6650_n2571), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][4]  (.Q(\ram[124][4] ), 
	.D(FE_PHN6696_n2570), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][3]  (.Q(\ram[124][3] ), 
	.D(FE_PHN2332_n2569), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[124][2]  (.Q(\ram[124][2] ), 
	.D(FE_PHN1544_n2568), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[124][1]  (.Q(\ram[124][1] ), 
	.D(FE_PHN1169_n2567), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[124][0]  (.Q(\ram[124][0] ), 
	.D(FE_PHN6555_n2566), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[120][15]  (.Q(\ram[120][15] ), 
	.D(FE_PHN2831_n2517), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[120][14]  (.Q(\ram[120][14] ), 
	.D(n2516), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[120][13]  (.Q(\ram[120][13] ), 
	.D(FE_PHN1928_n2515), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[120][12]  (.Q(\ram[120][12] ), 
	.D(FE_PHN1339_n2514), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[120][11]  (.Q(\ram[120][11] ), 
	.D(FE_PHN2130_n2513), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[120][10]  (.Q(\ram[120][10] ), 
	.D(FE_PHN2196_n2512), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][9]  (.Q(\ram[120][9] ), 
	.D(FE_PHN3166_n2511), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][8]  (.Q(\ram[120][8] ), 
	.D(FE_PHN2468_n2510), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][7]  (.Q(\ram[120][7] ), 
	.D(FE_PHN2098_n2509), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[120][6]  (.Q(\ram[120][6] ), 
	.D(FE_PHN628_n2508), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[120][5]  (.Q(\ram[120][5] ), 
	.D(FE_PHN671_n2507), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[120][4]  (.Q(\ram[120][4] ), 
	.D(FE_PHN2974_n2506), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[120][3]  (.Q(\ram[120][3] ), 
	.D(FE_PHN3175_n2505), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[120][2]  (.Q(\ram[120][2] ), 
	.D(FE_PHN2565_n2504), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[120][1]  (.Q(\ram[120][1] ), 
	.D(FE_PHN1361_n2503), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[120][0]  (.Q(\ram[120][0] ), 
	.D(FE_PHN2539_n2502), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[116][15]  (.Q(\ram[116][15] ), 
	.D(FE_PHN2857_n2453), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][14]  (.Q(\ram[116][14] ), 
	.D(FE_PHN1703_n2452), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][13]  (.Q(\ram[116][13] ), 
	.D(FE_PHN1886_n2451), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[116][12]  (.Q(\ram[116][12] ), 
	.D(FE_PHN1883_n2450), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[116][11]  (.Q(\ram[116][11] ), 
	.D(FE_PHN2016_n2449), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][10]  (.Q(\ram[116][10] ), 
	.D(FE_PHN2492_n2448), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[116][9]  (.Q(\ram[116][9] ), 
	.D(FE_PHN2683_n2447), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][8]  (.Q(\ram[116][8] ), 
	.D(FE_PHN3131_n2446), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[116][7]  (.Q(\ram[116][7] ), 
	.D(FE_PHN2968_n2445), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][6]  (.Q(\ram[116][6] ), 
	.D(FE_PHN629_n2444), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][5]  (.Q(\ram[116][5] ), 
	.D(FE_PHN2497_n2443), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[116][4]  (.Q(\ram[116][4] ), 
	.D(FE_PHN1128_n2442), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][3]  (.Q(\ram[116][3] ), 
	.D(FE_PHN731_n2441), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][2]  (.Q(\ram[116][2] ), 
	.D(FE_PHN972_n2440), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][1]  (.Q(\ram[116][1] ), 
	.D(FE_PHN886_n2439), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[116][0]  (.Q(\ram[116][0] ), 
	.D(FE_PHN2764_n2438), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[112][15]  (.Q(\ram[112][15] ), 
	.D(FE_PHN4138_n2389), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][14]  (.Q(\ram[112][14] ), 
	.D(FE_PHN4571_n2388), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[112][13]  (.Q(\ram[112][13] ), 
	.D(FE_PHN1022_n2387), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[112][12]  (.Q(\ram[112][12] ), 
	.D(FE_PHN5754_n2386), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][11]  (.Q(\ram[112][11] ), 
	.D(FE_PHN4506_n2385), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][10]  (.Q(\ram[112][10] ), 
	.D(FE_PHN4602_n2384), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][9]  (.Q(\ram[112][9] ), 
	.D(FE_PHN3887_n2383), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][8]  (.Q(\ram[112][8] ), 
	.D(FE_PHN5659_n2382), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][7]  (.Q(\ram[112][7] ), 
	.D(FE_PHN5742_n2381), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[112][6]  (.Q(\ram[112][6] ), 
	.D(FE_PHN5706_n2380), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][5]  (.Q(\ram[112][5] ), 
	.D(FE_PHN6685_n2379), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][4]  (.Q(\ram[112][4] ), 
	.D(FE_PHN6653_n2378), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][3]  (.Q(\ram[112][3] ), 
	.D(FE_PHN6643_n2377), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][2]  (.Q(\ram[112][2] ), 
	.D(FE_PHN5719_n2376), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[112][1]  (.Q(\ram[112][1] ), 
	.D(FE_PHN5654_n2375), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[112][0]  (.Q(\ram[112][0] ), 
	.D(FE_PHN4117_n2374), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[108][15]  (.Q(\ram[108][15] ), 
	.D(FE_PHN1140_n2325), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[108][14]  (.Q(\ram[108][14] ), 
	.D(FE_PHN2120_n2324), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[108][13]  (.Q(\ram[108][13] ), 
	.D(FE_PHN1624_n2323), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[108][12]  (.Q(\ram[108][12] ), 
	.D(FE_PHN2217_n2322), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][11]  (.Q(\ram[108][11] ), 
	.D(FE_PHN1507_n2321), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][10]  (.Q(\ram[108][10] ), 
	.D(FE_PHN2907_n2320), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[108][9]  (.Q(\ram[108][9] ), 
	.D(FE_PHN2183_n2319), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[108][8]  (.Q(\ram[108][8] ), 
	.D(FE_PHN2087_n2318), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][7]  (.Q(\ram[108][7] ), 
	.D(FE_PHN2875_n2317), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[108][6]  (.Q(\ram[108][6] ), 
	.D(FE_PHN1913_n2316), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][5]  (.Q(\ram[108][5] ), 
	.D(FE_PHN1457_n2315), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][4]  (.Q(\ram[108][4] ), 
	.D(FE_PHN2534_n2314), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[108][3]  (.Q(\ram[108][3] ), 
	.D(FE_PHN1600_n2313), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[108][2]  (.Q(\ram[108][2] ), 
	.D(FE_PHN897_n2312), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][1]  (.Q(\ram[108][1] ), 
	.D(FE_PHN1643_n2311), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[108][0]  (.Q(\ram[108][0] ), 
	.D(FE_PHN2883_n2310), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[104][15]  (.Q(\ram[104][15] ), 
	.D(FE_PHN2696_n2261), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][14]  (.Q(\ram[104][14] ), 
	.D(FE_PHN780_n2260), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][13]  (.Q(\ram[104][13] ), 
	.D(n2259), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][12]  (.Q(\ram[104][12] ), 
	.D(FE_PHN3972_n2258), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][11]  (.Q(\ram[104][11] ), 
	.D(FE_PHN5694_n2257), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][10]  (.Q(\ram[104][10] ), 
	.D(FE_PHN2740_n2256), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][9]  (.Q(\ram[104][9] ), 
	.D(FE_PHN1733_n2255), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][8]  (.Q(\ram[104][8] ), 
	.D(FE_PHN464_n2254), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[104][7]  (.Q(\ram[104][7] ), 
	.D(FE_PHN856_n2253), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[104][6]  (.Q(\ram[104][6] ), 
	.D(FE_PHN1999_n2252), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][5]  (.Q(\ram[104][5] ), 
	.D(FE_PHN5711_n2251), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[104][4]  (.Q(\ram[104][4] ), 
	.D(FE_PHN1290_n2250), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][3]  (.Q(\ram[104][3] ), 
	.D(FE_PHN2095_n2249), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][2]  (.Q(\ram[104][2] ), 
	.D(FE_PHN2678_n2248), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[104][1]  (.Q(\ram[104][1] ), 
	.D(FE_PHN2897_n2247), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[104][0]  (.Q(\ram[104][0] ), 
	.D(FE_PHN1631_n2246), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[100][15]  (.Q(\ram[100][15] ), 
	.D(FE_PHN896_n2197), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][14]  (.Q(\ram[100][14] ), 
	.D(FE_PHN3165_n2196), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][13]  (.Q(\ram[100][13] ), 
	.D(FE_PHN1086_n2195), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][12]  (.Q(\ram[100][12] ), 
	.D(FE_PHN1360_n2194), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][11]  (.Q(\ram[100][11] ), 
	.D(FE_PHN1091_n2193), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][10]  (.Q(\ram[100][10] ), 
	.D(FE_PHN1006_n2192), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][9]  (.Q(\ram[100][9] ), 
	.D(FE_PHN1663_n2191), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][8]  (.Q(\ram[100][8] ), 
	.D(FE_PHN1178_n2190), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[100][7]  (.Q(\ram[100][7] ), 
	.D(FE_PHN1068_n2189), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[100][6]  (.Q(\ram[100][6] ), 
	.D(FE_PHN1105_n2188), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][5]  (.Q(\ram[100][5] ), 
	.D(FE_PHN1535_n2187), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][4]  (.Q(\ram[100][4] ), 
	.D(FE_PHN2439_n2186), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][3]  (.Q(\ram[100][3] ), 
	.D(FE_PHN526_n2185), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[100][2]  (.Q(\ram[100][2] ), 
	.D(FE_PHN2518_n2184), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[100][1]  (.Q(\ram[100][1] ), 
	.D(FE_PHN544_n2183), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[100][0]  (.Q(\ram[100][0] ), 
	.D(FE_PHN1817_n2182), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[96][15]  (.Q(\ram[96][15] ), 
	.D(FE_PHN6711_n2133), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][14]  (.Q(\ram[96][14] ), 
	.D(FE_PHN6679_n2132), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][13]  (.Q(\ram[96][13] ), 
	.D(FE_PHN4471_n2131), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[96][12]  (.Q(\ram[96][12] ), 
	.D(FE_PHN4779_n2130), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[96][11]  (.Q(\ram[96][11] ), 
	.D(FE_PHN830_n2129), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[96][10]  (.Q(\ram[96][10] ), 
	.D(FE_PHN935_n2128), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][9]  (.Q(\ram[96][9] ), 
	.D(FE_PHN3371_n2127), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][8]  (.Q(\ram[96][8] ), 
	.D(FE_PHN6703_n2126), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[96][7]  (.Q(\ram[96][7] ), 
	.D(FE_PHN5724_n2125), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][6]  (.Q(\ram[96][6] ), 
	.D(FE_PHN5690_n2124), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[96][5]  (.Q(\ram[96][5] ), 
	.D(FE_PHN5658_n2123), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[96][4]  (.Q(\ram[96][4] ), 
	.D(FE_PHN5664_n2122), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[96][3]  (.Q(\ram[96][3] ), 
	.D(FE_PHN5657_n2121), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[96][2]  (.Q(\ram[96][2] ), 
	.D(FE_PHN6699_n2120), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[96][1]  (.Q(\ram[96][1] ), 
	.D(FE_PHN6671_n2119), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[96][0]  (.Q(\ram[96][0] ), 
	.D(FE_PHN7254_n2118), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[92][15]  (.Q(\ram[92][15] ), 
	.D(FE_PHN2668_n2069), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[92][14]  (.Q(\ram[92][14] ), 
	.D(FE_PHN2708_n2068), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][13]  (.Q(\ram[92][13] ), 
	.D(FE_PHN2578_n2067), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][12]  (.Q(\ram[92][12] ), 
	.D(FE_PHN2726_n2066), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][11]  (.Q(\ram[92][11] ), 
	.D(FE_PHN2893_n2065), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][10]  (.Q(\ram[92][10] ), 
	.D(FE_PHN1945_n2064), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][9]  (.Q(\ram[92][9] ), 
	.D(FE_PHN2426_n2063), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][8]  (.Q(\ram[92][8] ), 
	.D(FE_PHN2092_n2062), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[92][7]  (.Q(\ram[92][7] ), 
	.D(FE_PHN2222_n2061), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[92][6]  (.Q(\ram[92][6] ), 
	.D(FE_PHN2944_n2060), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][5]  (.Q(\ram[92][5] ), 
	.D(FE_PHN2686_n2059), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[92][4]  (.Q(\ram[92][4] ), 
	.D(FE_PHN1972_n2058), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[92][3]  (.Q(\ram[92][3] ), 
	.D(FE_PHN2629_n2057), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[92][2]  (.Q(\ram[92][2] ), 
	.D(FE_PHN2061_n2056), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[92][1]  (.Q(\ram[92][1] ), 
	.D(FE_PHN3026_n2055), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[92][0]  (.Q(\ram[92][0] ), 
	.D(FE_PHN2665_n2054), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[88][15]  (.Q(\ram[88][15] ), 
	.D(FE_PHN3226_n2005), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[88][14]  (.Q(\ram[88][14] ), 
	.D(FE_PHN2754_n2004), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[88][13]  (.Q(\ram[88][13] ), 
	.D(FE_PHN2760_n2003), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[88][12]  (.Q(\ram[88][12] ), 
	.D(FE_PHN2731_n2002), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[88][11]  (.Q(\ram[88][11] ), 
	.D(FE_PHN2886_n2001), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[88][10]  (.Q(\ram[88][10] ), 
	.D(FE_PHN1739_n2000), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[88][9]  (.Q(\ram[88][9] ), 
	.D(FE_PHN1969_n1999), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[88][8]  (.Q(\ram[88][8] ), 
	.D(FE_PHN2000_n1998), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][7]  (.Q(\ram[88][7] ), 
	.D(FE_PHN2389_n1997), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[88][6]  (.Q(\ram[88][6] ), 
	.D(FE_PHN2577_n1996), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][5]  (.Q(\ram[88][5] ), 
	.D(FE_PHN2051_n1995), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][4]  (.Q(\ram[88][4] ), 
	.D(FE_PHN2422_n1994), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[88][3]  (.Q(\ram[88][3] ), 
	.D(FE_PHN3187_n1993), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][2]  (.Q(\ram[88][2] ), 
	.D(FE_PHN2471_n1992), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[88][1]  (.Q(\ram[88][1] ), 
	.D(FE_PHN2593_n1991), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[88][0]  (.Q(\ram[88][0] ), 
	.D(FE_PHN2066_n1990), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[84][15]  (.Q(\ram[84][15] ), 
	.D(FE_PHN3022_n1941), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][14]  (.Q(\ram[84][14] ), 
	.D(FE_PHN2746_n1940), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][13]  (.Q(\ram[84][13] ), 
	.D(FE_PHN1666_n1939), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[84][12]  (.Q(\ram[84][12] ), 
	.D(FE_PHN2600_n1938), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[84][11]  (.Q(\ram[84][11] ), 
	.D(FE_PHN3143_n1937), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][10]  (.Q(\ram[84][10] ), 
	.D(FE_PHN2456_n1936), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[84][9]  (.Q(\ram[84][9] ), 
	.D(FE_PHN3087_n1935), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[84][8]  (.Q(\ram[84][8] ), 
	.D(FE_PHN2552_n1934), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[84][7]  (.Q(\ram[84][7] ), 
	.D(FE_PHN1867_n1933), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[84][6]  (.Q(\ram[84][6] ), 
	.D(FE_PHN1609_n1932), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][5]  (.Q(\ram[84][5] ), 
	.D(FE_PHN2707_n1931), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[84][4]  (.Q(\ram[84][4] ), 
	.D(FE_PHN1283_n1930), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][3]  (.Q(\ram[84][3] ), 
	.D(FE_PHN2507_n1929), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][2]  (.Q(\ram[84][2] ), 
	.D(FE_PHN1943_n1928), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[84][1]  (.Q(\ram[84][1] ), 
	.D(FE_PHN2664_n1927), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[84][0]  (.Q(\ram[84][0] ), 
	.D(FE_PHN2245_n1926), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[80][15]  (.Q(\ram[80][15] ), 
	.D(FE_PHN1126_n1877), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][14]  (.Q(\ram[80][14] ), 
	.D(FE_PHN2378_n1876), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][13]  (.Q(\ram[80][13] ), 
	.D(FE_PHN2613_n1875), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][12]  (.Q(\ram[80][12] ), 
	.D(FE_PHN4609_n1874), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][11]  (.Q(\ram[80][11] ), 
	.D(FE_PHN4251_n1873), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][10]  (.Q(\ram[80][10] ), 
	.D(FE_PHN4538_n1872), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[80][9]  (.Q(\ram[80][9] ), 
	.D(FE_PHN1364_n1871), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[80][8]  (.Q(\ram[80][8] ), 
	.D(FE_PHN4626_n1870), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[80][7]  (.Q(\ram[80][7] ), 
	.D(FE_PHN1698_n1869), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[80][6]  (.Q(\ram[80][6] ), 
	.D(FE_PHN2673_n1868), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][5]  (.Q(\ram[80][5] ), 
	.D(FE_PHN1226_n1867), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][4]  (.Q(\ram[80][4] ), 
	.D(FE_PHN2782_n1866), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][3]  (.Q(\ram[80][3] ), 
	.D(FE_PHN5757_n1865), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[80][2]  (.Q(\ram[80][2] ), 
	.D(FE_PHN4218_n1864), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[80][1]  (.Q(\ram[80][1] ), 
	.D(FE_PHN6674_n1863), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[80][0]  (.Q(\ram[80][0] ), 
	.D(FE_PHN1191_n1862), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[76][15]  (.Q(\ram[76][15] ), 
	.D(FE_PHN393_n1813), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][14]  (.Q(\ram[76][14] ), 
	.D(FE_PHN1480_n1812), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[76][13]  (.Q(\ram[76][13] ), 
	.D(FE_PHN885_n1811), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[76][12]  (.Q(\ram[76][12] ), 
	.D(FE_PHN1819_n1810), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[76][11]  (.Q(\ram[76][11] ), 
	.D(FE_PHN998_n1809), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][10]  (.Q(\ram[76][10] ), 
	.D(FE_PHN2595_n1808), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][9]  (.Q(\ram[76][9] ), 
	.D(FE_PHN2918_n1807), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][8]  (.Q(\ram[76][8] ), 
	.D(FE_PHN2890_n1806), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[76][7]  (.Q(\ram[76][7] ), 
	.D(FE_PHN1351_n1805), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[76][6]  (.Q(\ram[76][6] ), 
	.D(FE_PHN3141_n1804), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][5]  (.Q(\ram[76][5] ), 
	.D(FE_PHN1553_n1803), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[76][4]  (.Q(\ram[76][4] ), 
	.D(FE_PHN417_n1802), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][3]  (.Q(\ram[76][3] ), 
	.D(FE_PHN873_n1801), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][2]  (.Q(\ram[76][2] ), 
	.D(FE_PHN845_n1800), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[76][1]  (.Q(\ram[76][1] ), 
	.D(FE_PHN3185_n1799), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[76][0]  (.Q(\ram[76][0] ), 
	.D(FE_PHN630_n1798), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[72][15]  (.Q(\ram[72][15] ), 
	.D(FE_PHN2131_n1749), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][14]  (.Q(\ram[72][14] ), 
	.D(FE_PHN2898_n1748), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][13]  (.Q(\ram[72][13] ), 
	.D(FE_PHN2812_n1747), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[72][12]  (.Q(\ram[72][12] ), 
	.D(FE_PHN1661_n1746), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][11]  (.Q(\ram[72][11] ), 
	.D(FE_PHN915_n1745), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][10]  (.Q(\ram[72][10] ), 
	.D(FE_PHN2643_n1744), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][9]  (.Q(\ram[72][9] ), 
	.D(FE_PHN1606_n1743), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][8]  (.Q(\ram[72][8] ), 
	.D(FE_PHN1069_n1742), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[72][7]  (.Q(\ram[72][7] ), 
	.D(FE_PHN3105_n1741), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][6]  (.Q(\ram[72][6] ), 
	.D(FE_PHN659_n1740), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[72][5]  (.Q(\ram[72][5] ), 
	.D(FE_PHN2712_n1739), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][4]  (.Q(\ram[72][4] ), 
	.D(FE_PHN1822_n1738), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][3]  (.Q(\ram[72][3] ), 
	.D(FE_PHN3126_n1737), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[72][2]  (.Q(\ram[72][2] ), 
	.D(FE_PHN2023_n1736), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][1]  (.Q(\ram[72][1] ), 
	.D(FE_PHN538_n1735), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[72][0]  (.Q(\ram[72][0] ), 
	.D(FE_PHN2416_n1734), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[68][15]  (.Q(\ram[68][15] ), 
	.D(FE_PHN1200_n1685), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][14]  (.Q(\ram[68][14] ), 
	.D(FE_PHN2270_n1684), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][13]  (.Q(\ram[68][13] ), 
	.D(FE_PHN799_n1683), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][12]  (.Q(\ram[68][12] ), 
	.D(FE_PHN1645_n1682), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][11]  (.Q(\ram[68][11] ), 
	.D(FE_PHN3075_n1681), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][10]  (.Q(\ram[68][10] ), 
	.D(FE_PHN744_n1680), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][9]  (.Q(\ram[68][9] ), 
	.D(FE_PHN1893_n1679), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][8]  (.Q(\ram[68][8] ), 
	.D(FE_PHN1931_n1678), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][7]  (.Q(\ram[68][7] ), 
	.D(FE_PHN2220_n1677), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[68][6]  (.Q(\ram[68][6] ), 
	.D(FE_PHN3144_n1676), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][5]  (.Q(\ram[68][5] ), 
	.D(FE_PHN907_n1675), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][4]  (.Q(\ram[68][4] ), 
	.D(FE_PHN2557_n1674), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][3]  (.Q(\ram[68][3] ), 
	.D(FE_PHN1120_n1673), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[68][2]  (.Q(\ram[68][2] ), 
	.D(FE_PHN2648_n1672), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[68][1]  (.Q(\ram[68][1] ), 
	.D(FE_PHN2380_n1671), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[68][0]  (.Q(\ram[68][0] ), 
	.D(FE_PHN1205_n1670), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[64][15]  (.Q(\ram[64][15] ), 
	.D(FE_PHN1115_n1621), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][14]  (.Q(\ram[64][14] ), 
	.D(FE_PHN1981_n1620), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][13]  (.Q(\ram[64][13] ), 
	.D(FE_PHN2626_n1619), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[64][12]  (.Q(\ram[64][12] ), 
	.D(FE_PHN3042_n1618), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[64][11]  (.Q(\ram[64][11] ), 
	.D(FE_PHN2145_n1617), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][10]  (.Q(\ram[64][10] ), 
	.D(FE_PHN566_n1616), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][9]  (.Q(\ram[64][9] ), 
	.D(FE_PHN3059_n1615), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[64][8]  (.Q(\ram[64][8] ), 
	.D(FE_PHN2436_n1614), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][7]  (.Q(\ram[64][7] ), 
	.D(FE_PHN3029_n1613), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[64][6]  (.Q(\ram[64][6] ), 
	.D(FE_PHN797_n1612), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][5]  (.Q(\ram[64][5] ), 
	.D(FE_PHN536_n1611), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][4]  (.Q(\ram[64][4] ), 
	.D(FE_PHN2167_n1610), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][3]  (.Q(\ram[64][3] ), 
	.D(FE_PHN2982_n1609), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][2]  (.Q(\ram[64][2] ), 
	.D(FE_PHN716_n1608), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[64][1]  (.Q(\ram[64][1] ), 
	.D(FE_PHN1275_n1607), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[64][0]  (.Q(\ram[64][0] ), 
	.D(FE_PHN2137_n1606), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[60][15]  (.Q(\ram[60][15] ), 
	.D(FE_PHN2124_n1557), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][14]  (.Q(\ram[60][14] ), 
	.D(FE_PHN1511_n1556), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][13]  (.Q(\ram[60][13] ), 
	.D(FE_PHN2649_n1555), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[60][12]  (.Q(\ram[60][12] ), 
	.D(FE_PHN1107_n1554), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][11]  (.Q(\ram[60][11] ), 
	.D(FE_PHN2993_n1553), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][10]  (.Q(\ram[60][10] ), 
	.D(FE_PHN1618_n1552), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][9]  (.Q(\ram[60][9] ), 
	.D(FE_PHN2554_n1551), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[60][8]  (.Q(\ram[60][8] ), 
	.D(FE_PHN1269_n1550), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[60][7]  (.Q(\ram[60][7] ), 
	.D(FE_PHN1736_n1549), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[60][6]  (.Q(\ram[60][6] ), 
	.D(FE_PHN1547_n1548), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][5]  (.Q(\ram[60][5] ), 
	.D(FE_PHN611_n1547), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][4]  (.Q(\ram[60][4] ), 
	.D(FE_PHN2688_n1546), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][3]  (.Q(\ram[60][3] ), 
	.D(FE_PHN2887_n1545), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[60][2]  (.Q(\ram[60][2] ), 
	.D(FE_PHN1619_n1544), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[60][1]  (.Q(\ram[60][1] ), 
	.D(FE_PHN3048_n1543), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[60][0]  (.Q(\ram[60][0] ), 
	.D(FE_PHN1527_n1542), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[56][15]  (.Q(\ram[56][15] ), 
	.D(FE_PHN631_n1493), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[56][14]  (.Q(\ram[56][14] ), 
	.D(FE_PHN2776_n1492), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[56][13]  (.Q(\ram[56][13] ), 
	.D(FE_PHN3054_n1491), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][12]  (.Q(\ram[56][12] ), 
	.D(FE_PHN1556_n1490), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[56][11]  (.Q(\ram[56][11] ), 
	.D(FE_PHN3230_n1489), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][10]  (.Q(\ram[56][10] ), 
	.D(FE_PHN2899_n1488), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][9]  (.Q(\ram[56][9] ), 
	.D(FE_PHN2925_n1487), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[56][8]  (.Q(\ram[56][8] ), 
	.D(FE_PHN2417_n1486), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[56][7]  (.Q(\ram[56][7] ), 
	.D(FE_PHN1571_n1485), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][6]  (.Q(\ram[56][6] ), 
	.D(FE_PHN3067_n1484), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[56][5]  (.Q(\ram[56][5] ), 
	.D(FE_PHN2636_n1483), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][4]  (.Q(\ram[56][4] ), 
	.D(FE_PHN2259_n1482), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[56][3]  (.Q(\ram[56][3] ), 
	.D(FE_PHN2768_n1481), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[56][2]  (.Q(\ram[56][2] ), 
	.D(FE_PHN693_n1480), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[56][1]  (.Q(\ram[56][1] ), 
	.D(FE_PHN831_n1479), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[56][0]  (.Q(\ram[56][0] ), 
	.D(FE_PHN1540_n1478), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[52][15]  (.Q(\ram[52][15] ), 
	.D(n1429), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][14]  (.Q(\ram[52][14] ), 
	.D(FE_PHN2624_n1428), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][13]  (.Q(\ram[52][13] ), 
	.D(FE_PHN2330_n1427), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][12]  (.Q(\ram[52][12] ), 
	.D(FE_PHN3078_n1426), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][11]  (.Q(\ram[52][11] ), 
	.D(FE_PHN3216_n1425), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][10]  (.Q(\ram[52][10] ), 
	.D(FE_PHN2074_n1424), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][9]  (.Q(\ram[52][9] ), 
	.D(FE_PHN1433_n1423), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[52][8]  (.Q(\ram[52][8] ), 
	.D(FE_PHN3211_n1422), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][7]  (.Q(\ram[52][7] ), 
	.D(FE_PHN2608_n1421), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][6]  (.Q(\ram[52][6] ), 
	.D(FE_PHN2872_n1420), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][5]  (.Q(\ram[52][5] ), 
	.D(FE_PHN3041_n1419), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][4]  (.Q(\ram[52][4] ), 
	.D(FE_PHN1941_n1418), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][3]  (.Q(\ram[52][3] ), 
	.D(FE_PHN3014_n1417), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[52][2]  (.Q(\ram[52][2] ), 
	.D(FE_PHN2493_n1416), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][1]  (.Q(\ram[52][1] ), 
	.D(FE_PHN2041_n1415), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[52][0]  (.Q(\ram[52][0] ), 
	.D(FE_PHN2067_n1414), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[48][15]  (.Q(\ram[48][15] ), 
	.D(FE_PHN2771_n1365), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[48][14]  (.Q(\ram[48][14] ), 
	.D(FE_PHN1327_n1364), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[48][13]  (.Q(\ram[48][13] ), 
	.D(FE_PHN2830_n1363), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][12]  (.Q(\ram[48][12] ), 
	.D(FE_PHN2244_n1362), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][11]  (.Q(\ram[48][11] ), 
	.D(FE_PHN3010_n1361), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][10]  (.Q(\ram[48][10] ), 
	.D(FE_PHN1074_n1360), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][9]  (.Q(\ram[48][9] ), 
	.D(FE_PHN2681_n1359), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[48][8]  (.Q(\ram[48][8] ), 
	.D(FE_PHN3106_n1358), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[48][7]  (.Q(\ram[48][7] ), 
	.D(FE_PHN2226_n1357), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[48][6]  (.Q(\ram[48][6] ), 
	.D(FE_PHN2384_n1356), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[48][5]  (.Q(\ram[48][5] ), 
	.D(FE_PHN3109_n1355), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][4]  (.Q(\ram[48][4] ), 
	.D(FE_PHN3132_n1354), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][3]  (.Q(\ram[48][3] ), 
	.D(FE_PHN1528_n1353), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[48][2]  (.Q(\ram[48][2] ), 
	.D(FE_PHN2437_n1352), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[48][1]  (.Q(\ram[48][1] ), 
	.D(FE_PHN978_n1351), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[48][0]  (.Q(\ram[48][0] ), 
	.D(FE_PHN2987_n1350), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[44][15]  (.Q(\ram[44][15] ), 
	.D(FE_PHN3028_n1301), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[44][14]  (.Q(\ram[44][14] ), 
	.D(FE_PHN1617_n1300), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][13]  (.Q(\ram[44][13] ), 
	.D(FE_PHN2026_n1299), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[44][12]  (.Q(\ram[44][12] ), 
	.D(FE_PHN712_n1298), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[44][11]  (.Q(\ram[44][11] ), 
	.D(FE_PHN2136_n1297), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][10]  (.Q(\ram[44][10] ), 
	.D(FE_PHN2781_n1296), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[44][9]  (.Q(\ram[44][9] ), 
	.D(FE_PHN1725_n1295), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[44][8]  (.Q(\ram[44][8] ), 
	.D(FE_PHN2279_n1294), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[44][7]  (.Q(\ram[44][7] ), 
	.D(FE_PHN2804_n1293), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[44][6]  (.Q(\ram[44][6] ), 
	.D(FE_PHN2179_n1292), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][5]  (.Q(\ram[44][5] ), 
	.D(FE_PHN2197_n1291), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][4]  (.Q(\ram[44][4] ), 
	.D(FE_PHN2825_n1290), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][3]  (.Q(\ram[44][3] ), 
	.D(FE_PHN3007_n1289), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[44][2]  (.Q(\ram[44][2] ), 
	.D(FE_PHN1607_n1288), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][1]  (.Q(\ram[44][1] ), 
	.D(FE_PHN2566_n1287), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[44][0]  (.Q(\ram[44][0] ), 
	.D(FE_PHN5660_n1286), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[40][15]  (.Q(\ram[40][15] ), 
	.D(FE_PHN1918_n1237), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][14]  (.Q(\ram[40][14] ), 
	.D(FE_PHN3151_n1236), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][13]  (.Q(\ram[40][13] ), 
	.D(FE_PHN2420_n1235), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][12]  (.Q(\ram[40][12] ), 
	.D(FE_PHN1864_n1234), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[40][11]  (.Q(\ram[40][11] ), 
	.D(FE_PHN1273_n1233), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[40][10]  (.Q(\ram[40][10] ), 
	.D(FE_PHN2097_n1232), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][9]  (.Q(\ram[40][9] ), 
	.D(FE_PHN1186_n1231), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][8]  (.Q(\ram[40][8] ), 
	.D(FE_PHN1620_n1230), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[40][7]  (.Q(\ram[40][7] ), 
	.D(FE_PHN3070_n1229), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[40][6]  (.Q(\ram[40][6] ), 
	.D(FE_PHN2858_n1228), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[40][5]  (.Q(\ram[40][5] ), 
	.D(FE_PHN1625_n1227), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[40][4]  (.Q(\ram[40][4] ), 
	.D(FE_PHN1726_n1226), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][3]  (.Q(\ram[40][3] ), 
	.D(FE_PHN2902_n1225), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[40][2]  (.Q(\ram[40][2] ), 
	.D(FE_PHN2254_n1224), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][1]  (.Q(\ram[40][1] ), 
	.D(FE_PHN2277_n1223), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[40][0]  (.Q(\ram[40][0] ), 
	.D(FE_PHN2859_n1222), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[36][15]  (.Q(\ram[36][15] ), 
	.D(FE_PHN1794_n1173), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][14]  (.Q(\ram[36][14] ), 
	.D(FE_PHN1588_n1172), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[36][13]  (.Q(\ram[36][13] ), 
	.D(FE_PHN2470_n1171), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[36][12]  (.Q(\ram[36][12] ), 
	.D(FE_PHN835_n1170), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[36][11]  (.Q(\ram[36][11] ), 
	.D(FE_PHN2075_n1169), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][10]  (.Q(\ram[36][10] ), 
	.D(FE_PHN2084_n1168), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][9]  (.Q(\ram[36][9] ), 
	.D(FE_PHN2481_n1167), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][8]  (.Q(\ram[36][8] ), 
	.D(FE_PHN3083_n1166), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][7]  (.Q(\ram[36][7] ), 
	.D(FE_PHN932_n1165), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][6]  (.Q(\ram[36][6] ), 
	.D(FE_PHN2966_n1164), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][5]  (.Q(\ram[36][5] ), 
	.D(FE_PHN3080_n1163), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[36][4]  (.Q(\ram[36][4] ), 
	.D(FE_PHN2814_n1162), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[36][3]  (.Q(\ram[36][3] ), 
	.D(FE_PHN3064_n1161), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[36][2]  (.Q(\ram[36][2] ), 
	.D(FE_PHN614_n1160), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[36][1]  (.Q(\ram[36][1] ), 
	.D(FE_PHN1987_n1159), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[36][0]  (.Q(\ram[36][0] ), 
	.D(FE_PHN4836_n1158), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[32][15]  (.Q(\ram[32][15] ), 
	.D(FE_PHN2732_n1109), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][14]  (.Q(\ram[32][14] ), 
	.D(FE_PHN2106_n1108), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][13]  (.Q(\ram[32][13] ), 
	.D(FE_PHN2879_n1107), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][12]  (.Q(\ram[32][12] ), 
	.D(FE_PHN3715_n1106), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[32][11]  (.Q(\ram[32][11] ), 
	.D(FE_PHN750_n1105), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][10]  (.Q(\ram[32][10] ), 
	.D(FE_PHN3098_n1104), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[32][9]  (.Q(\ram[32][9] ), 
	.D(FE_PHN2971_n1103), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][8]  (.Q(\ram[32][8] ), 
	.D(FE_PHN1063_n1102), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][7]  (.Q(\ram[32][7] ), 
	.D(FE_PHN3065_n1101), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[32][6]  (.Q(\ram[32][6] ), 
	.D(FE_PHN899_n1100), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][5]  (.Q(\ram[32][5] ), 
	.D(FE_PHN3222_n1099), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][4]  (.Q(\ram[32][4] ), 
	.D(FE_PHN1649_n1098), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][3]  (.Q(\ram[32][3] ), 
	.D(FE_PHN2717_n1097), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[32][2]  (.Q(\ram[32][2] ), 
	.D(FE_PHN2264_n1096), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[32][1]  (.Q(\ram[32][1] ), 
	.D(FE_PHN2141_n1095), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[32][0]  (.Q(\ram[32][0] ), 
	.D(FE_PHN5729_n1094), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[28][15]  (.Q(\ram[28][15] ), 
	.D(FE_PHN4067_n1045), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[28][14]  (.Q(\ram[28][14] ), 
	.D(FE_PHN2553_n1044), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[28][13]  (.Q(\ram[28][13] ), 
	.D(FE_PHN3127_n1043), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[28][12]  (.Q(\ram[28][12] ), 
	.D(FE_PHN5444_n1042), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[28][11]  (.Q(\ram[28][11] ), 
	.D(FE_PHN1920_n1041), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][10]  (.Q(\ram[28][10] ), 
	.D(FE_PHN4182_n1040), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[28][9]  (.Q(\ram[28][9] ), 
	.D(FE_PHN1812_n1039), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[28][8]  (.Q(\ram[28][8] ), 
	.D(FE_PHN5143_n1038), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][7]  (.Q(\ram[28][7] ), 
	.D(FE_PHN4537_n1037), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[28][6]  (.Q(\ram[28][6] ), 
	.D(FE_PHN2219_n1036), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[28][5]  (.Q(\ram[28][5] ), 
	.D(FE_PHN648_n1035), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][4]  (.Q(\ram[28][4] ), 
	.D(FE_PHN5078_n1034), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[28][3]  (.Q(\ram[28][3] ), 
	.D(FE_PHN2178_n1033), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[28][2]  (.Q(\ram[28][2] ), 
	.D(FE_PHN4271_n1032), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[28][1]  (.Q(\ram[28][1] ), 
	.D(FE_PHN5717_n1031), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[28][0]  (.Q(\ram[28][0] ), 
	.D(FE_PHN4428_n1030), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[24][15]  (.Q(\ram[24][15] ), 
	.D(FE_PHN4904_n981), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][14]  (.Q(\ram[24][14] ), 
	.D(FE_PHN5696_n980), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][13]  (.Q(\ram[24][13] ), 
	.D(FE_PHN5669_n979), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[24][12]  (.Q(\ram[24][12] ), 
	.D(FE_PHN4241_n978), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[24][11]  (.Q(\ram[24][11] ), 
	.D(FE_PHN5725_n977), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[24][10]  (.Q(\ram[24][10] ), 
	.D(FE_PHN4399_n976), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[24][9]  (.Q(\ram[24][9] ), 
	.D(FE_PHN3527_n975), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[24][8]  (.Q(\ram[24][8] ), 
	.D(FE_PHN3391_n974), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][7]  (.Q(\ram[24][7] ), 
	.D(FE_PHN5745_n973), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][6]  (.Q(\ram[24][6] ), 
	.D(FE_PHN4542_n972), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[24][5]  (.Q(\ram[24][5] ), 
	.D(FE_PHN3506_n971), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[24][4]  (.Q(\ram[24][4] ), 
	.D(FE_PHN4027_n970), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[24][3]  (.Q(\ram[24][3] ), 
	.D(FE_PHN4622_n969), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][2]  (.Q(\ram[24][2] ), 
	.D(FE_PHN4545_n968), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[24][1]  (.Q(\ram[24][1] ), 
	.D(FE_PHN5677_n967), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[24][0]  (.Q(\ram[24][0] ), 
	.D(FE_PHN3956_n966), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[20][15]  (.Q(\ram[20][15] ), 
	.D(FE_PHN4508_n917), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][14]  (.Q(\ram[20][14] ), 
	.D(FE_PHN2634_n916), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][13]  (.Q(\ram[20][13] ), 
	.D(FE_PHN336_n915), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][12]  (.Q(\ram[20][12] ), 
	.D(FE_PHN4082_n914), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][11]  (.Q(\ram[20][11] ), 
	.D(FE_PHN4560_n913), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][10]  (.Q(\ram[20][10] ), 
	.D(n912), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[20][9]  (.Q(\ram[20][9] ), 
	.D(FE_PHN4681_n911), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][8]  (.Q(\ram[20][8] ), 
	.D(FE_PHN4593_n910), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][7]  (.Q(\ram[20][7] ), 
	.D(FE_PHN5555_n909), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][6]  (.Q(\ram[20][6] ), 
	.D(FE_PHN1082_n908), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[20][5]  (.Q(\ram[20][5] ), 
	.D(FE_PHN3088_n907), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[20][4]  (.Q(\ram[20][4] ), 
	.D(FE_PHN4361_n906), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[20][3]  (.Q(\ram[20][3] ), 
	.D(FE_PHN4557_n905), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][2]  (.Q(\ram[20][2] ), 
	.D(FE_PHN5033_n904), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[20][1]  (.Q(\ram[20][1] ), 
	.D(FE_PHN4667_n903), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[20][0]  (.Q(\ram[20][0] ), 
	.D(FE_PHN3865_n902), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[16][15]  (.Q(\ram[16][15] ), 
	.D(FE_PHN4331_n853), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[16][14]  (.Q(\ram[16][14] ), 
	.D(FE_PHN4261_n852), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][13]  (.Q(\ram[16][13] ), 
	.D(FE_PHN4333_n851), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[16][12]  (.Q(\ram[16][12] ), 
	.D(FE_PHN4647_n850), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[16][11]  (.Q(\ram[16][11] ), 
	.D(FE_PHN4491_n849), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][10]  (.Q(\ram[16][10] ), 
	.D(FE_PHN4221_n848), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][9]  (.Q(\ram[16][9] ), 
	.D(FE_PHN4588_n847), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][8]  (.Q(\ram[16][8] ), 
	.D(FE_PHN4267_n846), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][7]  (.Q(\ram[16][7] ), 
	.D(FE_PHN5494_n845), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[16][6]  (.Q(\ram[16][6] ), 
	.D(FE_PHN3863_n844), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[16][5]  (.Q(\ram[16][5] ), 
	.D(FE_PHN4696_n843), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[16][4]  (.Q(\ram[16][4] ), 
	.D(FE_PHN4217_n842), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[16][3]  (.Q(\ram[16][3] ), 
	.D(FE_PHN4605_n841), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[16][2]  (.Q(\ram[16][2] ), 
	.D(FE_PHN4324_n840), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[16][1]  (.Q(\ram[16][1] ), 
	.D(FE_PHN4698_n839), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[16][0]  (.Q(\ram[16][0] ), 
	.D(FE_PHN4722_n838), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[12][15]  (.Q(\ram[12][15] ), 
	.D(FE_PHN2353_n789), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[12][14]  (.Q(\ram[12][14] ), 
	.D(FE_PHN1454_n788), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[12][13]  (.Q(\ram[12][13] ), 
	.D(FE_PHN1872_n787), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][12]  (.Q(\ram[12][12] ), 
	.D(FE_PHN1587_n786), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[12][11]  (.Q(\ram[12][11] ), 
	.D(FE_PHN2998_n785), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][10]  (.Q(\ram[12][10] ), 
	.D(FE_PHN1064_n784), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[12][9]  (.Q(\ram[12][9] ), 
	.D(FE_PHN2170_n783), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][8]  (.Q(\ram[12][8] ), 
	.D(FE_PHN2573_n782), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][7]  (.Q(\ram[12][7] ), 
	.D(FE_PHN3114_n781), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][6]  (.Q(\ram[12][6] ), 
	.D(FE_PHN1482_n780), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][5]  (.Q(\ram[12][5] ), 
	.D(FE_PHN941_n779), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][4]  (.Q(\ram[12][4] ), 
	.D(FE_PHN2744_n778), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][3]  (.Q(\ram[12][3] ), 
	.D(FE_PHN2382_n777), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[12][2]  (.Q(\ram[12][2] ), 
	.D(FE_PHN1573_n776), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[12][1]  (.Q(\ram[12][1] ), 
	.D(FE_PHN874_n775), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[12][0]  (.Q(\ram[12][0] ), 
	.D(FE_PHN1399_n774), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[8][15]  (.Q(\ram[8][15] ), 
	.D(FE_PHN2135_n725), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[8][14]  (.Q(\ram[8][14] ), 
	.D(FE_PHN2465_n724), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[8][13]  (.Q(\ram[8][13] ), 
	.D(FE_PHN848_n723), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[8][12]  (.Q(\ram[8][12] ), 
	.D(FE_PHN1934_n722), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[8][11]  (.Q(\ram[8][11] ), 
	.D(FE_PHN3036_n721), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][10]  (.Q(\ram[8][10] ), 
	.D(FE_PHN1954_n720), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[8][9]  (.Q(\ram[8][9] ), 
	.D(FE_PHN2821_n719), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][8]  (.Q(\ram[8][8] ), 
	.D(FE_PHN1940_n718), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[8][7]  (.Q(\ram[8][7] ), 
	.D(FE_PHN3179_n717), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[8][6]  (.Q(\ram[8][6] ), 
	.D(FE_PHN2223_n716), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[8][5]  (.Q(\ram[8][5] ), 
	.D(FE_PHN3133_n715), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][4]  (.Q(\ram[8][4] ), 
	.D(FE_PHN1952_n714), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[8][3]  (.Q(\ram[8][3] ), 
	.D(FE_PHN3224_n713), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[8][2]  (.Q(\ram[8][2] ), 
	.D(FE_PHN1432_n712), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[8][1]  (.Q(\ram[8][1] ), 
	.D(FE_PHN2803_n711), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[8][0]  (.Q(\ram[8][0] ), 
	.D(FE_PHN2797_n710), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[4][15]  (.Q(\ram[4][15] ), 
	.D(FE_PHN2037_n661), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[4][14]  (.Q(\ram[4][14] ), 
	.D(FE_PHN1530_n660), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[4][13]  (.Q(\ram[4][13] ), 
	.D(FE_PHN1288_n659), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[4][12]  (.Q(\ram[4][12] ), 
	.D(FE_PHN2848_n658), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[4][11]  (.Q(\ram[4][11] ), 
	.D(FE_PHN2885_n657), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][10]  (.Q(\ram[4][10] ), 
	.D(FE_PHN2076_n656), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[4][9]  (.Q(\ram[4][9] ), 
	.D(FE_PHN2951_n655), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[4][8]  (.Q(\ram[4][8] ), 
	.D(FE_PHN2205_n654), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[4][7]  (.Q(\ram[4][7] ), 
	.D(FE_PHN2837_n653), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[4][6]  (.Q(\ram[4][6] ), 
	.D(FE_PHN2824_n652), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][5]  (.Q(\ram[4][5] ), 
	.D(FE_PHN3150_n651), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][4]  (.Q(\ram[4][4] ), 
	.D(FE_PHN2878_n650), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[4][3]  (.Q(\ram[4][3] ), 
	.D(FE_PHN3227_n649), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[4][2]  (.Q(\ram[4][2] ), 
	.D(FE_PHN2003_n648), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[4][1]  (.Q(\ram[4][1] ), 
	.D(FE_PHN1568_n647), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[4][0]  (.Q(\ram[4][0] ), 
	.D(FE_PHN2325_n646), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[0][15]  (.Q(\ram[0][15] ), 
	.D(FE_PHN2010_n597), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][14]  (.Q(\ram[0][14] ), 
	.D(FE_PHN3052_n596), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][13]  (.Q(\ram[0][13] ), 
	.D(FE_PHN2386_n595), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[0][12]  (.Q(\ram[0][12] ), 
	.D(FE_PHN3164_n594), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[0][11]  (.Q(\ram[0][11] ), 
	.D(FE_PHN2709_n593), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[0][10]  (.Q(\ram[0][10] ), 
	.D(FE_PHN3180_n592), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[0][9]  (.Q(\ram[0][9] ), 
	.D(FE_PHN1744_n591), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[0][8]  (.Q(\ram[0][8] ), 
	.D(FE_PHN3204_n590), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][7]  (.Q(\ram[0][7] ), 
	.D(FE_PHN2253_n589), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[0][6]  (.Q(\ram[0][6] ), 
	.D(FE_PHN2983_n588), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[0][5]  (.Q(\ram[0][5] ), 
	.D(FE_PHN1493_n587), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[0][4]  (.Q(\ram[0][4] ), 
	.D(FE_PHN2243_n586), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[0][3]  (.Q(\ram[0][3] ), 
	.D(FE_PHN3037_n585), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[0][2]  (.Q(\ram[0][2] ), 
	.D(FE_PHN2679_n584), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[0][1]  (.Q(\ram[0][1] ), 
	.D(FE_PHN2984_n583), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[0][0]  (.Q(\ram[0][0] ), 
	.D(FE_PHN1576_n582), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[255][15]  (.Q(\ram[255][15] ), 
	.D(FE_PHN1685_n4677), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[255][14]  (.Q(\ram[255][14] ), 
	.D(FE_PHN958_n4676), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[255][13]  (.Q(\ram[255][13] ), 
	.D(FE_PHN2435_n4675), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][12]  (.Q(\ram[255][12] ), 
	.D(FE_PHN1847_n4674), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[255][11]  (.Q(\ram[255][11] ), 
	.D(FE_PHN1134_n4673), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[255][10]  (.Q(\ram[255][10] ), 
	.D(FE_PHN1012_n4672), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][9]  (.Q(\ram[255][9] ), 
	.D(FE_PHN2144_n4671), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][8]  (.Q(\ram[255][8] ), 
	.D(FE_PHN3021_n4670), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][7]  (.Q(\ram[255][7] ), 
	.D(FE_PHN680_n4669), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[255][6]  (.Q(\ram[255][6] ), 
	.D(FE_PHN694_n4668), 
	.CK(clk));
   QDFFEHD \ram_reg[255][5]  (.Q(\ram[255][5] ), 
	.D(FE_PHN2942_n4667), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[255][4]  (.Q(\ram[255][4] ), 
	.D(FE_PHN1077_n4666), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[255][3]  (.Q(\ram[255][3] ), 
	.D(FE_PHN669_n4665), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[255][2]  (.Q(\ram[255][2] ), 
	.D(FE_PHN973_n4664), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[255][1]  (.Q(\ram[255][1] ), 
	.D(FE_PHN781_n4663), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[255][0]  (.Q(\ram[255][0] ), 
	.D(FE_PHN3044_n4662), 
	.CK(clk));
   QDFFEHD \ram_reg[251][15]  (.Q(\ram[251][15] ), 
	.D(FE_PHN339_n4613), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][14]  (.Q(\ram[251][14] ), 
	.D(FE_PHN1293_n4612), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][13]  (.Q(\ram[251][13] ), 
	.D(FE_PHN1246_n4611), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][12]  (.Q(\ram[251][12] ), 
	.D(FE_PHN2175_n4610), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][11]  (.Q(\ram[251][11] ), 
	.D(FE_PHN499_n4609), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][10]  (.Q(\ram[251][10] ), 
	.D(FE_PHN1756_n4608), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][9]  (.Q(\ram[251][9] ), 
	.D(FE_PHN1141_n4607), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][8]  (.Q(\ram[251][8] ), 
	.D(FE_PHN2901_n4606), 
	.CK(clk_m__L3_N5));
   QDFFEHD \ram_reg[251][7]  (.Q(\ram[251][7] ), 
	.D(FE_PHN2638_n4605), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][6]  (.Q(\ram[251][6] ), 
	.D(FE_PHN567_n4604), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][5]  (.Q(\ram[251][5] ), 
	.D(FE_PHN513_n4603), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][4]  (.Q(\ram[251][4] ), 
	.D(FE_PHN444_n4602), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[251][3]  (.Q(\ram[251][3] ), 
	.D(FE_PHN1626_n4601), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[251][2]  (.Q(\ram[251][2] ), 
	.D(FE_PHN227_n4600), 
	.CK(clk_m__L3_N9));
   QDFFEHD \ram_reg[251][1]  (.Q(\ram[251][1] ), 
	.D(FE_PHN625_n4599), 
	.CK(clk_m__L3_N29));
   QDFFEHD \ram_reg[251][0]  (.Q(\ram[251][0] ), 
	.D(FE_PHN1060_n4598), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[247][15]  (.Q(\ram[247][15] ), 
	.D(FE_PHN2351_n4549), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][14]  (.Q(\ram[247][14] ), 
	.D(FE_PHN478_n4548), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[247][13]  (.Q(\ram[247][13] ), 
	.D(FE_PHN2792_n4547), 
	.CK(clk));
   QDFFEHD \ram_reg[247][12]  (.Q(\ram[247][12] ), 
	.D(FE_PHN1212_n4546), 
	.CK(clk));
   QDFFEHD \ram_reg[247][11]  (.Q(\ram[247][11] ), 
	.D(FE_PHN861_n4545), 
	.CK(clk));
   QDFFEHD \ram_reg[247][10]  (.Q(\ram[247][10] ), 
	.D(FE_PHN2324_n4544), 
	.CK(clk));
   QDFFEHD \ram_reg[247][9]  (.Q(\ram[247][9] ), 
	.D(FE_PHN1460_n4543), 
	.CK(clk));
   QDFFEHD \ram_reg[247][8]  (.Q(\ram[247][8] ), 
	.D(FE_PHN3004_n4542), 
	.CK(clk));
   QDFFEHD \ram_reg[247][7]  (.Q(\ram[247][7] ), 
	.D(FE_PHN3202_n4541), 
	.CK(clk_m__L3_N8));
   QDFFEHD \ram_reg[247][6]  (.Q(\ram[247][6] ), 
	.D(FE_PHN3162_n4540), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][5]  (.Q(\ram[247][5] ), 
	.D(FE_PHN2415_n4539), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][4]  (.Q(\ram[247][4] ), 
	.D(FE_PHN2934_n4538), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][3]  (.Q(\ram[247][3] ), 
	.D(FE_PHN1065_n4537), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[247][2]  (.Q(\ram[247][2] ), 
	.D(FE_PHN2238_n4536), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[247][1]  (.Q(\ram[247][1] ), 
	.D(FE_PHN1302_n4535), 
	.CK(clk_m__L3_N4));
   QDFFEHD \ram_reg[247][0]  (.Q(\ram[247][0] ), 
	.D(FE_PHN1248_n4534), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[243][15]  (.Q(\ram[243][15] ), 
	.D(FE_PHN1510_n4485), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][14]  (.Q(\ram[243][14] ), 
	.D(FE_PHN1746_n4484), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][13]  (.Q(\ram[243][13] ), 
	.D(FE_PHN1256_n4483), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][12]  (.Q(\ram[243][12] ), 
	.D(FE_PHN2331_n4482), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[243][11]  (.Q(\ram[243][11] ), 
	.D(FE_PHN1486_n4481), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[243][10]  (.Q(\ram[243][10] ), 
	.D(FE_PHN2710_n4480), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][9]  (.Q(\ram[243][9] ), 
	.D(FE_PHN313_n4479), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[243][8]  (.Q(\ram[243][8] ), 
	.D(FE_PHN1030_n4478), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[243][7]  (.Q(\ram[243][7] ), 
	.D(FE_PHN263_n4477), 
	.CK(clk_m__L3_N7));
   QDFFEHD \ram_reg[243][6]  (.Q(\ram[243][6] ), 
	.D(FE_PHN1721_n4476), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][5]  (.Q(\ram[243][5] ), 
	.D(FE_PHN386_n4475), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][4]  (.Q(\ram[243][4] ), 
	.D(FE_PHN348_n4474), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][3]  (.Q(\ram[243][3] ), 
	.D(FE_PHN819_n4473), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][2]  (.Q(\ram[243][2] ), 
	.D(FE_PHN1599_n4472), 
	.CK(clk_m__L3_N3));
   QDFFEHD \ram_reg[243][1]  (.Q(\ram[243][1] ), 
	.D(FE_PHN434_n4471), 
	.CK(clk_m__L3_N6));
   QDFFEHD \ram_reg[243][0]  (.Q(\ram[243][0] ), 
	.D(FE_PHN1156_n4470), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[239][15]  (.Q(\ram[239][15] ), 
	.D(FE_PHN5042_n4421), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][14]  (.Q(\ram[239][14] ), 
	.D(FE_PHN4729_n4420), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][13]  (.Q(\ram[239][13] ), 
	.D(FE_PHN4463_n4419), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][12]  (.Q(\ram[239][12] ), 
	.D(FE_PHN4552_n4418), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][11]  (.Q(\ram[239][11] ), 
	.D(FE_PHN4201_n4417), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][10]  (.Q(\ram[239][10] ), 
	.D(FE_PHN4616_n4416), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[239][9]  (.Q(\ram[239][9] ), 
	.D(FE_PHN3643_n4415), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[239][8]  (.Q(\ram[239][8] ), 
	.D(FE_PHN4713_n4414), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[239][7]  (.Q(\ram[239][7] ), 
	.D(FE_PHN4159_n4413), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][6]  (.Q(\ram[239][6] ), 
	.D(FE_PHN4665_n4412), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[239][5]  (.Q(\ram[239][5] ), 
	.D(FE_PHN4366_n4411), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][4]  (.Q(\ram[239][4] ), 
	.D(FE_PHN4178_n4410), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][3]  (.Q(\ram[239][3] ), 
	.D(FE_PHN6705_n4409), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[239][2]  (.Q(\ram[239][2] ), 
	.D(FE_PHN4279_n4408), 
	.CK(clk_m__L3_N55));
   QDFFEHD \ram_reg[239][1]  (.Q(\ram[239][1] ), 
	.D(FE_PHN4362_n4407), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[239][0]  (.Q(\ram[239][0] ), 
	.D(FE_PHN4076_n4406), 
	.CK(clk_m__L3_N56));
   QDFFEHD \ram_reg[235][15]  (.Q(\ram[235][15] ), 
	.D(FE_PHN1933_n4357), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][14]  (.Q(\ram[235][14] ), 
	.D(FE_PHN4095_n4356), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[235][13]  (.Q(\ram[235][13] ), 
	.D(FE_PHN4498_n4355), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[235][12]  (.Q(\ram[235][12] ), 
	.D(FE_PHN1250_n4354), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][11]  (.Q(\ram[235][11] ), 
	.D(FE_PHN3177_n4353), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][10]  (.Q(\ram[235][10] ), 
	.D(FE_PHN492_n4352), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][9]  (.Q(\ram[235][9] ), 
	.D(FE_PHN1873_n4351), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][8]  (.Q(\ram[235][8] ), 
	.D(FE_PHN4487_n4350), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[235][7]  (.Q(\ram[235][7] ), 
	.D(FE_PHN725_n4349), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][6]  (.Q(\ram[235][6] ), 
	.D(FE_PHN1268_n4348), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][5]  (.Q(\ram[235][5] ), 
	.D(FE_PHN1440_n4347), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[235][4]  (.Q(\ram[235][4] ), 
	.D(FE_PHN2001_n4346), 
	.CK(clk_m__L3_N18));
   QDFFEHD \ram_reg[235][3]  (.Q(\ram[235][3] ), 
	.D(FE_PHN2303_n4345), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][2]  (.Q(\ram[235][2] ), 
	.D(FE_PHN2532_n4344), 
	.CK(clk_m__L3_N17));
   QDFFEHD \ram_reg[235][1]  (.Q(\ram[235][1] ), 
	.D(FE_PHN4992_n4343), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[235][0]  (.Q(\ram[235][0] ), 
	.D(FE_PHN3322_n4342), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[231][15]  (.Q(\ram[231][15] ), 
	.D(FE_PHN858_n4293), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][14]  (.Q(\ram[231][14] ), 
	.D(FE_PHN4199_n4292), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][13]  (.Q(\ram[231][13] ), 
	.D(FE_PHN4300_n4291), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][12]  (.Q(\ram[231][12] ), 
	.D(FE_PHN4237_n4290), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][11]  (.Q(\ram[231][11] ), 
	.D(FE_PHN4220_n4289), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[231][10]  (.Q(\ram[231][10] ), 
	.D(FE_PHN200_n4288), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][9]  (.Q(\ram[231][9] ), 
	.D(FE_PHN761_n4287), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][8]  (.Q(\ram[231][8] ), 
	.D(FE_PHN4293_n4286), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[231][7]  (.Q(\ram[231][7] ), 
	.D(FE_PHN3460_n4285), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][6]  (.Q(\ram[231][6] ), 
	.D(FE_PHN4642_n4284), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[231][5]  (.Q(\ram[231][5] ), 
	.D(FE_PHN4390_n4283), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][4]  (.Q(\ram[231][4] ), 
	.D(FE_PHN454_n4282), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[231][3]  (.Q(\ram[231][3] ), 
	.D(FE_PHN4649_n4281), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[231][2]  (.Q(\ram[231][2] ), 
	.D(FE_PHN624_n4280), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[231][1]  (.Q(\ram[231][1] ), 
	.D(FE_PHN4132_n4279), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[231][0]  (.Q(\ram[231][0] ), 
	.D(FE_PHN4620_n4278), 
	.CK(clk_m__L3_N45));
   QDFFEHD \ram_reg[227][15]  (.Q(\ram[227][15] ), 
	.D(FE_PHN3855_n4229), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][14]  (.Q(\ram[227][14] ), 
	.D(FE_PHN4574_n4228), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][13]  (.Q(\ram[227][13] ), 
	.D(FE_PHN3844_n4227), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[227][12]  (.Q(\ram[227][12] ), 
	.D(FE_PHN4684_n4226), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][11]  (.Q(\ram[227][11] ), 
	.D(FE_PHN5395_n4225), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][10]  (.Q(\ram[227][10] ), 
	.D(FE_PHN2025_n4224), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[227][9]  (.Q(\ram[227][9] ), 
	.D(FE_PHN1707_n4223), 
	.CK(clk_m__L3_N1));
   QDFFEHD \ram_reg[227][8]  (.Q(\ram[227][8] ), 
	.D(FE_PHN4682_n4222), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][7]  (.Q(\ram[227][7] ), 
	.D(FE_PHN2159_n4221), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[227][6]  (.Q(\ram[227][6] ), 
	.D(FE_PHN4272_n4220), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][5]  (.Q(\ram[227][5] ), 
	.D(FE_PHN3630_n4219), 
	.CK(clk_m__L3_N40));
   QDFFEHD \ram_reg[227][4]  (.Q(\ram[227][4] ), 
	.D(FE_PHN4437_n4218), 
	.CK(clk_m__L3_N44));
   QDFFEHD \ram_reg[227][3]  (.Q(\ram[227][3] ), 
	.D(FE_PHN4364_n4217), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][2]  (.Q(\ram[227][2] ), 
	.D(FE_PHN2867_n4216), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[227][1]  (.Q(\ram[227][1] ), 
	.D(FE_PHN3915_n4215), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[227][0]  (.Q(\ram[227][0] ), 
	.D(FE_PHN3353_n4214), 
	.CK(clk_m__L3_N41));
   QDFFEHD \ram_reg[223][15]  (.Q(\ram[223][15] ), 
	.D(FE_PHN2093_n4165), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[223][14]  (.Q(\ram[223][14] ), 
	.D(FE_PHN4689_n4164), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][13]  (.Q(\ram[223][13] ), 
	.D(FE_PHN6668_n4163), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][12]  (.Q(\ram[223][12] ), 
	.D(FE_PHN3210_n4162), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][11]  (.Q(\ram[223][11] ), 
	.D(FE_PHN616_n4161), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[223][10]  (.Q(\ram[223][10] ), 
	.D(FE_PHN1516_n4160), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[223][9]  (.Q(\ram[223][9] ), 
	.D(FE_PHN2365_n4159), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][8]  (.Q(\ram[223][8] ), 
	.D(FE_PHN5682_n4158), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[223][7]  (.Q(\ram[223][7] ), 
	.D(FE_PHN1280_n4157), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[223][6]  (.Q(\ram[223][6] ), 
	.D(FE_PHN924_n4156), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][5]  (.Q(\ram[223][5] ), 
	.D(FE_PHN6686_n4155), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][4]  (.Q(\ram[223][4] ), 
	.D(FE_PHN1503_n4154), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[223][3]  (.Q(\ram[223][3] ), 
	.D(FE_PHN6661_n4153), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][2]  (.Q(\ram[223][2] ), 
	.D(FE_PHN1769_n4152), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[223][1]  (.Q(\ram[223][1] ), 
	.D(FE_PHN5758_n4151), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[223][0]  (.Q(\ram[223][0] ), 
	.D(FE_PHN5753_n4150), 
	.CK(clk_m__L3_N74));
   QDFFEHD \ram_reg[219][15]  (.Q(\ram[219][15] ), 
	.D(FE_PHN1946_n4101), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][14]  (.Q(\ram[219][14] ), 
	.D(FE_PHN2234_n4100), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][13]  (.Q(\ram[219][13] ), 
	.D(FE_PHN843_n4099), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][12]  (.Q(\ram[219][12] ), 
	.D(FE_PHN2842_n4098), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][11]  (.Q(\ram[219][11] ), 
	.D(FE_PHN4744_n4097), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][10]  (.Q(\ram[219][10] ), 
	.D(FE_PHN3157_n4096), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[219][9]  (.Q(\ram[219][9] ), 
	.D(FE_PHN618_n4095), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][8]  (.Q(\ram[219][8] ), 
	.D(FE_PHN4745_n4094), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][7]  (.Q(\ram[219][7] ), 
	.D(FE_PHN2936_n4093), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][6]  (.Q(\ram[219][6] ), 
	.D(FE_PHN233_n4092), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[219][5]  (.Q(\ram[219][5] ), 
	.D(FE_PHN714_n4091), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][4]  (.Q(\ram[219][4] ), 
	.D(FE_PHN2622_n4090), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][3]  (.Q(\ram[219][3] ), 
	.D(FE_PHN1383_n4089), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][2]  (.Q(\ram[219][2] ), 
	.D(FE_PHN1032_n4088), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[219][1]  (.Q(\ram[219][1] ), 
	.D(FE_PHN4727_n4087), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[219][0]  (.Q(\ram[219][0] ), 
	.D(FE_PHN1031_n4086), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[215][15]  (.Q(\ram[215][15] ), 
	.D(FE_PHN4530_n4037), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][14]  (.Q(\ram[215][14] ), 
	.D(FE_PHN4337_n4036), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][13]  (.Q(\ram[215][13] ), 
	.D(FE_PHN4412_n4035), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[215][12]  (.Q(\ram[215][12] ), 
	.D(FE_PHN4296_n4034), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[215][11]  (.Q(\ram[215][11] ), 
	.D(FE_PHN4181_n4033), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][10]  (.Q(\ram[215][10] ), 
	.D(FE_PHN6462_n4032), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][9]  (.Q(\ram[215][9] ), 
	.D(FE_PHN4149_n4031), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[215][8]  (.Q(\ram[215][8] ), 
	.D(FE_PHN4515_n4030), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[215][7]  (.Q(\ram[215][7] ), 
	.D(FE_PHN4668_n4029), 
	.CK(clk_m__L3_N54));
   QDFFEHD \ram_reg[215][6]  (.Q(\ram[215][6] ), 
	.D(FE_PHN4160_n4028), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[215][5]  (.Q(\ram[215][5] ), 
	.D(FE_PHN6450_n4027), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[215][4]  (.Q(\ram[215][4] ), 
	.D(FE_PHN4548_n4026), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][3]  (.Q(\ram[215][3] ), 
	.D(FE_PHN4344_n4025), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][2]  (.Q(\ram[215][2] ), 
	.D(FE_PHN250_n4024), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][1]  (.Q(\ram[215][1] ), 
	.D(FE_PHN4262_n4023), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[215][0]  (.Q(\ram[215][0] ), 
	.D(FE_PHN4157_n4022), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[211][15]  (.Q(\ram[211][15] ), 
	.D(FE_PHN621_n3973), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[211][14]  (.Q(\ram[211][14] ), 
	.D(FE_PHN5430_n3972), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[211][13]  (.Q(\ram[211][13] ), 
	.D(FE_PHN4501_n3971), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][12]  (.Q(\ram[211][12] ), 
	.D(FE_PHN3565_n3970), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][11]  (.Q(\ram[211][11] ), 
	.D(FE_PHN4425_n3969), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[211][10]  (.Q(\ram[211][10] ), 
	.D(FE_PHN6654_n3968), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][9]  (.Q(\ram[211][9] ), 
	.D(FE_PHN332_n3967), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][8]  (.Q(\ram[211][8] ), 
	.D(FE_PHN4253_n3966), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][7]  (.Q(\ram[211][7] ), 
	.D(FE_PHN3775_n3965), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][6]  (.Q(\ram[211][6] ), 
	.D(FE_PHN3704_n3964), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][5]  (.Q(\ram[211][5] ), 
	.D(FE_PHN4461_n3963), 
	.CK(clk_m__L3_N39));
   QDFFEHD \ram_reg[211][4]  (.Q(\ram[211][4] ), 
	.D(FE_PHN4594_n3962), 
	.CK(clk_m__L3_N42));
   QDFFEHD \ram_reg[211][3]  (.Q(\ram[211][3] ), 
	.D(FE_PHN4365_n3961), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[211][2]  (.Q(\ram[211][2] ), 
	.D(FE_PHN6675_n3960), 
	.CK(clk_m__L3_N43));
   QDFFEHD \ram_reg[211][1]  (.Q(\ram[211][1] ), 
	.D(FE_PHN3352_n3959), 
	.CK(clk_m__L3_N57));
   QDFFEHD \ram_reg[211][0]  (.Q(\ram[211][0] ), 
	.D(FE_PHN4613_n3958), 
	.CK(clk_m__L3_N58));
   QDFFEHD \ram_reg[207][15]  (.Q(\ram[207][15] ), 
	.D(FE_PHN610_n3909), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][14]  (.Q(\ram[207][14] ), 
	.D(FE_PHN3057_n3908), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][13]  (.Q(\ram[207][13] ), 
	.D(FE_PHN898_n3907), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[207][12]  (.Q(\ram[207][12] ), 
	.D(FE_PHN1876_n3906), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][11]  (.Q(\ram[207][11] ), 
	.D(FE_PHN196_n3905), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][10]  (.Q(\ram[207][10] ), 
	.D(FE_PHN1890_n3904), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][9]  (.Q(\ram[207][9] ), 
	.D(FE_PHN2483_n3903), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[207][8]  (.Q(\ram[207][8] ), 
	.D(FE_PHN1970_n3902), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[207][7]  (.Q(\ram[207][7] ), 
	.D(FE_PHN2133_n3901), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][6]  (.Q(\ram[207][6] ), 
	.D(FE_PHN1800_n3900), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[207][5]  (.Q(\ram[207][5] ), 
	.D(FE_PHN1166_n3899), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][4]  (.Q(\ram[207][4] ), 
	.D(FE_PHN2548_n3898), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][3]  (.Q(\ram[207][3] ), 
	.D(FE_PHN2290_n3897), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][2]  (.Q(\ram[207][2] ), 
	.D(FE_PHN2816_n3896), 
	.CK(clk_m__L3_N37));
   QDFFEHD \ram_reg[207][1]  (.Q(\ram[207][1] ), 
	.D(FE_PHN2479_n3895), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[207][0]  (.Q(\ram[207][0] ), 
	.D(FE_PHN2421_n3894), 
	.CK(clk_m__L3_N48));
   QDFFEHD \ram_reg[203][15]  (.Q(\ram[203][15] ), 
	.D(FE_PHN1203_n3845), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[203][14]  (.Q(\ram[203][14] ), 
	.D(FE_PHN2484_n3844), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][13]  (.Q(\ram[203][13] ), 
	.D(FE_PHN3174_n3843), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[203][12]  (.Q(\ram[203][12] ), 
	.D(FE_PHN461_n3842), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[203][11]  (.Q(\ram[203][11] ), 
	.D(FE_PHN1201_n3841), 
	.CK(clk_m__L3_N34));
   QDFFEHD \ram_reg[203][10]  (.Q(\ram[203][10] ), 
	.D(FE_PHN2276_n3840), 
	.CK(clk_m__L3_N32));
   QDFFEHD \ram_reg[203][9]  (.Q(\ram[203][9] ), 
	.D(FE_PHN955_n3839), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][8]  (.Q(\ram[203][8] ), 
	.D(FE_PHN511_n3838), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][7]  (.Q(\ram[203][7] ), 
	.D(FE_PHN1345_n3837), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][6]  (.Q(\ram[203][6] ), 
	.D(FE_PHN1562_n3836), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][5]  (.Q(\ram[203][5] ), 
	.D(FE_PHN1131_n3835), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][4]  (.Q(\ram[203][4] ), 
	.D(FE_PHN1341_n3834), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][3]  (.Q(\ram[203][3] ), 
	.D(FE_PHN1912_n3833), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][2]  (.Q(\ram[203][2] ), 
	.D(FE_PHN879_n3832), 
	.CK(clk_m__L3_N35));
   QDFFEHD \ram_reg[203][1]  (.Q(\ram[203][1] ), 
	.D(FE_PHN1215_n3831), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[203][0]  (.Q(\ram[203][0] ), 
	.D(FE_PHN2840_n3830), 
	.CK(clk_m__L3_N47));
   QDFFEHD \ram_reg[199][15]  (.Q(\ram[199][15] ), 
	.D(FE_PHN578_n3781), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][14]  (.Q(\ram[199][14] ), 
	.D(FE_PHN1358_n3780), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][13]  (.Q(\ram[199][13] ), 
	.D(FE_PHN2268_n3779), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[199][12]  (.Q(\ram[199][12] ), 
	.D(FE_PHN3040_n3778), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[199][11]  (.Q(\ram[199][11] ), 
	.D(FE_PHN3123_n3777), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][10]  (.Q(\ram[199][10] ), 
	.D(FE_PHN2322_n3776), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[199][9]  (.Q(\ram[199][9] ), 
	.D(FE_PHN1992_n3775), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[199][8]  (.Q(\ram[199][8] ), 
	.D(FE_PHN1443_n3774), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][7]  (.Q(\ram[199][7] ), 
	.D(FE_PHN1518_n3773), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][6]  (.Q(\ram[199][6] ), 
	.D(FE_PHN265_n3772), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][5]  (.Q(\ram[199][5] ), 
	.D(n3771), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][4]  (.Q(\ram[199][4] ), 
	.D(FE_PHN2150_n3770), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][3]  (.Q(\ram[199][3] ), 
	.D(FE_PHN3171_n3769), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[199][2]  (.Q(\ram[199][2] ), 
	.D(FE_PHN315_n3768), 
	.CK(clk_m__L3_N36));
   QDFFEHD \ram_reg[199][1]  (.Q(\ram[199][1] ), 
	.D(FE_PHN913_n3767), 
	.CK(clk_m__L3_N66));
   QDFFEHD \ram_reg[199][0]  (.Q(\ram[199][0] ), 
	.D(FE_PHN1145_n3766), 
	.CK(clk_m__L3_N60));
   QDFFEHD \ram_reg[195][15]  (.Q(\ram[195][15] ), 
	.D(FE_PHN1297_n3717), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][14]  (.Q(\ram[195][14] ), 
	.D(FE_PHN2192_n3716), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][13]  (.Q(\ram[195][13] ), 
	.D(FE_PHN1976_n3715), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[195][12]  (.Q(\ram[195][12] ), 
	.D(FE_PHN2970_n3714), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[195][11]  (.Q(\ram[195][11] ), 
	.D(FE_PHN1428_n3713), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][10]  (.Q(\ram[195][10] ), 
	.D(FE_PHN1582_n3712), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][9]  (.Q(\ram[195][9] ), 
	.D(FE_PHN1690_n3711), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][8]  (.Q(\ram[195][8] ), 
	.D(FE_PHN779_n3710), 
	.CK(clk_m__L3_N30));
   QDFFEHD \ram_reg[195][7]  (.Q(\ram[195][7] ), 
	.D(FE_PHN1692_n3709), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][6]  (.Q(\ram[195][6] ), 
	.D(FE_PHN772_n3708), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][5]  (.Q(\ram[195][5] ), 
	.D(FE_PHN2343_n3707), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][4]  (.Q(\ram[195][4] ), 
	.D(FE_PHN1048_n3706), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][3]  (.Q(\ram[195][3] ), 
	.D(FE_PHN1427_n3705), 
	.CK(clk_m__L3_N46));
   QDFFEHD \ram_reg[195][2]  (.Q(\ram[195][2] ), 
	.D(FE_PHN2561_n3704), 
	.CK(clk_m__L3_N38));
   QDFFEHD \ram_reg[195][1]  (.Q(\ram[195][1] ), 
	.D(FE_PHN1371_n3703), 
	.CK(clk_m__L3_N33));
   QDFFEHD \ram_reg[195][0]  (.Q(\ram[195][0] ), 
	.D(FE_PHN666_n3702), 
	.CK(clk_m__L3_N31));
   QDFFEHD \ram_reg[191][15]  (.Q(\ram[191][15] ), 
	.D(FE_PHN2045_n3653), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[191][14]  (.Q(\ram[191][14] ), 
	.D(FE_PHN1531_n3652), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[191][13]  (.Q(\ram[191][13] ), 
	.D(FE_PHN707_n3651), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[191][12]  (.Q(\ram[191][12] ), 
	.D(FE_PHN1320_n3650), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[191][11]  (.Q(\ram[191][11] ), 
	.D(FE_PHN2410_n3649), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[191][10]  (.Q(\ram[191][10] ), 
	.D(FE_PHN936_n3648), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][9]  (.Q(\ram[191][9] ), 
	.D(FE_PHN2579_n3647), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[191][8]  (.Q(\ram[191][8] ), 
	.D(FE_PHN1000_n3646), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][7]  (.Q(\ram[191][7] ), 
	.D(FE_PHN754_n3645), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][6]  (.Q(\ram[191][6] ), 
	.D(FE_PHN1392_n3644), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[191][5]  (.Q(\ram[191][5] ), 
	.D(FE_PHN827_n3643), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[191][4]  (.Q(\ram[191][4] ), 
	.D(FE_PHN1843_n3642), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][3]  (.Q(\ram[191][3] ), 
	.D(FE_PHN2919_n3641), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[191][2]  (.Q(\ram[191][2] ), 
	.D(FE_PHN3146_n3640), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[191][1]  (.Q(\ram[191][1] ), 
	.D(FE_PHN3001_n3639), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[191][0]  (.Q(\ram[191][0] ), 
	.D(FE_PHN2488_n3638), 
	.CK(clk_m__L3_N105));
   QDFFEHD \ram_reg[187][15]  (.Q(\ram[187][15] ), 
	.D(FE_PHN963_n3589), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][14]  (.Q(\ram[187][14] ), 
	.D(FE_PHN1093_n3588), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][13]  (.Q(\ram[187][13] ), 
	.D(FE_PHN767_n3587), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[187][12]  (.Q(\ram[187][12] ), 
	.D(FE_PHN1764_n3586), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[187][11]  (.Q(\ram[187][11] ), 
	.D(FE_PHN1823_n3585), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[187][10]  (.Q(\ram[187][10] ), 
	.D(FE_PHN111_n3584), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[187][9]  (.Q(\ram[187][9] ), 
	.D(FE_PHN1199_n3583), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[187][8]  (.Q(\ram[187][8] ), 
	.D(FE_PHN1438_n3582), 
	.CK(clk_m__L3_N102));
   QDFFEHD \ram_reg[187][7]  (.Q(\ram[187][7] ), 
	.D(FE_PHN1217_n3581), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[187][6]  (.Q(\ram[187][6] ), 
	.D(FE_PHN167_n3580), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[187][5]  (.Q(\ram[187][5] ), 
	.D(FE_PHN446_n3579), 
	.CK(clk_m__L3_N106));
   QDFFEHD \ram_reg[187][4]  (.Q(\ram[187][4] ), 
	.D(FE_PHN1465_n3578), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[187][3]  (.Q(\ram[187][3] ), 
	.D(FE_PHN2424_n3577), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[187][2]  (.Q(\ram[187][2] ), 
	.D(FE_PHN917_n3576), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][1]  (.Q(\ram[187][1] ), 
	.D(FE_PHN704_n3575), 
	.CK(clk_m__L3_N101));
   QDFFEHD \ram_reg[187][0]  (.Q(\ram[187][0] ), 
	.D(FE_PHN331_n3574), 
	.CK(clk_m__N0));
   QDFFEHD \ram_reg[183][15]  (.Q(\ram[183][15] ), 
	.D(FE_PHN2657_n3525), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[183][14]  (.Q(\ram[183][14] ), 
	.D(FE_PHN2530_n3524), 
	.CK(clk_m__L3_N100));
   QDFFEHD \ram_reg[183][13]  (.Q(\ram[183][13] ), 
	.D(FE_PHN2477_n3523), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[183][12]  (.Q(\ram[183][12] ), 
	.D(FE_PHN2523_n3522), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][11]  (.Q(\ram[183][11] ), 
	.D(FE_PHN1260_n3521), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[183][10]  (.Q(\ram[183][10] ), 
	.D(FE_PHN3212_n3520), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][9]  (.Q(\ram[183][9] ), 
	.D(FE_PHN3173_n3519), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][8]  (.Q(\ram[183][8] ), 
	.D(FE_PHN2819_n3518), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][7]  (.Q(\ram[183][7] ), 
	.D(FE_PHN2147_n3517), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[183][6]  (.Q(\ram[183][6] ), 
	.D(FE_PHN1957_n3516), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[183][5]  (.Q(\ram[183][5] ), 
	.D(FE_PHN1436_n3515), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[183][4]  (.Q(\ram[183][4] ), 
	.D(FE_PHN1570_n3514), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][3]  (.Q(\ram[183][3] ), 
	.D(FE_PHN636_n3513), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[183][2]  (.Q(\ram[183][2] ), 
	.D(FE_PHN488_n3512), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][1]  (.Q(\ram[183][1] ), 
	.D(FE_PHN711_n3511), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[183][0]  (.Q(\ram[183][0] ), 
	.D(FE_PHN579_n3510), 
	.CK(clk_m__L3_N104));
   QDFFEHD \ram_reg[179][15]  (.Q(\ram[179][15] ), 
	.D(FE_PHN3219_n3461), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][14]  (.Q(\ram[179][14] ), 
	.D(FE_PHN1832_n3460), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][13]  (.Q(\ram[179][13] ), 
	.D(FE_PHN3082_n3459), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[179][12]  (.Q(\ram[179][12] ), 
	.D(FE_PHN2855_n3458), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][11]  (.Q(\ram[179][11] ), 
	.D(FE_PHN2556_n3457), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][10]  (.Q(\ram[179][10] ), 
	.D(FE_PHN2329_n3456), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][9]  (.Q(\ram[179][9] ), 
	.D(FE_PHN2809_n3455), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][8]  (.Q(\ram[179][8] ), 
	.D(FE_PHN2581_n3454), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[179][7]  (.Q(\ram[179][7] ), 
	.D(FE_PHN3094_n3453), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][6]  (.Q(\ram[179][6] ), 
	.D(FE_PHN1771_n3452), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[179][5]  (.Q(\ram[179][5] ), 
	.D(FE_PHN3229_n3451), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[179][4]  (.Q(\ram[179][4] ), 
	.D(FE_PHN1722_n3450), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][3]  (.Q(\ram[179][3] ), 
	.D(FE_PHN1033_n3449), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[179][2]  (.Q(\ram[179][2] ), 
	.D(FE_PHN2778_n3448), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[179][1]  (.Q(\ram[179][1] ), 
	.D(FE_PHN2937_n3447), 
	.CK(clk_m__L3_N117));
   QDFFEHD \ram_reg[179][0]  (.Q(\ram[179][0] ), 
	.D(FE_PHN1765_n3446), 
	.CK(clk_m__L3_N115));
   QDFFEHD \ram_reg[175][15]  (.Q(\ram[175][15] ), 
	.D(FE_PHN1386_n3397), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][14]  (.Q(\ram[175][14] ), 
	.D(FE_PHN1037_n3396), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][13]  (.Q(\ram[175][13] ), 
	.D(FE_PHN1380_n3395), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[175][12]  (.Q(\ram[175][12] ), 
	.D(FE_PHN2651_n3394), 
	.CK(clk));
   QDFFEHD \ram_reg[175][11]  (.Q(\ram[175][11] ), 
	.D(FE_PHN1441_n3393), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][10]  (.Q(\ram[175][10] ), 
	.D(FE_PHN2947_n3392), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][9]  (.Q(\ram[175][9] ), 
	.D(FE_PHN1362_n3391), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][8]  (.Q(\ram[175][8] ), 
	.D(FE_PHN2086_n3390), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][7]  (.Q(\ram[175][7] ), 
	.D(FE_PHN482_n3389), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][6]  (.Q(\ram[175][6] ), 
	.D(FE_PHN3172_n3388), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][5]  (.Q(\ram[175][5] ), 
	.D(FE_PHN2959_n3387), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][4]  (.Q(\ram[175][4] ), 
	.D(FE_PHN584_n3386), 
	.CK(clk_m__L3_N2));
   QDFFEHD \ram_reg[175][3]  (.Q(\ram[175][3] ), 
	.D(FE_PHN2155_n3385), 
	.CK(clk_m__L3_N19));
   QDFFEHD \ram_reg[175][2]  (.Q(\ram[175][2] ), 
	.D(FE_PHN994_n3384), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][1]  (.Q(\ram[175][1] ), 
	.D(FE_PHN1437_n3383), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[175][0]  (.Q(\ram[175][0] ), 
	.D(FE_PHN1991_n3382), 
	.CK(clk_m__L3_N16));
   QDFFEHD \ram_reg[171][15]  (.Q(\ram[171][15] ), 
	.D(FE_PHN1309_n3333), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][14]  (.Q(\ram[171][14] ), 
	.D(FE_PHN3089_n3332), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][13]  (.Q(\ram[171][13] ), 
	.D(FE_PHN2783_n3331), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][12]  (.Q(\ram[171][12] ), 
	.D(FE_PHN1543_n3330), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][11]  (.Q(\ram[171][11] ), 
	.D(FE_PHN532_n3329), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][10]  (.Q(\ram[171][10] ), 
	.D(FE_PHN3090_n3328), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][9]  (.Q(\ram[171][9] ), 
	.D(FE_PHN502_n3327), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][8]  (.Q(\ram[171][8] ), 
	.D(FE_PHN1002_n3326), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][7]  (.Q(\ram[171][7] ), 
	.D(FE_PHN1154_n3325), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][6]  (.Q(\ram[171][6] ), 
	.D(FE_PHN763_n3324), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][5]  (.Q(\ram[171][5] ), 
	.D(FE_PHN508_n3323), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][4]  (.Q(\ram[171][4] ), 
	.D(FE_PHN1354_n3322), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[171][3]  (.Q(\ram[171][3] ), 
	.D(FE_PHN2961_n3321), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][2]  (.Q(\ram[171][2] ), 
	.D(FE_PHN2810_n3320), 
	.CK(clk_m__L3_N15));
   QDFFEHD \ram_reg[171][1]  (.Q(\ram[171][1] ), 
	.D(FE_PHN3072_n3319), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[171][0]  (.Q(\ram[171][0] ), 
	.D(FE_PHN1331_n3318), 
	.CK(clk_m__L3_N11));
   QDFFEHD \ram_reg[167][15]  (.Q(\ram[167][15] ), 
	.D(FE_PHN2019_n3269), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[167][14]  (.Q(\ram[167][14] ), 
	.D(FE_PHN1466_n3268), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][13]  (.Q(\ram[167][13] ), 
	.D(FE_PHN705_n3267), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][12]  (.Q(\ram[167][12] ), 
	.D(FE_PHN1381_n3266), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][11]  (.Q(\ram[167][11] ), 
	.D(FE_PHN4968_n3265), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][10]  (.Q(\ram[167][10] ), 
	.D(FE_PHN1195_n3264), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][9]  (.Q(\ram[167][9] ), 
	.D(FE_PHN4369_n3263), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][8]  (.Q(\ram[167][8] ), 
	.D(FE_PHN4446_n3262), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][7]  (.Q(\ram[167][7] ), 
	.D(FE_PHN3025_n3261), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[167][6]  (.Q(\ram[167][6] ), 
	.D(FE_PHN4069_n3260), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][5]  (.Q(\ram[167][5] ), 
	.D(FE_PHN2514_n3259), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][4]  (.Q(\ram[167][4] ), 
	.D(FE_PHN4686_n3258), 
	.CK(clk_m__L3_N12));
   QDFFEHD \ram_reg[167][3]  (.Q(\ram[167][3] ), 
	.D(FE_PHN4580_n3257), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][2]  (.Q(\ram[167][2] ), 
	.D(FE_PHN1741_n3256), 
	.CK(clk_m__L3_N14));
   QDFFEHD \ram_reg[167][1]  (.Q(\ram[167][1] ), 
	.D(FE_PHN4652_n3255), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[167][0]  (.Q(\ram[167][0] ), 
	.D(FE_PHN945_n3254), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[163][15]  (.Q(\ram[163][15] ), 
	.D(FE_PHN2770_n3205), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][14]  (.Q(\ram[163][14] ), 
	.D(FE_PHN2056_n3204), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][13]  (.Q(\ram[163][13] ), 
	.D(FE_PHN2302_n3203), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][12]  (.Q(\ram[163][12] ), 
	.D(FE_PHN939_n3202), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][11]  (.Q(\ram[163][11] ), 
	.D(FE_PHN829_n3201), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][10]  (.Q(\ram[163][10] ), 
	.D(FE_PHN1204_n3200), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][9]  (.Q(\ram[163][9] ), 
	.D(FE_PHN1667_n3199), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][8]  (.Q(\ram[163][8] ), 
	.D(FE_PHN1411_n3198), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][7]  (.Q(\ram[163][7] ), 
	.D(FE_PHN1171_n3197), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[163][6]  (.Q(\ram[163][6] ), 
	.D(FE_PHN1359_n3196), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[163][5]  (.Q(\ram[163][5] ), 
	.D(FE_PHN948_n3195), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][4]  (.Q(\ram[163][4] ), 
	.D(FE_PHN732_n3194), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][3]  (.Q(\ram[163][3] ), 
	.D(FE_PHN1871_n3193), 
	.CK(clk_m__L3_N10));
   QDFFEHD \ram_reg[163][2]  (.Q(\ram[163][2] ), 
	.D(FE_PHN1118_n3192), 
	.CK(clk_m__L3_N13));
   QDFFEHD \ram_reg[163][1]  (.Q(\ram[163][1] ), 
	.D(FE_PHN3107_n3191), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[163][0]  (.Q(\ram[163][0] ), 
	.D(FE_PHN2398_n3190), 
	.CK(clk_m__L3_N27));
   QDFFEHD \ram_reg[159][15]  (.Q(\ram[159][15] ), 
	.D(FE_PHN4465_n3141), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[159][14]  (.Q(\ram[159][14] ), 
	.D(FE_PHN4525_n3140), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][13]  (.Q(\ram[159][13] ), 
	.D(FE_PHN4591_n3139), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][12]  (.Q(\ram[159][12] ), 
	.D(FE_PHN4210_n3138), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][11]  (.Q(\ram[159][11] ), 
	.D(FE_PHN3553_n3137), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[159][10]  (.Q(\ram[159][10] ), 
	.D(FE_PHN4627_n3136), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[159][9]  (.Q(\ram[159][9] ), 
	.D(FE_PHN4731_n3135), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[159][8]  (.Q(\ram[159][8] ), 
	.D(FE_PHN4110_n3134), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[159][7]  (.Q(\ram[159][7] ), 
	.D(FE_PHN4184_n3133), 
	.CK(clk_m__L3_N26));
   QDFFEHD \ram_reg[159][6]  (.Q(\ram[159][6] ), 
	.D(FE_PHN4270_n3132), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[159][5]  (.Q(\ram[159][5] ), 
	.D(FE_PHN4658_n3131), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[159][4]  (.Q(\ram[159][4] ), 
	.D(FE_PHN4632_n3130), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[159][3]  (.Q(\ram[159][3] ), 
	.D(FE_PHN3881_n3129), 
	.CK(clk_m__L3_N28));
   QDFFEHD \ram_reg[159][2]  (.Q(\ram[159][2] ), 
	.D(FE_PHN4065_n3128), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[159][1]  (.Q(\ram[159][1] ), 
	.D(FE_PHN5545_n3127), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[159][0]  (.Q(\ram[159][0] ), 
	.D(FE_PHN4692_n3126), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[155][15]  (.Q(\ram[155][15] ), 
	.D(FE_PHN4196_n3077), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[155][14]  (.Q(\ram[155][14] ), 
	.D(FE_PHN4478_n3076), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][13]  (.Q(\ram[155][13] ), 
	.D(FE_PHN4421_n3075), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][12]  (.Q(\ram[155][12] ), 
	.D(FE_PHN4385_n3074), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][11]  (.Q(\ram[155][11] ), 
	.D(FE_PHN4227_n3073), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][10]  (.Q(\ram[155][10] ), 
	.D(FE_PHN3679_n3072), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[155][9]  (.Q(\ram[155][9] ), 
	.D(FE_PHN4276_n3071), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[155][8]  (.Q(\ram[155][8] ), 
	.D(FE_PHN4202_n3070), 
	.CK(clk_m__L3_N93));
   QDFFEHD \ram_reg[155][7]  (.Q(\ram[155][7] ), 
	.D(FE_PHN4512_n3069), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][6]  (.Q(\ram[155][6] ), 
	.D(FE_PHN5777_n3068), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][5]  (.Q(\ram[155][5] ), 
	.D(FE_PHN3906_n3067), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[155][4]  (.Q(\ram[155][4] ), 
	.D(FE_PHN4551_n3066), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[155][3]  (.Q(\ram[155][3] ), 
	.D(FE_PHN4509_n3065), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][2]  (.Q(\ram[155][2] ), 
	.D(FE_PHN3334_n3064), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][1]  (.Q(\ram[155][1] ), 
	.D(FE_PHN4388_n3063), 
	.CK(clk_m__L3_N22));
   QDFFEHD \ram_reg[155][0]  (.Q(\ram[155][0] ), 
	.D(FE_PHN4723_n3062), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[151][15]  (.Q(\ram[151][15] ), 
	.D(FE_PHN4482_n3013), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][14]  (.Q(\ram[151][14] ), 
	.D(FE_PHN4195_n3012), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][13]  (.Q(\ram[151][13] ), 
	.D(FE_PHN4420_n3011), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][12]  (.Q(\ram[151][12] ), 
	.D(FE_PHN4106_n3010), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[151][11]  (.Q(\ram[151][11] ), 
	.D(FE_PHN4126_n3009), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[151][10]  (.Q(\ram[151][10] ), 
	.D(FE_PHN4725_n3008), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[151][9]  (.Q(\ram[151][9] ), 
	.D(FE_PHN4214_n3007), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[151][8]  (.Q(\ram[151][8] ), 
	.D(FE_PHN4404_n3006), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[151][7]  (.Q(\ram[151][7] ), 
	.D(FE_PHN3749_n3005), 
	.CK(clk_m__L3_N127));
   QDFFEHD \ram_reg[151][6]  (.Q(\ram[151][6] ), 
	.D(FE_PHN5680_n3004), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[151][5]  (.Q(\ram[151][5] ), 
	.D(FE_PHN4158_n3003), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[151][4]  (.Q(\ram[151][4] ), 
	.D(FE_PHN3520_n3002), 
	.CK(clk_m__L3_N52));
   QDFFEHD \ram_reg[151][3]  (.Q(\ram[151][3] ), 
	.D(FE_PHN5502_n3001), 
	.CK(clk_m__L3_N53));
   QDFFEHD \ram_reg[151][2]  (.Q(\ram[151][2] ), 
	.D(FE_PHN4174_n3000), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[151][1]  (.Q(\ram[151][1] ), 
	.D(FE_PHN4175_n2999), 
	.CK(clk_m__L3_N49));
   QDFFEHD \ram_reg[151][0]  (.Q(\ram[151][0] ), 
	.D(FE_PHN4466_n2998), 
	.CK(clk_m__L3_N126));
   QDFFEHD \ram_reg[147][15]  (.Q(\ram[147][15] ), 
	.D(FE_PHN3147_n2949), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[147][14]  (.Q(\ram[147][14] ), 
	.D(FE_PHN498_n2948), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[147][13]  (.Q(\ram[147][13] ), 
	.D(FE_PHN806_n2947), 
	.CK(clk_m__L3_N89));
   QDFFEHD \ram_reg[147][12]  (.Q(\ram[147][12] ), 
	.D(FE_PHN4483_n2946), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][11]  (.Q(\ram[147][11] ), 
	.D(FE_PHN4376_n2945), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][10]  (.Q(\ram[147][10] ), 
	.D(FE_PHN3996_n2944), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[147][9]  (.Q(\ram[147][9] ), 
	.D(FE_PHN4702_n2943), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][8]  (.Q(\ram[147][8] ), 
	.D(FE_PHN540_n2942), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[147][7]  (.Q(\ram[147][7] ), 
	.D(FE_PHN5738_n2941), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][6]  (.Q(\ram[147][6] ), 
	.D(FE_PHN1324_n2940), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][5]  (.Q(\ram[147][5] ), 
	.D(FE_PHN833_n2939), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][4]  (.Q(\ram[147][4] ), 
	.D(FE_PHN4810_n2938), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][3]  (.Q(\ram[147][3] ), 
	.D(FE_PHN524_n2937), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][2]  (.Q(\ram[147][2] ), 
	.D(FE_PHN4651_n2936), 
	.CK(clk_m__L3_N95));
   QDFFEHD \ram_reg[147][1]  (.Q(\ram[147][1] ), 
	.D(FE_PHN6487_n2935), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[147][0]  (.Q(\ram[147][0] ), 
	.D(FE_PHN5459_n2934), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[143][15]  (.Q(\ram[143][15] ), 
	.D(FE_PHN3024_n2885), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[143][14]  (.Q(\ram[143][14] ), 
	.D(FE_PHN2015_n2884), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[143][13]  (.Q(\ram[143][13] ), 
	.D(FE_PHN2358_n2883), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[143][12]  (.Q(\ram[143][12] ), 
	.D(FE_PHN2603_n2882), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[143][11]  (.Q(\ram[143][11] ), 
	.D(FE_PHN1526_n2881), 
	.CK(clk_m__L3_N108));
   QDFFEHD \ram_reg[143][10]  (.Q(\ram[143][10] ), 
	.D(n2880), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[143][9]  (.Q(\ram[143][9] ), 
	.D(FE_PHN1754_n2879), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[143][8]  (.Q(\ram[143][8] ), 
	.D(FE_PHN1842_n2878), 
	.CK(clk_m__L3_N107));
   QDFFEHD \ram_reg[143][7]  (.Q(\ram[143][7] ), 
	.D(FE_PHN1492_n2877), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[143][6]  (.Q(\ram[143][6] ), 
	.D(FE_PHN5681_n2876), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[143][5]  (.Q(\ram[143][5] ), 
	.D(FE_PHN2741_n2875), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[143][4]  (.Q(\ram[143][4] ), 
	.D(FE_PHN1995_n2874), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[143][3]  (.Q(\ram[143][3] ), 
	.D(FE_PHN6593_n2873), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[143][2]  (.Q(\ram[143][2] ), 
	.D(FE_PHN2697_n2872), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[143][1]  (.Q(\ram[143][1] ), 
	.D(FE_PHN2625_n2871), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[143][0]  (.Q(\ram[143][0] ), 
	.D(FE_PHN3181_n2870), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[139][15]  (.Q(\ram[139][15] ), 
	.D(FE_PHN2091_n2821), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][14]  (.Q(\ram[139][14] ), 
	.D(FE_PHN2448_n2820), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][13]  (.Q(\ram[139][13] ), 
	.D(FE_PHN1335_n2819), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][12]  (.Q(\ram[139][12] ), 
	.D(FE_PHN467_n2818), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][11]  (.Q(\ram[139][11] ), 
	.D(FE_PHN2823_n2817), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][10]  (.Q(\ram[139][10] ), 
	.D(FE_PHN1139_n2816), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][9]  (.Q(\ram[139][9] ), 
	.D(FE_PHN3081_n2815), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[139][8]  (.Q(\ram[139][8] ), 
	.D(FE_PHN2140_n2814), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][7]  (.Q(\ram[139][7] ), 
	.D(FE_PHN2247_n2813), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][6]  (.Q(\ram[139][6] ), 
	.D(FE_PHN1372_n2812), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[139][5]  (.Q(\ram[139][5] ), 
	.D(FE_PHN688_n2811), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[139][4]  (.Q(\ram[139][4] ), 
	.D(FE_PHN1902_n2810), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[139][3]  (.Q(\ram[139][3] ), 
	.D(FE_PHN872_n2809), 
	.CK(clk_m__L3_N25));
   QDFFEHD \ram_reg[139][2]  (.Q(\ram[139][2] ), 
	.D(FE_PHN901_n2808), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[139][1]  (.Q(\ram[139][1] ), 
	.D(FE_PHN1100_n2807), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[139][0]  (.Q(\ram[139][0] ), 
	.D(FE_PHN2173_n2806), 
	.CK(clk_m__L3_N92));
   QDFFEHD \ram_reg[135][15]  (.Q(\ram[135][15] ), 
	.D(FE_PHN2721_n2757), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[135][14]  (.Q(\ram[135][14] ), 
	.D(FE_PHN2844_n2756), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[135][13]  (.Q(\ram[135][13] ), 
	.D(FE_PHN2252_n2755), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[135][12]  (.Q(\ram[135][12] ), 
	.D(FE_PHN3622_n2754), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][11]  (.Q(\ram[135][11] ), 
	.D(FE_PHN3856_n2753), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[135][10]  (.Q(\ram[135][10] ), 
	.D(FE_PHN1947_n2752), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][9]  (.Q(\ram[135][9] ), 
	.D(FE_PHN880_n2751), 
	.CK(clk_m__L3_N94));
   QDFFEHD \ram_reg[135][8]  (.Q(\ram[135][8] ), 
	.D(FE_PHN5663_n2750), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][7]  (.Q(\ram[135][7] ), 
	.D(FE_PHN5686_n2749), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][6]  (.Q(\ram[135][6] ), 
	.D(FE_PHN1968_n2748), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][5]  (.Q(\ram[135][5] ), 
	.D(FE_PHN5727_n2747), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][4]  (.Q(\ram[135][4] ), 
	.D(FE_PHN3035_n2746), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][3]  (.Q(\ram[135][3] ), 
	.D(FE_PHN1229_n2745), 
	.CK(clk_m__L3_N21));
   QDFFEHD \ram_reg[135][2]  (.Q(\ram[135][2] ), 
	.D(FE_PHN533_n2744), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[135][1]  (.Q(\ram[135][1] ), 
	.D(FE_PHN5689_n2743), 
	.CK(clk_m__L3_N24));
   QDFFEHD \ram_reg[135][0]  (.Q(\ram[135][0] ), 
	.D(FE_PHN1821_n2742), 
	.CK(clk_m__L3_N97));
   QDFFEHD \ram_reg[131][15]  (.Q(\ram[131][15] ), 
	.D(FE_PHN2472_n2693), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][14]  (.Q(\ram[131][14] ), 
	.D(FE_PHN3101_n2692), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][13]  (.Q(\ram[131][13] ), 
	.D(FE_PHN563_n2691), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][12]  (.Q(\ram[131][12] ), 
	.D(FE_PHN2052_n2690), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[131][11]  (.Q(\ram[131][11] ), 
	.D(FE_PHN1906_n2689), 
	.CK(clk_m__L3_N91));
   QDFFEHD \ram_reg[131][10]  (.Q(\ram[131][10] ), 
	.D(FE_PHN2176_n2688), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[131][9]  (.Q(\ram[131][9] ), 
	.D(FE_PHN1227_n2687), 
	.CK(clk_m__L3_N90));
   QDFFEHD \ram_reg[131][8]  (.Q(\ram[131][8] ), 
	.D(FE_PHN1776_n2686), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[131][7]  (.Q(\ram[131][7] ), 
	.D(FE_PHN1152_n2685), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[131][6]  (.Q(\ram[131][6] ), 
	.D(FE_PHN1263_n2684), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][5]  (.Q(\ram[131][5] ), 
	.D(FE_PHN575_n2683), 
	.CK(clk_m__L3_N20));
   QDFFEHD \ram_reg[131][4]  (.Q(\ram[131][4] ), 
	.D(FE_PHN1072_n2682), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][3]  (.Q(\ram[131][3] ), 
	.D(FE_PHN1123_n2681), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][2]  (.Q(\ram[131][2] ), 
	.D(FE_PHN1340_n2680), 
	.CK(clk_m__L3_N96));
   QDFFEHD \ram_reg[131][1]  (.Q(\ram[131][1] ), 
	.D(FE_PHN1190_n2679), 
	.CK(clk_m__L3_N23));
   QDFFEHD \ram_reg[131][0]  (.Q(\ram[131][0] ), 
	.D(FE_PHN788_n2678), 
	.CK(clk_m__L3_N98));
   QDFFEHD \ram_reg[127][15]  (.Q(\ram[127][15] ), 
	.D(FE_PHN2647_n2629), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[127][14]  (.Q(\ram[127][14] ), 
	.D(FE_PHN6667_n2628), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[127][13]  (.Q(\ram[127][13] ), 
	.D(FE_PHN2198_n2627), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[127][12]  (.Q(\ram[127][12] ), 
	.D(FE_PHN5751_n2626), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][11]  (.Q(\ram[127][11] ), 
	.D(FE_PHN6681_n2625), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][10]  (.Q(\ram[127][10] ), 
	.D(FE_PHN5755_n2624), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][9]  (.Q(\ram[127][9] ), 
	.D(FE_PHN4486_n2623), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[127][8]  (.Q(\ram[127][8] ), 
	.D(FE_PHN5700_n2622), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][7]  (.Q(\ram[127][7] ), 
	.D(FE_PHN4353_n2621), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][6]  (.Q(\ram[127][6] ), 
	.D(FE_PHN1238_n2620), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[127][5]  (.Q(\ram[127][5] ), 
	.D(FE_PHN4901_n2619), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][4]  (.Q(\ram[127][4] ), 
	.D(FE_PHN5728_n2618), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[127][3]  (.Q(\ram[127][3] ), 
	.D(FE_PHN1494_n2617), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[127][2]  (.Q(\ram[127][2] ), 
	.D(FE_PHN5667_n2616), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[127][1]  (.Q(\ram[127][1] ), 
	.D(FE_PHN5701_n2615), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[127][0]  (.Q(\ram[127][0] ), 
	.D(FE_PHN6697_n2614), 
	.CK(clk_m__L3_N156));
   QDFFEHD \ram_reg[123][15]  (.Q(\ram[123][15] ), 
	.D(FE_PHN2896_n2565), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][14]  (.Q(\ram[123][14] ), 
	.D(FE_PHN4694_n2564), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][13]  (.Q(\ram[123][13] ), 
	.D(FE_PHN1462_n2563), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[123][12]  (.Q(\ram[123][12] ), 
	.D(FE_PHN2408_n2562), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][11]  (.Q(\ram[123][11] ), 
	.D(FE_PHN2877_n2561), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[123][10]  (.Q(\ram[123][10] ), 
	.D(FE_PHN2644_n2560), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[123][9]  (.Q(\ram[123][9] ), 
	.D(FE_PHN2428_n2559), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[123][8]  (.Q(\ram[123][8] ), 
	.D(FE_PHN2171_n2558), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[123][7]  (.Q(\ram[123][7] ), 
	.D(FE_PHN1430_n2557), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[123][6]  (.Q(\ram[123][6] ), 
	.D(FE_PHN1997_n2556), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[123][5]  (.Q(\ram[123][5] ), 
	.D(FE_PHN2412_n2555), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[123][4]  (.Q(\ram[123][4] ), 
	.D(FE_PHN4564_n2554), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[123][3]  (.Q(\ram[123][3] ), 
	.D(FE_PHN592_n2553), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[123][2]  (.Q(\ram[123][2] ), 
	.D(FE_PHN1973_n2552), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[123][1]  (.Q(\ram[123][1] ), 
	.D(FE_PHN2174_n2551), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[123][0]  (.Q(\ram[123][0] ), 
	.D(FE_PHN2319_n2550), 
	.CK(clk_m__L3_N152));
   QDFFEHD \ram_reg[119][15]  (.Q(\ram[119][15] ), 
	.D(FE_PHN2632_n2501), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[119][14]  (.Q(\ram[119][14] ), 
	.D(FE_PHN2736_n2500), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][13]  (.Q(\ram[119][13] ), 
	.D(FE_PHN3091_n2499), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[119][12]  (.Q(\ram[119][12] ), 
	.D(FE_PHN1499_n2498), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[119][11]  (.Q(\ram[119][11] ), 
	.D(FE_PHN2119_n2497), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][10]  (.Q(\ram[119][10] ), 
	.D(FE_PHN1701_n2496), 
	.CK(clk_m__L3_N151));
   QDFFEHD \ram_reg[119][9]  (.Q(\ram[119][9] ), 
	.D(FE_PHN2510_n2495), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][8]  (.Q(\ram[119][8] ), 
	.D(FE_PHN1452_n2494), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][7]  (.Q(\ram[119][7] ), 
	.D(FE_PHN1041_n2493), 
	.CK(clk_m__L3_N153));
   QDFFEHD \ram_reg[119][6]  (.Q(\ram[119][6] ), 
	.D(FE_PHN2187_n2492), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][5]  (.Q(\ram[119][5] ), 
	.D(FE_PHN1225_n2491), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[119][4]  (.Q(\ram[119][4] ), 
	.D(FE_PHN1453_n2490), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][3]  (.Q(\ram[119][3] ), 
	.D(FE_PHN292_n2489), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][2]  (.Q(\ram[119][2] ), 
	.D(FE_PHN798_n2488), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[119][1]  (.Q(\ram[119][1] ), 
	.D(FE_PHN2524_n2487), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[119][0]  (.Q(\ram[119][0] ), 
	.D(FE_PHN1451_n2486), 
	.CK(clk_m__L3_N157));
   QDFFEHD \ram_reg[115][15]  (.Q(\ram[115][15] ), 
	.D(FE_PHN4317_n2437), 
	.CK(clk_m__L3_N124));
   QDFFEHD \ram_reg[115][14]  (.Q(\ram[115][14] ), 
	.D(FE_PHN756_n2436), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[115][13]  (.Q(\ram[115][13] ), 
	.D(FE_PHN408_n2435), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[115][12]  (.Q(\ram[115][12] ), 
	.D(FE_PHN6657_n2434), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][11]  (.Q(\ram[115][11] ), 
	.D(FE_PHN4280_n2433), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][10]  (.Q(\ram[115][10] ), 
	.D(FE_PHN4321_n2432), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[115][9]  (.Q(\ram[115][9] ), 
	.D(FE_PHN4062_n2431), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[115][8]  (.Q(\ram[115][8] ), 
	.D(FE_PHN4422_n2430), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][7]  (.Q(\ram[115][7] ), 
	.D(FE_PHN6556_n2429), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][6]  (.Q(\ram[115][6] ), 
	.D(FE_PHN5650_n2428), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[115][5]  (.Q(\ram[115][5] ), 
	.D(FE_PHN6670_n2427), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[115][4]  (.Q(\ram[115][4] ), 
	.D(FE_PHN6655_n2426), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[115][3]  (.Q(\ram[115][3] ), 
	.D(FE_PHN6647_n2425), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[115][2]  (.Q(\ram[115][2] ), 
	.D(FE_PHN5720_n2424), 
	.CK(clk_m__L3_N154));
   QDFFEHD \ram_reg[115][1]  (.Q(\ram[115][1] ), 
	.D(FE_PHN5714_n2423), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[115][0]  (.Q(\ram[115][0] ), 
	.D(FE_PHN4869_n2422), 
	.CK(clk_m__L3_N155));
   QDFFEHD \ram_reg[111][15]  (.Q(\ram[111][15] ), 
	.D(FE_PHN1814_n2373), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][14]  (.Q(\ram[111][14] ), 
	.D(FE_PHN1944_n2372), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][13]  (.Q(\ram[111][13] ), 
	.D(FE_PHN1860_n2371), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][12]  (.Q(\ram[111][12] ), 
	.D(FE_PHN2870_n2370), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][11]  (.Q(\ram[111][11] ), 
	.D(FE_PHN2575_n2369), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][10]  (.Q(\ram[111][10] ), 
	.D(FE_PHN2716_n2368), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][9]  (.Q(\ram[111][9] ), 
	.D(FE_PHN2714_n2367), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][8]  (.Q(\ram[111][8] ), 
	.D(FE_PHN2659_n2366), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][7]  (.Q(\ram[111][7] ), 
	.D(FE_PHN428_n2365), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[111][6]  (.Q(\ram[111][6] ), 
	.D(FE_PHN1623_n2364), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][5]  (.Q(\ram[111][5] ), 
	.D(FE_PHN1312_n2363), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][4]  (.Q(\ram[111][4] ), 
	.D(FE_PHN2766_n2362), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][3]  (.Q(\ram[111][3] ), 
	.D(FE_PHN409_n2361), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[111][2]  (.Q(\ram[111][2] ), 
	.D(FE_PHN3200_n2360), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][1]  (.Q(\ram[111][1] ), 
	.D(FE_PHN2704_n2359), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[111][0]  (.Q(\ram[111][0] ), 
	.D(FE_PHN3136_n2358), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[107][15]  (.Q(\ram[107][15] ), 
	.D(FE_PHN2655_n2309), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][14]  (.Q(\ram[107][14] ), 
	.D(FE_PHN1173_n2308), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[107][13]  (.Q(\ram[107][13] ), 
	.D(FE_PHN820_n2307), 
	.CK(clk_m__L3_N73));
   QDFFEHD \ram_reg[107][12]  (.Q(\ram[107][12] ), 
	.D(FE_PHN2930_n2306), 
	.CK(clk_m__L3_N72));
   QDFFEHD \ram_reg[107][11]  (.Q(\ram[107][11] ), 
	.D(FE_PHN1678_n2305), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[107][10]  (.Q(\ram[107][10] ), 
	.D(FE_PHN3062_n2304), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][9]  (.Q(\ram[107][9] ), 
	.D(FE_PHN1616_n2303), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][8]  (.Q(\ram[107][8] ), 
	.D(FE_PHN2306_n2302), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[107][7]  (.Q(\ram[107][7] ), 
	.D(FE_PHN1875_n2301), 
	.CK(clk_m__L3_N82));
   QDFFEHD \ram_reg[107][6]  (.Q(\ram[107][6] ), 
	.D(FE_PHN1206_n2300), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][5]  (.Q(\ram[107][5] ), 
	.D(FE_PHN415_n2299), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[107][4]  (.Q(\ram[107][4] ), 
	.D(FE_PHN1978_n2298), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][3]  (.Q(\ram[107][3] ), 
	.D(FE_PHN4672_n2297), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[107][2]  (.Q(\ram[107][2] ), 
	.D(FE_PHN1262_n2296), 
	.CK(clk_m__L3_N69));
   QDFFEHD \ram_reg[107][1]  (.Q(\ram[107][1] ), 
	.D(FE_PHN1854_n2295), 
	.CK(clk_m__L3_N83));
   QDFFEHD \ram_reg[107][0]  (.Q(\ram[107][0] ), 
	.D(FE_PHN349_n2294), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[103][15]  (.Q(\ram[103][15] ), 
	.D(FE_PHN400_n2245), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[103][14]  (.Q(\ram[103][14] ), 
	.D(FE_PHN1596_n2244), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[103][13]  (.Q(\ram[103][13] ), 
	.D(FE_PHN970_n2243), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][12]  (.Q(\ram[103][12] ), 
	.D(FE_PHN2650_n2242), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][11]  (.Q(\ram[103][11] ), 
	.D(FE_PHN2652_n2241), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][10]  (.Q(\ram[103][10] ), 
	.D(FE_PHN3016_n2240), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][9]  (.Q(\ram[103][9] ), 
	.D(FE_PHN2203_n2239), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][8]  (.Q(\ram[103][8] ), 
	.D(FE_PHN622_n2238), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][7]  (.Q(\ram[103][7] ), 
	.D(FE_PHN2034_n2237), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[103][6]  (.Q(\ram[103][6] ), 
	.D(FE_PHN430_n2236), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][5]  (.Q(\ram[103][5] ), 
	.D(FE_PHN2777_n2235), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][4]  (.Q(\ram[103][4] ), 
	.D(FE_PHN2305_n2234), 
	.CK(clk_m__L3_N71));
   QDFFEHD \ram_reg[103][3]  (.Q(\ram[103][3] ), 
	.D(FE_PHN1564_n2233), 
	.CK(clk_m__L3_N81));
   QDFFEHD \ram_reg[103][2]  (.Q(\ram[103][2] ), 
	.D(FE_PHN2235_n2232), 
	.CK(clk_m__L3_N87));
   QDFFEHD \ram_reg[103][1]  (.Q(\ram[103][1] ), 
	.D(FE_PHN1149_n2231), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[103][0]  (.Q(\ram[103][0] ), 
	.D(FE_PHN1369_n2230), 
	.CK(clk_m__L3_N86));
   QDFFEHD \ram_reg[99][15]  (.Q(\ram[99][15] ), 
	.D(FE_PHN5737_n2181), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[99][14]  (.Q(\ram[99][14] ), 
	.D(FE_PHN4922_n2180), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][13]  (.Q(\ram[99][13] ), 
	.D(FE_PHN4785_n2179), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[99][12]  (.Q(\ram[99][12] ), 
	.D(FE_PHN3435_n2178), 
	.CK(clk_m__L3_N70));
   QDFFEHD \ram_reg[99][11]  (.Q(\ram[99][11] ), 
	.D(FE_PHN5666_n2177), 
	.CK(clk_m__L3_N84));
   QDFFEHD \ram_reg[99][10]  (.Q(\ram[99][10] ), 
	.D(FE_PHN5662_n2176), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][9]  (.Q(\ram[99][9] ), 
	.D(FE_PHN6694_n2175), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][8]  (.Q(\ram[99][8] ), 
	.D(FE_PHN242_n2174), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][7]  (.Q(\ram[99][7] ), 
	.D(FE_PHN715_n2173), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[99][6]  (.Q(\ram[99][6] ), 
	.D(FE_PHN5736_n2172), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][5]  (.Q(\ram[99][5] ), 
	.D(FE_PHN5652_n2171), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][4]  (.Q(\ram[99][4] ), 
	.D(FE_PHN6660_n2170), 
	.CK(clk_m__L3_N85));
   QDFFEHD \ram_reg[99][3]  (.Q(\ram[99][3] ), 
	.D(FE_PHN6662_n2169), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[99][2]  (.Q(\ram[99][2] ), 
	.D(FE_PHN6644_n2168), 
	.CK(clk_m__L3_N88));
   QDFFEHD \ram_reg[99][1]  (.Q(\ram[99][1] ), 
	.D(FE_PHN6707_n2167), 
	.CK(clk_m__L3_N80));
   QDFFEHD \ram_reg[99][0]  (.Q(\ram[99][0] ), 
	.D(FE_PHN6708_n2166), 
	.CK(clk_m__L3_N79));
   QDFFEHD \ram_reg[95][15]  (.Q(\ram[95][15] ), 
	.D(FE_PHN2599_n2117), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][14]  (.Q(\ram[95][14] ), 
	.D(FE_PHN2807_n2116), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[95][13]  (.Q(\ram[95][13] ), 
	.D(FE_PHN2607_n2115), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][12]  (.Q(\ram[95][12] ), 
	.D(FE_PHN1841_n2114), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[95][11]  (.Q(\ram[95][11] ), 
	.D(FE_PHN2737_n2113), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[95][10]  (.Q(\ram[95][10] ), 
	.D(FE_PHN3100_n2112), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][9]  (.Q(\ram[95][9] ), 
	.D(FE_PHN2980_n2111), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][8]  (.Q(\ram[95][8] ), 
	.D(FE_PHN2011_n2110), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[95][7]  (.Q(\ram[95][7] ), 
	.D(FE_PHN2805_n2109), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][6]  (.Q(\ram[95][6] ), 
	.D(FE_PHN1808_n2108), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[95][5]  (.Q(\ram[95][5] ), 
	.D(FE_PHN796_n2107), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[95][4]  (.Q(\ram[95][4] ), 
	.D(FE_PHN1921_n2106), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][3]  (.Q(\ram[95][3] ), 
	.D(FE_PHN2969_n2105), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[95][2]  (.Q(\ram[95][2] ), 
	.D(FE_PHN3221_n2104), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][1]  (.Q(\ram[95][1] ), 
	.D(FE_PHN2920_n2103), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[95][0]  (.Q(\ram[95][0] ), 
	.D(FE_PHN2758_n2102), 
	.CK(clk_m__L3_N166));
   QDFFEHD \ram_reg[91][15]  (.Q(\ram[91][15] ), 
	.D(FE_PHN3046_n2053), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][14]  (.Q(\ram[91][14] ), 
	.D(FE_PHN3102_n2052), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[91][13]  (.Q(\ram[91][13] ), 
	.D(FE_PHN3006_n2051), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][12]  (.Q(\ram[91][12] ), 
	.D(FE_PHN2794_n2050), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][11]  (.Q(\ram[91][11] ), 
	.D(FE_PHN2339_n2049), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][10]  (.Q(\ram[91][10] ), 
	.D(FE_PHN2909_n2048), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][9]  (.Q(\ram[91][9] ), 
	.D(FE_PHN2442_n2047), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][8]  (.Q(\ram[91][8] ), 
	.D(FE_PHN1326_n2046), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][7]  (.Q(\ram[91][7] ), 
	.D(FE_PHN1861_n2045), 
	.CK(clk_m__L3_N160));
   QDFFEHD \ram_reg[91][6]  (.Q(\ram[91][6] ), 
	.D(FE_PHN2459_n2044), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][5]  (.Q(\ram[91][5] ), 
	.D(FE_PHN2876_n2043), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][4]  (.Q(\ram[91][4] ), 
	.D(FE_PHN980_n2042), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[91][3]  (.Q(\ram[91][3] ), 
	.D(FE_PHN3071_n2041), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][2]  (.Q(\ram[91][2] ), 
	.D(FE_PHN2555_n2040), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][1]  (.Q(\ram[91][1] ), 
	.D(FE_PHN2660_n2039), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[91][0]  (.Q(\ram[91][0] ), 
	.D(FE_PHN2676_n2038), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[87][15]  (.Q(\ram[87][15] ), 
	.D(FE_PHN1656_n1989), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][14]  (.Q(\ram[87][14] ), 
	.D(FE_PHN2427_n1988), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][13]  (.Q(\ram[87][13] ), 
	.D(FE_PHN2377_n1987), 
	.CK(clk_m__L3_N163));
   QDFFEHD \ram_reg[87][12]  (.Q(\ram[87][12] ), 
	.D(FE_PHN1887_n1986), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[87][11]  (.Q(\ram[87][11] ), 
	.D(FE_PHN1431_n1985), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][10]  (.Q(\ram[87][10] ), 
	.D(FE_PHN2994_n1984), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][9]  (.Q(\ram[87][9] ), 
	.D(FE_PHN2462_n1983), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][8]  (.Q(\ram[87][8] ), 
	.D(FE_PHN1328_n1982), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][7]  (.Q(\ram[87][7] ), 
	.D(FE_PHN2083_n1981), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][6]  (.Q(\ram[87][6] ), 
	.D(FE_PHN983_n1980), 
	.CK(clk_m__L3_N167));
   QDFFEHD \ram_reg[87][5]  (.Q(\ram[87][5] ), 
	.D(FE_PHN1939_n1979), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][4]  (.Q(\ram[87][4] ), 
	.D(FE_PHN3190_n1978), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][3]  (.Q(\ram[87][3] ), 
	.D(FE_PHN2908_n1977), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][2]  (.Q(\ram[87][2] ), 
	.D(FE_PHN1112_n1976), 
	.CK(clk_m__L3_N162));
   QDFFEHD \ram_reg[87][1]  (.Q(\ram[87][1] ), 
	.D(FE_PHN2434_n1975), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[87][0]  (.Q(\ram[87][0] ), 
	.D(FE_PHN2348_n1974), 
	.CK(clk_m__L3_N148));
   QDFFEHD \ram_reg[83][15]  (.Q(\ram[83][15] ), 
	.D(FE_PHN1888_n1925), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][14]  (.Q(\ram[83][14] ), 
	.D(FE_PHN2653_n1924), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][13]  (.Q(\ram[83][13] ), 
	.D(FE_PHN1073_n1923), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][12]  (.Q(\ram[83][12] ), 
	.D(FE_PHN3840_n1922), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][11]  (.Q(\ram[83][11] ), 
	.D(FE_PHN4186_n1921), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[83][10]  (.Q(\ram[83][10] ), 
	.D(FE_PHN4664_n1920), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][9]  (.Q(\ram[83][9] ), 
	.D(FE_PHN4250_n1919), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][8]  (.Q(\ram[83][8] ), 
	.D(FE_PHN4476_n1918), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[83][7]  (.Q(\ram[83][7] ), 
	.D(FE_PHN2906_n1917), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][6]  (.Q(\ram[83][6] ), 
	.D(FE_PHN4363_n1916), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][5]  (.Q(\ram[83][5] ), 
	.D(FE_PHN2202_n1915), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[83][4]  (.Q(\ram[83][4] ), 
	.D(FE_PHN2964_n1914), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[83][3]  (.Q(\ram[83][3] ), 
	.D(FE_PHN5765_n1913), 
	.CK(clk_m__L3_N164));
   QDFFEHD \ram_reg[83][2]  (.Q(\ram[83][2] ), 
	.D(FE_PHN2698_n1912), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[83][1]  (.Q(\ram[83][1] ), 
	.D(FE_PHN4239_n1911), 
	.CK(clk_m__L3_N150));
   QDFFEHD \ram_reg[83][0]  (.Q(\ram[83][0] ), 
	.D(FE_PHN1106_n1910), 
	.CK(clk_m__L3_N149));
   QDFFEHD \ram_reg[79][15]  (.Q(\ram[79][15] ), 
	.D(FE_PHN617_n1861), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][14]  (.Q(\ram[79][14] ), 
	.D(FE_PHN1903_n1860), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][13]  (.Q(\ram[79][13] ), 
	.D(FE_PHN3023_n1859), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][12]  (.Q(\ram[79][12] ), 
	.D(FE_PHN1373_n1858), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][11]  (.Q(\ram[79][11] ), 
	.D(FE_PHN2381_n1857), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][10]  (.Q(\ram[79][10] ), 
	.D(FE_PHN3019_n1856), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[79][9]  (.Q(\ram[79][9] ), 
	.D(FE_PHN1042_n1855), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][8]  (.Q(\ram[79][8] ), 
	.D(FE_PHN1459_n1854), 
	.CK(clk_m__L3_N59));
   QDFFEHD \ram_reg[79][7]  (.Q(\ram[79][7] ), 
	.D(FE_PHN1671_n1853), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[79][6]  (.Q(\ram[79][6] ), 
	.D(FE_PHN1848_n1852), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][5]  (.Q(\ram[79][5] ), 
	.D(FE_PHN950_n1851), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][4]  (.Q(\ram[79][4] ), 
	.D(FE_PHN3097_n1850), 
	.CK(clk_m__L3_N65));
   QDFFEHD \ram_reg[79][3]  (.Q(\ram[79][3] ), 
	.D(FE_PHN1222_n1849), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[79][2]  (.Q(\ram[79][2] ), 
	.D(FE_PHN2847_n1848), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[79][1]  (.Q(\ram[79][1] ), 
	.D(FE_PHN1349_n1847), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[79][0]  (.Q(\ram[79][0] ), 
	.D(FE_PHN1286_n1846), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[75][15]  (.Q(\ram[75][15] ), 
	.D(FE_PHN1481_n1797), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][14]  (.Q(\ram[75][14] ), 
	.D(FE_PHN2298_n1796), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][13]  (.Q(\ram[75][13] ), 
	.D(FE_PHN243_n1795), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][12]  (.Q(\ram[75][12] ), 
	.D(FE_PHN2200_n1794), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][11]  (.Q(\ram[75][11] ), 
	.D(FE_PHN1775_n1793), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][10]  (.Q(\ram[75][10] ), 
	.D(FE_PHN347_n1792), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][9]  (.Q(\ram[75][9] ), 
	.D(FE_PHN2667_n1791), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][8]  (.Q(\ram[75][8] ), 
	.D(FE_PHN545_n1790), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[75][7]  (.Q(\ram[75][7] ), 
	.D(FE_PHN2725_n1789), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][6]  (.Q(\ram[75][6] ), 
	.D(FE_PHN2271_n1788), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][5]  (.Q(\ram[75][5] ), 
	.D(FE_PHN3039_n1787), 
	.CK(clk_m__L3_N68));
   QDFFEHD \ram_reg[75][4]  (.Q(\ram[75][4] ), 
	.D(FE_PHN2635_n1786), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][3]  (.Q(\ram[75][3] ), 
	.D(FE_PHN1054_n1785), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[75][2]  (.Q(\ram[75][2] ), 
	.D(FE_PHN3055_n1784), 
	.CK(clk_m__L3_N67));
   QDFFEHD \ram_reg[75][1]  (.Q(\ram[75][1] ), 
	.D(FE_PHN1533_n1783), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[75][0]  (.Q(\ram[75][0] ), 
	.D(FE_PHN316_n1782), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[71][15]  (.Q(\ram[71][15] ), 
	.D(FE_PHN1379_n1733), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][14]  (.Q(\ram[71][14] ), 
	.D(FE_PHN1150_n1732), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][13]  (.Q(\ram[71][13] ), 
	.D(FE_PHN3085_n1731), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][12]  (.Q(\ram[71][12] ), 
	.D(FE_PHN389_n1730), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][11]  (.Q(\ram[71][11] ), 
	.D(FE_PHN1889_n1729), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][10]  (.Q(\ram[71][10] ), 
	.D(FE_PHN1249_n1728), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][9]  (.Q(\ram[71][9] ), 
	.D(FE_PHN2957_n1727), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][8]  (.Q(\ram[71][8] ), 
	.D(FE_PHN3038_n1726), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[71][7]  (.Q(\ram[71][7] ), 
	.D(FE_PHN2948_n1725), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][6]  (.Q(\ram[71][6] ), 
	.D(FE_PHN1758_n1724), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][5]  (.Q(\ram[71][5] ), 
	.D(FE_PHN2551_n1723), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][4]  (.Q(\ram[71][4] ), 
	.D(FE_PHN605_n1722), 
	.CK(clk_m__L3_N64));
   QDFFEHD \ram_reg[71][3]  (.Q(\ram[71][3] ), 
	.D(FE_PHN1580_n1721), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[71][2]  (.Q(\ram[71][2] ), 
	.D(FE_PHN760_n1720), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[71][1]  (.Q(\ram[71][1] ), 
	.D(FE_PHN2755_n1719), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[71][0]  (.Q(\ram[71][0] ), 
	.D(FE_PHN1016_n1718), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[67][15]  (.Q(\ram[67][15] ), 
	.D(FE_PHN992_n1669), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[67][14]  (.Q(\ram[67][14] ), 
	.D(FE_PHN1257_n1668), 
	.CK(clk_m__L3_N75));
   QDFFEHD \ram_reg[67][13]  (.Q(\ram[67][13] ), 
	.D(FE_PHN911_n1667), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[67][12]  (.Q(\ram[67][12] ), 
	.D(FE_PHN1240_n1666), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[67][11]  (.Q(\ram[67][11] ), 
	.D(FE_PHN2393_n1665), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][10]  (.Q(\ram[67][10] ), 
	.D(FE_PHN1835_n1664), 
	.CK(clk_m__L3_N78));
   QDFFEHD \ram_reg[67][9]  (.Q(\ram[67][9] ), 
	.D(n1663), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[67][8]  (.Q(\ram[67][8] ), 
	.D(FE_PHN2516_n1662), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][7]  (.Q(\ram[67][7] ), 
	.D(FE_PHN1124_n1661), 
	.CK(clk_m__L3_N63));
   QDFFEHD \ram_reg[67][6]  (.Q(\ram[67][6] ), 
	.D(FE_PHN2246_n1660), 
	.CK(clk_m__L3_N61));
   QDFFEHD \ram_reg[67][5]  (.Q(\ram[67][5] ), 
	.D(FE_PHN2044_n1659), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][4]  (.Q(\ram[67][4] ), 
	.D(FE_PHN2151_n1658), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][3]  (.Q(\ram[67][3] ), 
	.D(FE_PHN748_n1657), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[67][2]  (.Q(\ram[67][2] ), 
	.D(FE_PHN559_n1656), 
	.CK(clk_m__L3_N62));
   QDFFEHD \ram_reg[67][1]  (.Q(\ram[67][1] ), 
	.D(FE_PHN1581_n1655), 
	.CK(clk_m__L3_N76));
   QDFFEHD \ram_reg[67][0]  (.Q(\ram[67][0] ), 
	.D(FE_PHN2617_n1654), 
	.CK(clk_m__L3_N77));
   QDFFEHD \ram_reg[63][15]  (.Q(\ram[63][15] ), 
	.D(FE_PHN1986_n1605), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][14]  (.Q(\ram[63][14] ), 
	.D(FE_PHN734_n1604), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][13]  (.Q(\ram[63][13] ), 
	.D(FE_PHN1170_n1603), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][12]  (.Q(\ram[63][12] ), 
	.D(FE_PHN2854_n1602), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[63][11]  (.Q(\ram[63][11] ), 
	.D(FE_PHN3184_n1601), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[63][10]  (.Q(\ram[63][10] ), 
	.D(FE_PHN3047_n1600), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][9]  (.Q(\ram[63][9] ), 
	.D(FE_PHN1675_n1599), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[63][8]  (.Q(\ram[63][8] ), 
	.D(FE_PHN2272_n1598), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][7]  (.Q(\ram[63][7] ), 
	.D(FE_PHN774_n1597), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[63][6]  (.Q(\ram[63][6] ), 
	.D(FE_PHN2852_n1596), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][5]  (.Q(\ram[63][5] ), 
	.D(n1595), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][4]  (.Q(\ram[63][4] ), 
	.D(FE_PHN2121_n1594), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[63][3]  (.Q(\ram[63][3] ), 
	.D(FE_PHN3125_n1593), 
	.CK(clk_m__L3_N169));
   QDFFEHD \ram_reg[63][2]  (.Q(\ram[63][2] ), 
	.D(FE_PHN2291_n1592), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[63][1]  (.Q(\ram[63][1] ), 
	.D(FE_PHN2292_n1591), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[63][0]  (.Q(\ram[63][0] ), 
	.D(FE_PHN2013_n1590), 
	.CK(clk_m__L3_N175));
   QDFFEHD \ram_reg[59][15]  (.Q(\ram[59][15] ), 
	.D(FE_PHN1409_n1541), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][14]  (.Q(\ram[59][14] ), 
	.D(FE_PHN3009_n1540), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][13]  (.Q(\ram[59][13] ), 
	.D(FE_PHN1868_n1539), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][12]  (.Q(\ram[59][12] ), 
	.D(FE_PHN2574_n1538), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[59][11]  (.Q(\ram[59][11] ), 
	.D(FE_PHN2064_n1537), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][10]  (.Q(\ram[59][10] ), 
	.D(FE_PHN3220_n1536), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][9]  (.Q(\ram[59][9] ), 
	.D(FE_PHN1836_n1535), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][8]  (.Q(\ram[59][8] ), 
	.D(FE_PHN2188_n1534), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][7]  (.Q(\ram[59][7] ), 
	.D(FE_PHN2903_n1533), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][6]  (.Q(\ram[59][6] ), 
	.D(FE_PHN2735_n1532), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][5]  (.Q(\ram[59][5] ), 
	.D(FE_PHN2833_n1531), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[59][4]  (.Q(\ram[59][4] ), 
	.D(FE_PHN2340_n1530), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[59][3]  (.Q(\ram[59][3] ), 
	.D(FE_PHN3140_n1529), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[59][2]  (.Q(\ram[59][2] ), 
	.D(FE_PHN990_n1528), 
	.CK(clk_m__L3_N172));
   QDFFEHD \ram_reg[59][1]  (.Q(\ram[59][1] ), 
	.D(FE_PHN1967_n1527), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[59][0]  (.Q(\ram[59][0] ), 
	.D(FE_PHN823_n1526), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[55][15]  (.Q(\ram[55][15] ), 
	.D(FE_PHN1763_n1477), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][14]  (.Q(\ram[55][14] ), 
	.D(FE_PHN2808_n1476), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][13]  (.Q(\ram[55][13] ), 
	.D(FE_PHN751_n1475), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][12]  (.Q(\ram[55][12] ), 
	.D(FE_PHN2527_n1474), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[55][11]  (.Q(\ram[55][11] ), 
	.D(FE_PHN1826_n1473), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][10]  (.Q(\ram[55][10] ), 
	.D(FE_PHN2881_n1472), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][9]  (.Q(\ram[55][9] ), 
	.D(FE_PHN1524_n1471), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][8]  (.Q(\ram[55][8] ), 
	.D(FE_PHN3096_n1470), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][7]  (.Q(\ram[55][7] ), 
	.D(FE_PHN2449_n1469), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][6]  (.Q(\ram[55][6] ), 
	.D(FE_PHN2986_n1468), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][5]  (.Q(\ram[55][5] ), 
	.D(FE_PHN2711_n1467), 
	.CK(clk_m__L3_N170));
   QDFFEHD \ram_reg[55][4]  (.Q(\ram[55][4] ), 
	.D(FE_PHN1338_n1466), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][3]  (.Q(\ram[55][3] ), 
	.D(FE_PHN2546_n1465), 
	.CK(clk_m__L3_N173));
   QDFFEHD \ram_reg[55][2]  (.Q(\ram[55][2] ), 
	.D(FE_PHN2469_n1464), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][1]  (.Q(\ram[55][1] ), 
	.D(FE_PHN2757_n1463), 
	.CK(clk_m__L3_N174));
   QDFFEHD \ram_reg[55][0]  (.Q(\ram[55][0] ), 
	.D(FE_PHN2549_n1462), 
	.CK(clk_m__L3_N158));
   QDFFEHD \ram_reg[51][15]  (.Q(\ram[51][15] ), 
	.D(FE_PHN3058_n1413), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[51][14]  (.Q(\ram[51][14] ), 
	.D(FE_PHN1829_n1412), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][13]  (.Q(\ram[51][13] ), 
	.D(FE_PHN1330_n1411), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][12]  (.Q(\ram[51][12] ), 
	.D(FE_PHN1897_n1410), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[51][11]  (.Q(\ram[51][11] ), 
	.D(FE_PHN1291_n1409), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][10]  (.Q(\ram[51][10] ), 
	.D(FE_PHN981_n1408), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][9]  (.Q(\ram[51][9] ), 
	.D(FE_PHN2924_n1407), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[51][8]  (.Q(\ram[51][8] ), 
	.D(FE_PHN436_n1406), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][7]  (.Q(\ram[51][7] ), 
	.D(FE_PHN3156_n1405), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[51][6]  (.Q(\ram[51][6] ), 
	.D(FE_PHN2684_n1404), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[51][5]  (.Q(\ram[51][5] ), 
	.D(FE_PHN2504_n1403), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][4]  (.Q(\ram[51][4] ), 
	.D(FE_PHN2204_n1402), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][3]  (.Q(\ram[51][3] ), 
	.D(FE_PHN3196_n1401), 
	.CK(clk_m__L3_N159));
   QDFFEHD \ram_reg[51][2]  (.Q(\ram[51][2] ), 
	.D(FE_PHN2505_n1400), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[51][1]  (.Q(\ram[51][1] ), 
	.D(FE_PHN2785_n1399), 
	.CK(clk_m__L3_N177));
   QDFFEHD \ram_reg[51][0]  (.Q(\ram[51][0] ), 
	.D(FE_PHN2661_n1398), 
	.CK(clk_m__L3_N161));
   QDFFEHD \ram_reg[47][15]  (.Q(\ram[47][15] ), 
	.D(FE_PHN3063_n1349), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[47][14]  (.Q(\ram[47][14] ), 
	.D(FE_PHN1221_n1348), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][13]  (.Q(\ram[47][13] ), 
	.D(FE_PHN2547_n1347), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[47][12]  (.Q(\ram[47][12] ), 
	.D(FE_PHN2115_n1346), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][11]  (.Q(\ram[47][11] ), 
	.D(FE_PHN2451_n1345), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][10]  (.Q(\ram[47][10] ), 
	.D(FE_PHN2784_n1344), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][9]  (.Q(\ram[47][9] ), 
	.D(FE_PHN2525_n1343), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[47][8]  (.Q(\ram[47][8] ), 
	.D(FE_PHN2739_n1342), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[47][7]  (.Q(\ram[47][7] ), 
	.D(FE_PHN2780_n1341), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][6]  (.Q(\ram[47][6] ), 
	.D(FE_PHN1271_n1340), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][5]  (.Q(\ram[47][5] ), 
	.D(FE_PHN2032_n1339), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][4]  (.Q(\ram[47][4] ), 
	.D(FE_PHN2156_n1338), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][3]  (.Q(\ram[47][3] ), 
	.D(FE_PHN2767_n1337), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[47][2]  (.Q(\ram[47][2] ), 
	.D(FE_PHN2965_n1336), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][1]  (.Q(\ram[47][1] ), 
	.D(FE_PHN1495_n1335), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[47][0]  (.Q(\ram[47][0] ), 
	.D(FE_PHN1977_n1334), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[43][15]  (.Q(\ram[43][15] ), 
	.D(FE_PHN1993_n1285), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][14]  (.Q(\ram[43][14] ), 
	.D(FE_PHN2405_n1284), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[43][13]  (.Q(\ram[43][13] ), 
	.D(FE_PHN2519_n1283), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[43][12]  (.Q(\ram[43][12] ), 
	.D(FE_PHN1747_n1282), 
	.CK(clk_m__L3_N176));
   QDFFEHD \ram_reg[43][11]  (.Q(\ram[43][11] ), 
	.D(FE_PHN2938_n1281), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[43][10]  (.Q(\ram[43][10] ), 
	.D(FE_PHN2864_n1280), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][9]  (.Q(\ram[43][9] ), 
	.D(FE_PHN3170_n1279), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][8]  (.Q(\ram[43][8] ), 
	.D(FE_PHN2640_n1278), 
	.CK(clk_m__L3_N143));
   QDFFEHD \ram_reg[43][7]  (.Q(\ram[43][7] ), 
	.D(FE_PHN3160_n1277), 
	.CK(clk_m__L3_N171));
   QDFFEHD \ram_reg[43][6]  (.Q(\ram[43][6] ), 
	.D(FE_PHN1682_n1276), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[43][5]  (.Q(\ram[43][5] ), 
	.D(FE_PHN1799_n1275), 
	.CK(clk_m__L3_N168));
   QDFFEHD \ram_reg[43][4]  (.Q(\ram[43][4] ), 
	.D(FE_PHN2671_n1274), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[43][3]  (.Q(\ram[43][3] ), 
	.D(FE_PHN1501_n1273), 
	.CK(clk_m__L3_N139));
   QDFFEHD \ram_reg[43][2]  (.Q(\ram[43][2] ), 
	.D(FE_PHN2311_n1272), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[43][1]  (.Q(\ram[43][1] ), 
	.D(FE_PHN2945_n1271), 
	.CK(clk_m__L3_N146));
   QDFFEHD \ram_reg[43][0]  (.Q(\ram[43][0] ), 
	.D(FE_PHN2116_n1270), 
	.CK(clk_m__L3_N129));
   QDFFEHD \ram_reg[39][15]  (.Q(\ram[39][15] ), 
	.D(FE_PHN2251_n1221), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][14]  (.Q(\ram[39][14] ), 
	.D(FE_PHN2082_n1220), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[39][13]  (.Q(\ram[39][13] ), 
	.D(FE_PHN2473_n1219), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[39][12]  (.Q(\ram[39][12] ), 
	.D(FE_PHN1296_n1218), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[39][11]  (.Q(\ram[39][11] ), 
	.D(FE_PHN1311_n1217), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[39][10]  (.Q(\ram[39][10] ), 
	.D(FE_PHN2628_n1216), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][9]  (.Q(\ram[39][9] ), 
	.D(FE_PHN2705_n1215), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][8]  (.Q(\ram[39][8] ), 
	.D(FE_PHN1310_n1214), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[39][7]  (.Q(\ram[39][7] ), 
	.D(FE_PHN2935_n1213), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[39][6]  (.Q(\ram[39][6] ), 
	.D(FE_PHN3111_n1212), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[39][5]  (.Q(\ram[39][5] ), 
	.D(FE_PHN1394_n1211), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[39][4]  (.Q(\ram[39][4] ), 
	.D(FE_PHN2070_n1210), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[39][3]  (.Q(\ram[39][3] ), 
	.D(FE_PHN2029_n1209), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[39][2]  (.Q(\ram[39][2] ), 
	.D(FE_PHN2282_n1208), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[39][1]  (.Q(\ram[39][1] ), 
	.D(FE_PHN1496_n1207), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[39][0]  (.Q(\ram[39][0] ), 
	.D(FE_PHN4754_n1206), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[35][15]  (.Q(\ram[35][15] ), 
	.D(FE_PHN2391_n1157), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[35][14]  (.Q(\ram[35][14] ), 
	.D(FE_PHN2528_n1156), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][13]  (.Q(\ram[35][13] ), 
	.D(FE_PHN2669_n1155), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][12]  (.Q(\ram[35][12] ), 
	.D(FE_PHN5674_n1154), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][11]  (.Q(\ram[35][11] ), 
	.D(FE_PHN2604_n1153), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][10]  (.Q(\ram[35][10] ), 
	.D(FE_PHN937_n1152), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][9]  (.Q(\ram[35][9] ), 
	.D(FE_PHN2108_n1151), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[35][8]  (.Q(\ram[35][8] ), 
	.D(FE_PHN3093_n1150), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][7]  (.Q(\ram[35][7] ), 
	.D(FE_PHN2501_n1149), 
	.CK(clk_m__L3_N144));
   QDFFEHD \ram_reg[35][6]  (.Q(\ram[35][6] ), 
	.D(FE_PHN2645_n1148), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][5]  (.Q(\ram[35][5] ), 
	.D(FE_PHN2956_n1147), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][4]  (.Q(\ram[35][4] ), 
	.D(FE_PHN256_n1146), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][3]  (.Q(\ram[35][3] ), 
	.D(FE_PHN749_n1145), 
	.CK(clk_m__L3_N138));
   QDFFEHD \ram_reg[35][2]  (.Q(\ram[35][2] ), 
	.D(FE_PHN713_n1144), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][1]  (.Q(\ram[35][1] ), 
	.D(FE_PHN4556_n1143), 
	.CK(clk_m__L3_N147));
   QDFFEHD \ram_reg[35][0]  (.Q(\ram[35][0] ), 
	.D(FE_PHN5731_n1142), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[31][15]  (.Q(\ram[31][15] ), 
	.D(FE_PHN4977_n1093), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[31][14]  (.Q(\ram[31][14] ), 
	.D(FE_PHN1505_n1092), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][13]  (.Q(\ram[31][13] ), 
	.D(FE_PHN1998_n1091), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[31][12]  (.Q(\ram[31][12] ), 
	.D(FE_PHN4969_n1090), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[31][11]  (.Q(\ram[31][11] ), 
	.D(FE_PHN837_n1089), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][10]  (.Q(\ram[31][10] ), 
	.D(FE_PHN4152_n1088), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[31][9]  (.Q(\ram[31][9] ), 
	.D(FE_PHN4988_n1087), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][8]  (.Q(\ram[31][8] ), 
	.D(FE_PHN5693_n1086), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][7]  (.Q(\ram[31][7] ), 
	.D(FE_PHN572_n1085), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][6]  (.Q(\ram[31][6] ), 
	.D(FE_PHN1144_n1084), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][5]  (.Q(\ram[31][5] ), 
	.D(FE_PHN2861_n1083), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][4]  (.Q(\ram[31][4] ), 
	.D(FE_PHN3676_n1082), 
	.CK(clk_m__L3_N121));
   QDFFEHD \ram_reg[31][3]  (.Q(\ram[31][3] ), 
	.D(FE_PHN966_n1081), 
	.CK(clk_m__L3_N103));
   QDFFEHD \ram_reg[31][2]  (.Q(\ram[31][2] ), 
	.D(n1080), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[31][1]  (.Q(\ram[31][1] ), 
	.D(FE_PHN5277_n1079), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[31][0]  (.Q(\ram[31][0] ), 
	.D(FE_PHN4962_n1078), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[27][15]  (.Q(\ram[27][15] ), 
	.D(FE_PHN4346_n1029), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[27][14]  (.Q(\ram[27][14] ), 
	.D(FE_PHN5739_n1028), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][13]  (.Q(\ram[27][13] ), 
	.D(FE_PHN3672_n1027), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[27][12]  (.Q(\ram[27][12] ), 
	.D(FE_PHN4313_n1026), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[27][11]  (.Q(\ram[27][11] ), 
	.D(FE_PHN4286_n1025), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][10]  (.Q(\ram[27][10] ), 
	.D(FE_PHN4371_n1024), 
	.CK(clk_m__L3_N125));
   QDFFEHD \ram_reg[27][9]  (.Q(\ram[27][9] ), 
	.D(FE_PHN4621_n1023), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][8]  (.Q(\ram[27][8] ), 
	.D(FE_PHN3431_n1022), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][7]  (.Q(\ram[27][7] ), 
	.D(FE_PHN4606_n1021), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[27][6]  (.Q(\ram[27][6] ), 
	.D(FE_PHN3745_n1020), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][5]  (.Q(\ram[27][5] ), 
	.D(FE_PHN5723_n1019), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[27][4]  (.Q(\ram[27][4] ), 
	.D(FE_PHN3623_n1018), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[27][3]  (.Q(\ram[27][3] ), 
	.D(FE_PHN3454_n1017), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[27][2]  (.Q(\ram[27][2] ), 
	.D(FE_PHN4411_n1016), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[27][1]  (.Q(\ram[27][1] ), 
	.D(FE_PHN5671_n1015), 
	.CK(clk_m__L3_N136));
   QDFFEHD \ram_reg[27][0]  (.Q(\ram[27][0] ), 
	.D(FE_PHN3375_n1014), 
	.CK(clk_m__L3_N120));
   QDFFEHD \ram_reg[23][15]  (.Q(\ram[23][15] ), 
	.D(FE_PHN4454_n965), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][14]  (.Q(\ram[23][14] ), 
	.D(FE_PHN4380_n964), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][13]  (.Q(\ram[23][13] ), 
	.D(FE_PHN1183_n963), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[23][12]  (.Q(\ram[23][12] ), 
	.D(FE_PHN4663_n962), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][11]  (.Q(\ram[23][11] ), 
	.D(FE_PHN4183_n961), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[23][10]  (.Q(\ram[23][10] ), 
	.D(FE_PHN4046_n960), 
	.CK(clk_m__L3_N165));
   QDFFEHD \ram_reg[23][9]  (.Q(\ram[23][9] ), 
	.D(FE_PHN5330_n959), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][8]  (.Q(\ram[23][8] ), 
	.D(FE_PHN4104_n958), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[23][7]  (.Q(\ram[23][7] ), 
	.D(FE_PHN3682_n957), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][6]  (.Q(\ram[23][6] ), 
	.D(FE_PHN2068_n956), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[23][5]  (.Q(\ram[23][5] ), 
	.D(FE_PHN2304_n955), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[23][4]  (.Q(\ram[23][4] ), 
	.D(FE_PHN4309_n954), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][3]  (.Q(\ram[23][3] ), 
	.D(FE_PHN5705_n953), 
	.CK(clk_m__L3_N134));
   QDFFEHD \ram_reg[23][2]  (.Q(\ram[23][2] ), 
	.D(FE_PHN4198_n952), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[23][1]  (.Q(\ram[23][1] ), 
	.D(FE_PHN5041_n951), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[23][0]  (.Q(\ram[23][0] ), 
	.D(FE_PHN6473_n950), 
	.CK(clk_m__L3_N137));
   QDFFEHD \ram_reg[19][15]  (.Q(\ram[19][15] ), 
	.D(FE_PHN4154_n901), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[19][14]  (.Q(\ram[19][14] ), 
	.D(FE_PHN5465_n900), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][13]  (.Q(\ram[19][13] ), 
	.D(FE_PHN4022_n899), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[19][12]  (.Q(\ram[19][12] ), 
	.D(FE_PHN4628_n898), 
	.CK(clk_m__L3_N123));
   QDFFEHD \ram_reg[19][11]  (.Q(\ram[19][11] ), 
	.D(FE_PHN4467_n897), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][10]  (.Q(\ram[19][10] ), 
	.D(FE_PHN4687_n896), 
	.CK(clk_m__L3_N122));
   QDFFEHD \ram_reg[19][9]  (.Q(\ram[19][9] ), 
	.D(FE_PHN4707_n895), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][8]  (.Q(\ram[19][8] ), 
	.D(FE_PHN3522_n894), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[19][7]  (.Q(\ram[19][7] ), 
	.D(FE_PHN4194_n893), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][6]  (.Q(\ram[19][6] ), 
	.D(FE_PHN4699_n892), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[19][5]  (.Q(\ram[19][5] ), 
	.D(FE_PHN4339_n891), 
	.CK(clk_m__L3_N132));
   QDFFEHD \ram_reg[19][4]  (.Q(\ram[19][4] ), 
	.D(FE_PHN4374_n890), 
	.CK(clk_m__L3_N118));
   QDFFEHD \ram_reg[19][3]  (.Q(\ram[19][3] ), 
	.D(FE_PHN4008_n889), 
	.CK(clk_m__L3_N133));
   QDFFEHD \ram_reg[19][2]  (.Q(\ram[19][2] ), 
	.D(FE_PHN4488_n888), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[19][1]  (.Q(\ram[19][1] ), 
	.D(FE_PHN4266_n887), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[19][0]  (.Q(\ram[19][0] ), 
	.D(FE_PHN4679_n886), 
	.CK(clk_m__L3_N119));
   QDFFEHD \ram_reg[15][15]  (.Q(\ram[15][15] ), 
	.D(FE_PHN2895_n837), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][14]  (.Q(\ram[15][14] ), 
	.D(FE_PHN1714_n836), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[15][13]  (.Q(\ram[15][13] ), 
	.D(FE_PHN1572_n835), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][12]  (.Q(\ram[15][12] ), 
	.D(FE_PHN2385_n834), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[15][11]  (.Q(\ram[15][11] ), 
	.D(FE_PHN1165_n833), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[15][10]  (.Q(\ram[15][10] ), 
	.D(FE_PHN3176_n832), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[15][9]  (.Q(\ram[15][9] ), 
	.D(FE_PHN2672_n831), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][8]  (.Q(\ram[15][8] ), 
	.D(FE_PHN2788_n830), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[15][7]  (.Q(\ram[15][7] ), 
	.D(FE_PHN2241_n829), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[15][6]  (.Q(\ram[15][6] ), 
	.D(FE_PHN3034_n828), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[15][5]  (.Q(\ram[15][5] ), 
	.D(FE_PHN1274_n827), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[15][4]  (.Q(\ram[15][4] ), 
	.D(FE_PHN1417_n826), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[15][3]  (.Q(\ram[15][3] ), 
	.D(FE_PHN1545_n825), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[15][2]  (.Q(\ram[15][2] ), 
	.D(FE_PHN1824_n824), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[15][1]  (.Q(\ram[15][1] ), 
	.D(FE_PHN1026_n823), 
	.CK(clk_m__L3_N99));
   QDFFEHD \ram_reg[15][0]  (.Q(\ram[15][0] ), 
	.D(FE_PHN1975_n822), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][15]  (.Q(\ram[11][15] ), 
	.D(FE_PHN2835_n773), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[11][14]  (.Q(\ram[11][14] ), 
	.D(FE_PHN1791_n772), 
	.CK(clk_m__L3_N113));
   QDFFEHD \ram_reg[11][13]  (.Q(\ram[11][13] ), 
	.D(FE_PHN1658_n771), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[11][12]  (.Q(\ram[11][12] ), 
	.D(FE_PHN3149_n770), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][11]  (.Q(\ram[11][11] ), 
	.D(FE_PHN465_n769), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][10]  (.Q(\ram[11][10] ), 
	.D(FE_PHN3209_n768), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[11][9]  (.Q(\ram[11][9] ), 
	.D(FE_PHN1589_n767), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][8]  (.Q(\ram[11][8] ), 
	.D(FE_PHN2592_n766), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[11][7]  (.Q(\ram[11][7] ), 
	.D(FE_PHN1385_n765), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[11][6]  (.Q(\ram[11][6] ), 
	.D(FE_PHN1669_n764), 
	.CK(clk_m__L3_N111));
   QDFFEHD \ram_reg[11][5]  (.Q(\ram[11][5] ), 
	.D(FE_PHN245_n763), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][4]  (.Q(\ram[11][4] ), 
	.D(FE_PHN1996_n762), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][3]  (.Q(\ram[11][3] ), 
	.D(FE_PHN2926_n761), 
	.CK(clk_m__L3_N110));
   QDFFEHD \ram_reg[11][2]  (.Q(\ram[11][2] ), 
	.D(FE_PHN2242_n760), 
	.CK(clk_m__L3_N114));
   QDFFEHD \ram_reg[11][1]  (.Q(\ram[11][1] ), 
	.D(FE_PHN2028_n759), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[11][0]  (.Q(\ram[11][0] ), 
	.D(FE_PHN3137_n758), 
	.CK(clk_m__L3_N116));
   QDFFEHD \ram_reg[7][15]  (.Q(\ram[7][15] ), 
	.D(FE_PHN2035_n709), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][14]  (.Q(\ram[7][14] ), 
	.D(FE_PHN1638_n708), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][13]  (.Q(\ram[7][13] ), 
	.D(FE_PHN1621_n707), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[7][12]  (.Q(\ram[7][12] ), 
	.D(FE_PHN3195_n706), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[7][11]  (.Q(\ram[7][11] ), 
	.D(FE_PHN2266_n705), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][10]  (.Q(\ram[7][10] ), 
	.D(FE_PHN1786_n704), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][9]  (.Q(\ram[7][9] ), 
	.D(FE_PHN2031_n703), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[7][8]  (.Q(\ram[7][8] ), 
	.D(FE_PHN2891_n702), 
	.CK(clk_m__L3_N145));
   QDFFEHD \ram_reg[7][7]  (.Q(\ram[7][7] ), 
	.D(FE_PHN2255_n701), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][6]  (.Q(\ram[7][6] ), 
	.D(FE_PHN2430_n700), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[7][5]  (.Q(\ram[7][5] ), 
	.D(FE_PHN2975_n699), 
	.CK(clk_m__L3_N141));
   QDFFEHD \ram_reg[7][4]  (.Q(\ram[7][4] ), 
	.D(FE_PHN1550_n698), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][3]  (.Q(\ram[7][3] ), 
	.D(FE_PHN1329_n697), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[7][2]  (.Q(\ram[7][2] ), 
	.D(FE_PHN1684_n696), 
	.CK(clk_m__L3_N128));
   QDFFEHD \ram_reg[7][1]  (.Q(\ram[7][1] ), 
	.D(FE_PHN1956_n695), 
	.CK(clk_m__L3_N130));
   QDFFEHD \ram_reg[7][0]  (.Q(\ram[7][0] ), 
	.D(FE_PHN982_n694), 
	.CK(clk_m__L3_N135));
   QDFFEHD \ram_reg[3][15]  (.Q(\ram[3][15] ), 
	.D(FE_PHN2836_n645), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][14]  (.Q(\ram[3][14] ), 
	.D(FE_PHN1727_n644), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][13]  (.Q(\ram[3][13] ), 
	.D(FE_PHN2880_n643), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][12]  (.Q(\ram[3][12] ), 
	.D(FE_PHN2478_n642), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][11]  (.Q(\ram[3][11] ), 
	.D(FE_PHN3084_n641), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[3][10]  (.Q(\ram[3][10] ), 
	.D(FE_PHN753_n640), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[3][9]  (.Q(\ram[3][9] ), 
	.D(FE_PHN2419_n639), 
	.CK(clk_m__L3_N142));
   QDFFEHD \ram_reg[3][8]  (.Q(\ram[3][8] ), 
	.D(FE_PHN2396_n638), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][7]  (.Q(\ram[3][7] ), 
	.D(FE_PHN2117_n637), 
	.CK(clk_m__L3_N112));
   QDFFEHD \ram_reg[3][6]  (.Q(\ram[3][6] ), 
	.D(FE_PHN2105_n636), 
	.CK(clk_m__L3_N140));
   QDFFEHD \ram_reg[3][5]  (.Q(\ram[3][5] ), 
	.D(FE_PHN2383_n635), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[3][4]  (.Q(\ram[3][4] ), 
	.D(FE_PHN2639_n634), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][3]  (.Q(\ram[3][3] ), 
	.D(FE_PHN2871_n633), 
	.CK(clk_m__L3_N109));
   QDFFEHD \ram_reg[3][2]  (.Q(\ram[3][2] ), 
	.D(FE_PHN2284_n632), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][1]  (.Q(\ram[3][1] ), 
	.D(FE_PHN3043_n631), 
	.CK(clk_m__L3_N131));
   QDFFEHD \ram_reg[3][0]  (.Q(\ram[3][0] ), 
	.D(FE_PHN1837_n630), 
	.CK(clk_m__L3_N131));
   AN2EHD U2 (.O(n1), 
	.I2(n545), 
	.I1(n544));
   AN2EHD U3 (.O(n2), 
	.I2(n544), 
	.I1(n548));
   AN2HHD U4 (.O(n3), 
	.I2(n545), 
	.I1(n557));
   AN2HHD U5 (.O(n4), 
	.I2(n548), 
	.I1(n557));
   AN2HHD U6 (.O(n5), 
	.I2(n551), 
	.I1(n557));
   AN2HHD U7 (.O(n7), 
	.I2(n554), 
	.I1(n557));
   AN2HHD U8 (.O(n24), 
	.I2(n545), 
	.I1(n566));
   AN2HHD U9 (.O(n25), 
	.I2(n545), 
	.I1(n575));
   AN2EHD U10 (.O(n26), 
	.I2(n544), 
	.I1(n551));
   AN2EHD U11 (.O(n28), 
	.I2(n544), 
	.I1(n554));
   AN2HHD U12 (.O(n29), 
	.I2(n548), 
	.I1(n566));
   AN2EHD U13 (.O(n31), 
	.I2(n548), 
	.I1(n575));
   AN2HHD U14 (.O(n32), 
	.I2(n551), 
	.I1(n566));
   AN2HHD U15 (.O(n34), 
	.I2(n554), 
	.I1(n566));
   AN2EHD U16 (.O(n35), 
	.I2(n551), 
	.I1(n575));
   AN2HHD U17 (.O(n37), 
	.I2(n554), 
	.I1(n575));
   AN2EHD U18 (.O(n38), 
	.I2(n72), 
	.I1(n208));
   AN2EHD U19 (.O(n40), 
	.I2(n106), 
	.I1(n208));
   AN2EHD U20 (.O(n41), 
	.I2(n140), 
	.I1(n208));
   AN2EHD U21 (.O(n43), 
	.I2(n174), 
	.I1(n208));
   AN2EHD U22 (.O(n44), 
	.I2(n72), 
	.I1(n341));
   AN2EHD U23 (.O(n46), 
	.I2(n72), 
	.I1(n474));
   AN2EHD U24 (.O(n47), 
	.I2(n106), 
	.I1(n341));
   AN2EHD U25 (.O(n49), 
	.I2(n106), 
	.I1(n474));
   AN2EHD U26 (.O(n50), 
	.I2(n140), 
	.I1(n341));
   AN2EHD U27 (.O(n52), 
	.I2(n174), 
	.I1(n341));
   AN2EHD U28 (.O(n53), 
	.I2(n140), 
	.I1(n474));
   AN2EHD U29 (.O(n55), 
	.I2(n174), 
	.I1(n474));
   AN2EHD U30 (.O(n56), 
	.I2(n1), 
	.I1(n38));
   AN2EHD U31 (.O(n58), 
	.I2(n2), 
	.I1(n38));
   AN2EHD U32 (.O(n59), 
	.I2(n26), 
	.I1(n38));
   AN2EHD U33 (.O(n61), 
	.I2(n28), 
	.I1(n38));
   AN2EHD U34 (.O(n62), 
	.I2(n3), 
	.I1(n38));
   AN2EHD U35 (.O(n64), 
	.I2(n4), 
	.I1(n38));
   AN2EHD U36 (.O(n65), 
	.I2(n5), 
	.I1(n38));
   AN2EHD U37 (.O(n67), 
	.I2(n7), 
	.I1(n38));
   AN2EHD U38 (.O(n68), 
	.I2(n24), 
	.I1(n38));
   AN2EHD U39 (.O(n70), 
	.I2(n29), 
	.I1(n38));
   AN2EHD U40 (.O(n73), 
	.I2(n32), 
	.I1(n38));
   AN2EHD U41 (.O(n75), 
	.I2(n34), 
	.I1(n38));
   AN2EHD U42 (.O(n76), 
	.I2(n25), 
	.I1(n38));
   AN2EHD U43 (.O(n78), 
	.I2(n31), 
	.I1(n38));
   AN2EHD U44 (.O(n80), 
	.I2(n35), 
	.I1(n38));
   AN2EHD U45 (.O(n82), 
	.I2(n37), 
	.I1(n38));
   AN2EHD U46 (.O(n84), 
	.I2(n1), 
	.I1(n40));
   AN2EHD U47 (.O(n86), 
	.I2(n2), 
	.I1(n40));
   AN2EHD U48 (.O(n88), 
	.I2(n26), 
	.I1(n40));
   AN2EHD U49 (.O(n90), 
	.I2(n28), 
	.I1(n40));
   AN2EHD U50 (.O(n92), 
	.I2(n3), 
	.I1(n40));
   AN2EHD U51 (.O(n94), 
	.I2(n4), 
	.I1(n40));
   AN2EHD U52 (.O(n96), 
	.I2(n5), 
	.I1(n40));
   AN2EHD U53 (.O(n98), 
	.I2(n7), 
	.I1(n40));
   AN2EHD U54 (.O(n100), 
	.I2(n24), 
	.I1(n40));
   AN2EHD U55 (.O(n102), 
	.I2(n29), 
	.I1(n40));
   AN2EHD U56 (.O(n104), 
	.I2(n32), 
	.I1(n40));
   AN2EHD U57 (.O(n107), 
	.I2(n34), 
	.I1(n40));
   AN2EHD U58 (.O(n109), 
	.I2(n25), 
	.I1(n40));
   AN2EHD U59 (.O(n110), 
	.I2(n31), 
	.I1(n40));
   AN2EHD U60 (.O(n112), 
	.I2(n35), 
	.I1(n40));
   AN2EHD U61 (.O(n114), 
	.I2(n37), 
	.I1(n40));
   AN2EHD U62 (.O(n116), 
	.I2(n1), 
	.I1(n41));
   AN2EHD U63 (.O(n118), 
	.I2(n2), 
	.I1(n41));
   AN2EHD U64 (.O(n120), 
	.I2(n26), 
	.I1(n41));
   AN2EHD U65 (.O(n122), 
	.I2(n28), 
	.I1(n41));
   AN2EHD U66 (.O(n124), 
	.I2(n3), 
	.I1(n41));
   AN2EHD U67 (.O(n126), 
	.I2(n4), 
	.I1(n41));
   AN2EHD U68 (.O(n128), 
	.I2(n5), 
	.I1(n41));
   AN2EHD U69 (.O(n130), 
	.I2(n7), 
	.I1(n41));
   AN2EHD U70 (.O(n132), 
	.I2(n24), 
	.I1(n41));
   AN2EHD U71 (.O(n134), 
	.I2(n29), 
	.I1(n41));
   AN2EHD U72 (.O(n136), 
	.I2(n32), 
	.I1(n41));
   AN2EHD U73 (.O(n138), 
	.I2(n34), 
	.I1(n41));
   AN2EHD U74 (.O(n141), 
	.I2(n25), 
	.I1(n41));
   AN2EHD U75 (.O(n143), 
	.I2(n31), 
	.I1(n41));
   AN2EHD U76 (.O(n144), 
	.I2(n35), 
	.I1(n41));
   AN2EHD U77 (.O(n146), 
	.I2(n37), 
	.I1(n41));
   AN2EHD U78 (.O(n148), 
	.I2(n1), 
	.I1(n43));
   AN2EHD U79 (.O(n150), 
	.I2(n2), 
	.I1(n43));
   AN2EHD U80 (.O(n152), 
	.I2(n26), 
	.I1(n43));
   AN2EHD U81 (.O(n154), 
	.I2(n28), 
	.I1(n43));
   AN2EHD U82 (.O(n156), 
	.I2(n3), 
	.I1(n43));
   AN2EHD U83 (.O(n158), 
	.I2(n4), 
	.I1(n43));
   AN2EHD U84 (.O(n160), 
	.I2(n5), 
	.I1(n43));
   AN2EHD U85 (.O(n162), 
	.I2(n7), 
	.I1(n43));
   AN2EHD U86 (.O(n164), 
	.I2(n24), 
	.I1(n43));
   AN2EHD U87 (.O(n166), 
	.I2(n29), 
	.I1(n43));
   AN2EHD U88 (.O(n168), 
	.I2(n32), 
	.I1(n43));
   AN2EHD U89 (.O(n170), 
	.I2(n34), 
	.I1(n43));
   AN2EHD U90 (.O(n172), 
	.I2(n25), 
	.I1(n43));
   AN2EHD U91 (.O(n175), 
	.I2(n31), 
	.I1(n43));
   AN2EHD U92 (.O(n177), 
	.I2(n35), 
	.I1(n43));
   AN2EHD U93 (.O(n178), 
	.I2(n37), 
	.I1(n43));
   AN2EHD U94 (.O(n180), 
	.I2(n1), 
	.I1(n44));
   AN2EHD U95 (.O(n182), 
	.I2(n2), 
	.I1(n44));
   AN2EHD U96 (.O(n184), 
	.I2(n26), 
	.I1(n44));
   AN2EHD U97 (.O(n186), 
	.I2(n28), 
	.I1(n44));
   AN2EHD U98 (.O(n188), 
	.I2(n3), 
	.I1(n44));
   AN2EHD U99 (.O(n190), 
	.I2(n4), 
	.I1(n44));
   AN2EHD U100 (.O(n192), 
	.I2(n5), 
	.I1(n44));
   AN2EHD U101 (.O(n194), 
	.I2(n7), 
	.I1(n44));
   AN2EHD U102 (.O(n196), 
	.I2(n24), 
	.I1(n44));
   AN2EHD U103 (.O(n198), 
	.I2(n29), 
	.I1(n44));
   AN2EHD U104 (.O(n200), 
	.I2(n32), 
	.I1(n44));
   AN2EHD U105 (.O(n202), 
	.I2(n34), 
	.I1(n44));
   AN2EHD U106 (.O(n204), 
	.I2(n25), 
	.I1(n44));
   AN2EHD U107 (.O(n206), 
	.I2(n31), 
	.I1(n44));
   AN2EHD U108 (.O(n209), 
	.I2(n35), 
	.I1(n44));
   AN2EHD U109 (.O(n211), 
	.I2(n37), 
	.I1(n44));
   AN2EHD U110 (.O(n212), 
	.I2(n1), 
	.I1(n47));
   AN2EHD U111 (.O(n214), 
	.I2(n2), 
	.I1(n47));
   AN2EHD U112 (.O(n216), 
	.I2(n26), 
	.I1(n47));
   AN2EHD U113 (.O(n218), 
	.I2(n28), 
	.I1(n47));
   AN2EHD U114 (.O(n220), 
	.I2(n3), 
	.I1(n47));
   AN2EHD U115 (.O(n222), 
	.I2(n4), 
	.I1(n47));
   AN2EHD U116 (.O(n224), 
	.I2(n5), 
	.I1(n47));
   AN2EHD U117 (.O(n226), 
	.I2(n7), 
	.I1(n47));
   AN2EHD U118 (.O(n228), 
	.I2(n24), 
	.I1(n47));
   AN2EHD U119 (.O(n230), 
	.I2(n29), 
	.I1(n47));
   AN2EHD U120 (.O(n232), 
	.I2(n32), 
	.I1(n47));
   AN2EHD U121 (.O(n234), 
	.I2(n34), 
	.I1(n47));
   AN2EHD U122 (.O(n236), 
	.I2(n25), 
	.I1(n47));
   AN2EHD U123 (.O(n238), 
	.I2(n31), 
	.I1(n47));
   AN2EHD U124 (.O(n240), 
	.I2(n35), 
	.I1(n47));
   AN2EHD U125 (.O(n242), 
	.I2(n37), 
	.I1(n47));
   AN2EHD U126 (.O(n244), 
	.I2(n1), 
	.I1(n50));
   AN2EHD U127 (.O(n245), 
	.I2(n2), 
	.I1(n50));
   AN2EHD U128 (.O(n247), 
	.I2(n26), 
	.I1(n50));
   AN2EHD U129 (.O(n249), 
	.I2(n28), 
	.I1(n50));
   AN2EHD U130 (.O(n251), 
	.I2(n3), 
	.I1(n50));
   AN2EHD U131 (.O(n253), 
	.I2(n4), 
	.I1(n50));
   AN2EHD U132 (.O(n255), 
	.I2(n5), 
	.I1(n50));
   AN2EHD U133 (.O(n257), 
	.I2(n7), 
	.I1(n50));
   AN2EHD U134 (.O(n259), 
	.I2(n24), 
	.I1(n50));
   AN2EHD U135 (.O(n261), 
	.I2(n29), 
	.I1(n50));
   AN2EHD U136 (.O(n263), 
	.I2(n32), 
	.I1(n50));
   AN2EHD U137 (.O(n265), 
	.I2(n34), 
	.I1(n50));
   AN2EHD U138 (.O(n267), 
	.I2(n25), 
	.I1(n50));
   AN2EHD U139 (.O(n269), 
	.I2(n31), 
	.I1(n50));
   AN2EHD U140 (.O(n271), 
	.I2(n35), 
	.I1(n50));
   AN2EHD U141 (.O(n273), 
	.I2(n37), 
	.I1(n50));
   AN2EHD U142 (.O(n275), 
	.I2(n1), 
	.I1(n52));
   AN2EHD U143 (.O(n277), 
	.I2(n2), 
	.I1(n52));
   AN2EHD U144 (.O(n278), 
	.I2(n26), 
	.I1(n52));
   AN2EHD U145 (.O(n280), 
	.I2(n28), 
	.I1(n52));
   AN2EHD U146 (.O(n282), 
	.I2(n3), 
	.I1(n52));
   AN2EHD U147 (.O(n284), 
	.I2(n4), 
	.I1(n52));
   AN2EHD U148 (.O(n286), 
	.I2(n5), 
	.I1(n52));
   AN2EHD U149 (.O(n288), 
	.I2(n7), 
	.I1(n52));
   AN2EHD U150 (.O(n290), 
	.I2(n24), 
	.I1(n52));
   AN2EHD U151 (.O(n292), 
	.I2(n29), 
	.I1(n52));
   AN2EHD U152 (.O(n294), 
	.I2(n32), 
	.I1(n52));
   AN2EHD U153 (.O(n296), 
	.I2(n34), 
	.I1(n52));
   AN2EHD U154 (.O(n298), 
	.I2(n25), 
	.I1(n52));
   AN2EHD U155 (.O(n300), 
	.I2(n31), 
	.I1(n52));
   AN2EHD U156 (.O(n302), 
	.I2(n35), 
	.I1(n52));
   AN2EHD U157 (.O(n304), 
	.I2(n37), 
	.I1(n52));
   AN2EHD U158 (.O(n306), 
	.I2(n1), 
	.I1(n46));
   AN2EHD U159 (.O(n308), 
	.I2(n2), 
	.I1(n46));
   AN2EHD U160 (.O(n310), 
	.I2(n26), 
	.I1(n46));
   AN2EHD U161 (.O(n311), 
	.I2(n28), 
	.I1(n46));
   AN2EHD U162 (.O(n313), 
	.I2(n3), 
	.I1(n46));
   AN2EHD U163 (.O(n315), 
	.I2(n4), 
	.I1(n46));
   AN2EHD U164 (.O(n317), 
	.I2(n5), 
	.I1(n46));
   AN2EHD U165 (.O(n319), 
	.I2(n7), 
	.I1(n46));
   AN2EHD U166 (.O(n321), 
	.I2(n24), 
	.I1(n46));
   AN2EHD U167 (.O(n323), 
	.I2(n29), 
	.I1(n46));
   AN2EHD U168 (.O(n325), 
	.I2(n32), 
	.I1(n46));
   AN2EHD U169 (.O(n327), 
	.I2(n34), 
	.I1(n46));
   AN2EHD U170 (.O(n329), 
	.I2(n25), 
	.I1(n46));
   AN2EHD U171 (.O(n331), 
	.I2(n31), 
	.I1(n46));
   AN2EHD U172 (.O(n333), 
	.I2(n35), 
	.I1(n46));
   AN2EHD U173 (.O(n335), 
	.I2(n37), 
	.I1(n46));
   AN2EHD U174 (.O(n337), 
	.I2(n1), 
	.I1(n49));
   AN2EHD U175 (.O(n339), 
	.I2(n2), 
	.I1(n49));
   AN2EHD U176 (.O(n342), 
	.I2(n26), 
	.I1(n49));
   AN2EHD U177 (.O(n344), 
	.I2(n28), 
	.I1(n49));
   AN2EHD U178 (.O(n345), 
	.I2(n3), 
	.I1(n49));
   AN2EHD U179 (.O(n347), 
	.I2(n4), 
	.I1(n49));
   AN2EHD U180 (.O(n349), 
	.I2(n5), 
	.I1(n49));
   AN2EHD U181 (.O(n351), 
	.I2(n7), 
	.I1(n49));
   AN2EHD U182 (.O(n353), 
	.I2(n24), 
	.I1(n49));
   AN2EHD U183 (.O(n355), 
	.I2(n29), 
	.I1(n49));
   AN2EHD U184 (.O(n357), 
	.I2(n32), 
	.I1(n49));
   AN2EHD U185 (.O(n359), 
	.I2(n34), 
	.I1(n49));
   AN2EHD U186 (.O(n361), 
	.I2(n25), 
	.I1(n49));
   AN2EHD U187 (.O(n363), 
	.I2(n31), 
	.I1(n49));
   AN2EHD U188 (.O(n365), 
	.I2(n35), 
	.I1(n49));
   AN2EHD U189 (.O(n367), 
	.I2(n37), 
	.I1(n49));
   AN2EHD U190 (.O(n369), 
	.I2(n1), 
	.I1(n53));
   AN2EHD U191 (.O(n371), 
	.I2(n2), 
	.I1(n53));
   AN2EHD U192 (.O(n373), 
	.I2(n26), 
	.I1(n53));
   AN2EHD U193 (.O(n375), 
	.I2(n28), 
	.I1(n53));
   AN2EHD U194 (.O(n377), 
	.I2(n3), 
	.I1(n53));
   AN2EHD U195 (.O(n378), 
	.I2(n4), 
	.I1(n53));
   AN2EHD U196 (.O(n380), 
	.I2(n5), 
	.I1(n53));
   AN2EHD U197 (.O(n382), 
	.I2(n7), 
	.I1(n53));
   AN2EHD U198 (.O(n384), 
	.I2(n24), 
	.I1(n53));
   AN2EHD U199 (.O(n386), 
	.I2(n29), 
	.I1(n53));
   AN2EHD U200 (.O(n388), 
	.I2(n32), 
	.I1(n53));
   AN2EHD U201 (.O(n390), 
	.I2(n34), 
	.I1(n53));
   AN2EHD U202 (.O(n392), 
	.I2(n25), 
	.I1(n53));
   AN2EHD U203 (.O(n394), 
	.I2(n31), 
	.I1(n53));
   AN2EHD U204 (.O(n396), 
	.I2(n35), 
	.I1(n53));
   AN2EHD U205 (.O(n398), 
	.I2(n37), 
	.I1(n53));
   AN2EHD U206 (.O(n400), 
	.I2(n1), 
	.I1(n55));
   AN2EHD U207 (.O(n402), 
	.I2(n2), 
	.I1(n55));
   AN2EHD U208 (.O(n404), 
	.I2(n26), 
	.I1(n55));
   AN2EHD U209 (.O(n406), 
	.I2(n28), 
	.I1(n55));
   AN2EHD U210 (.O(n408), 
	.I2(n3), 
	.I1(n55));
   AN2EHD U211 (.O(n410), 
	.I2(n4), 
	.I1(n55));
   AN2EHD U212 (.O(n411), 
	.I2(n5), 
	.I1(n55));
   AN2EHD U213 (.O(n413), 
	.I2(n7), 
	.I1(n55));
   AN2EHD U214 (.O(n415), 
	.I2(n24), 
	.I1(n55));
   AN2EHD U215 (.O(n417), 
	.I2(n29), 
	.I1(n55));
   AN2EHD U216 (.O(n419), 
	.I2(n32), 
	.I1(n55));
   AN2EHD U217 (.O(n421), 
	.I2(n34), 
	.I1(n55));
   AN2EHD U218 (.O(n423), 
	.I2(n25), 
	.I1(n55));
   AN2EHD U219 (.O(n425), 
	.I2(n31), 
	.I1(n55));
   AN2EHD U220 (.O(n427), 
	.I2(n35), 
	.I1(n55));
   AN2EHD U221 (.O(n429), 
	.I2(n37), 
	.I1(n55));
   AN2EHD U222 (.O(n431), 
	.I2(n72), 
	.I1(n71));
   AN2EHD U223 (.O(n433), 
	.I2(n431), 
	.I1(n1));
   AN2EHD U224 (.O(n435), 
	.I2(n71), 
	.I1(n106));
   AN2EHD U225 (.O(n437), 
	.I2(n71), 
	.I1(n140));
   AN2EHD U226 (.O(n439), 
	.I2(n71), 
	.I1(n174));
   AN2EHD U227 (.O(n441), 
	.I2(n431), 
	.I1(n2));
   AN2EHD U228 (.O(n443), 
	.I2(n431), 
	.I1(n26));
   AN2EHD U229 (.O(n444), 
	.I2(n431), 
	.I1(n28));
   AN2EHD U230 (.O(n446), 
	.I2(n431), 
	.I1(n3));
   AN2EHD U231 (.O(n448), 
	.I2(n431), 
	.I1(n4));
   AN2EHD U232 (.O(n450), 
	.I2(n431), 
	.I1(n5));
   AN2EHD U233 (.O(n452), 
	.I2(n431), 
	.I1(n7));
   AN2EHD U234 (.O(n454), 
	.I2(n431), 
	.I1(n24));
   AN2EHD U235 (.O(n456), 
	.I2(n431), 
	.I1(n29));
   AN2EHD U236 (.O(n458), 
	.I2(n431), 
	.I1(n32));
   AN2EHD U237 (.O(n460), 
	.I2(n431), 
	.I1(n34));
   AN2EHD U238 (.O(n462), 
	.I2(n431), 
	.I1(n25));
   AN2EHD U239 (.O(n464), 
	.I2(n431), 
	.I1(n31));
   AN2EHD U240 (.O(n466), 
	.I2(n431), 
	.I1(n35));
   AN2EHD U241 (.O(n468), 
	.I2(n431), 
	.I1(n37));
   AN2EHD U242 (.O(n470), 
	.I2(n1), 
	.I1(n435));
   AN2EHD U243 (.O(n472), 
	.I2(n2), 
	.I1(n435));
   AN2EHD U244 (.O(n475), 
	.I2(n26), 
	.I1(n435));
   AN2EHD U245 (.O(n477), 
	.I2(n28), 
	.I1(n435));
   AN2EHD U246 (.O(n478), 
	.I2(n3), 
	.I1(n435));
   AN2EHD U247 (.O(n480), 
	.I2(n4), 
	.I1(n435));
   AN2EHD U248 (.O(n482), 
	.I2(n5), 
	.I1(n435));
   AN2EHD U249 (.O(n484), 
	.I2(n7), 
	.I1(n435));
   AN2EHD U250 (.O(n486), 
	.I2(n24), 
	.I1(n435));
   AN2EHD U251 (.O(n488), 
	.I2(n29), 
	.I1(n435));
   AN2EHD U252 (.O(n490), 
	.I2(n32), 
	.I1(n435));
   AN2EHD U253 (.O(n492), 
	.I2(n34), 
	.I1(n435));
   AN2EHD U254 (.O(n494), 
	.I2(n25), 
	.I1(n435));
   AN2EHD U255 (.O(n496), 
	.I2(n31), 
	.I1(n435));
   AN2EHD U256 (.O(n498), 
	.I2(n35), 
	.I1(n435));
   AN2EHD U257 (.O(n500), 
	.I2(n37), 
	.I1(n435));
   AN2EHD U258 (.O(n502), 
	.I2(n1), 
	.I1(n437));
   AN2EHD U259 (.O(n504), 
	.I2(n2), 
	.I1(n437));
   AN2EHD U260 (.O(n506), 
	.I2(n26), 
	.I1(n437));
   AN2EHD U261 (.O(n508), 
	.I2(n28), 
	.I1(n437));
   AN2EHD U262 (.O(n510), 
	.I2(n3), 
	.I1(n437));
   AN2EHD U263 (.O(n511), 
	.I2(n4), 
	.I1(n437));
   AN2EHD U264 (.O(n513), 
	.I2(n5), 
	.I1(n437));
   AN2EHD U265 (.O(n515), 
	.I2(n7), 
	.I1(n437));
   AN2EHD U266 (.O(n517), 
	.I2(n24), 
	.I1(n437));
   AN2EHD U267 (.O(n519), 
	.I2(n29), 
	.I1(n437));
   AN2EHD U268 (.O(n521), 
	.I2(n32), 
	.I1(n437));
   AN2EHD U269 (.O(n523), 
	.I2(n34), 
	.I1(n437));
   AN2EHD U270 (.O(n525), 
	.I2(n25), 
	.I1(n437));
   AN2EHD U271 (.O(n527), 
	.I2(n31), 
	.I1(n437));
   AN2EHD U272 (.O(n529), 
	.I2(n35), 
	.I1(n437));
   AN2EHD U273 (.O(n531), 
	.I2(n37), 
	.I1(n437));
   AN2EHD U274 (.O(n533), 
	.I2(n1), 
	.I1(n439));
   AN2EHD U275 (.O(n535), 
	.I2(n2), 
	.I1(n439));
   AN2EHD U276 (.O(n537), 
	.I2(n26), 
	.I1(n439));
   AN2EHD U277 (.O(n539), 
	.I2(n28), 
	.I1(n439));
   AN2EHD U278 (.O(n541), 
	.I2(n3), 
	.I1(n439));
   AN2EHD U279 (.O(n543), 
	.I2(n4), 
	.I1(n439));
   AN2EHD U280 (.O(n546), 
	.I2(n5), 
	.I1(n439));
   AN2EHD U281 (.O(n549), 
	.I2(n7), 
	.I1(n439));
   AN2EHD U282 (.O(n552), 
	.I2(n24), 
	.I1(n439));
   AN2EHD U283 (.O(n555), 
	.I2(n29), 
	.I1(n439));
   AN2EHD U284 (.O(n558), 
	.I2(n32), 
	.I1(n439));
   AN2EHD U285 (.O(n560), 
	.I2(n34), 
	.I1(n439));
   AN2EHD U286 (.O(n562), 
	.I2(n25), 
	.I1(n439));
   AN2EHD U287 (.O(n564), 
	.I2(n31), 
	.I1(n439));
   AN2EHD U288 (.O(n567), 
	.I2(n35), 
	.I1(n439));
   AN2EHD U289 (.O(n569), 
	.I2(n37), 
	.I1(n439));
   ND2DHD U751 (.O(n27), 
	.I2(mem_write_en), 
	.I1(n441));
   ND2DHD U753 (.O(n30), 
	.I2(mem_write_en), 
	.I1(n443));
   ND2DHD U755 (.O(n33), 
	.I2(mem_write_en), 
	.I1(n444));
   ND2DHD U757 (.O(n36), 
	.I2(mem_write_en), 
	.I1(n446));
   ND2DHD U759 (.O(n39), 
	.I2(mem_write_en), 
	.I1(n448));
   ND2DHD U761 (.O(n42), 
	.I2(mem_write_en), 
	.I1(n450));
   ND2DHD U763 (.O(n45), 
	.I2(mem_write_en), 
	.I1(n452));
   ND2DHD U765 (.O(n48), 
	.I2(mem_write_en), 
	.I1(n454));
   ND2DHD U767 (.O(n51), 
	.I2(mem_write_en), 
	.I1(n456));
   ND2DHD U769 (.O(n54), 
	.I2(mem_write_en), 
	.I1(n458));
   ND2DHD U771 (.O(n57), 
	.I2(mem_write_en), 
	.I1(n460));
   ND2DHD U773 (.O(n60), 
	.I2(mem_write_en), 
	.I1(n462));
   ND2DHD U775 (.O(n63), 
	.I2(mem_write_en), 
	.I1(n464));
   ND2DHD U777 (.O(n66), 
	.I2(mem_write_en), 
	.I1(n466));
   ND2DHD U779 (.O(n69), 
	.I2(mem_write_en), 
	.I1(n468));
   ND2DHD U781 (.O(n74), 
	.I2(mem_write_en), 
	.I1(n470));
   ND2DHD U783 (.O(n77), 
	.I2(mem_write_en), 
	.I1(n472));
   ND2DHD U785 (.O(n79), 
	.I2(mem_write_en), 
	.I1(n475));
   ND2DHD U787 (.O(n81), 
	.I2(mem_write_en), 
	.I1(n477));
   ND2DHD U789 (.O(n83), 
	.I2(FE_OFN94_mem_write), 
	.I1(n478));
   ND2DHD U791 (.O(n85), 
	.I2(FE_OFN94_mem_write), 
	.I1(n480));
   ND2DHD U793 (.O(n87), 
	.I2(FE_OFN94_mem_write), 
	.I1(n482));
   ND2DHD U795 (.O(n89), 
	.I2(FE_OFN94_mem_write), 
	.I1(n484));
   ND2DHD U797 (.O(n91), 
	.I2(mem_write_en), 
	.I1(n486));
   ND2DHD U799 (.O(n93), 
	.I2(mem_write_en), 
	.I1(n488));
   ND2DHD U801 (.O(n95), 
	.I2(mem_write_en), 
	.I1(n490));
   ND2DHD U803 (.O(n97), 
	.I2(mem_write_en), 
	.I1(n492));
   ND2DHD U805 (.O(n99), 
	.I2(mem_write_en), 
	.I1(n494));
   ND2DHD U807 (.O(n101), 
	.I2(mem_write_en), 
	.I1(n496));
   ND2DHD U809 (.O(n103), 
	.I2(mem_write_en), 
	.I1(n498));
   ND2DHD U811 (.O(n105), 
	.I2(mem_write_en), 
	.I1(n500));
   ND2DHD U813 (.O(n108), 
	.I2(mem_write_en), 
	.I1(n502));
   ND2DHD U815 (.O(n111), 
	.I2(mem_write_en), 
	.I1(n504));
   ND2DHD U817 (.O(n113), 
	.I2(mem_write_en), 
	.I1(n506));
   ND2DHD U819 (.O(n115), 
	.I2(mem_write_en), 
	.I1(n508));
   ND2DHD U821 (.O(n117), 
	.I2(mem_write_en), 
	.I1(n510));
   ND2DHD U823 (.O(n119), 
	.I2(mem_write_en), 
	.I1(n511));
   ND2DHD U825 (.O(n121), 
	.I2(mem_write_en), 
	.I1(n513));
   ND2DHD U827 (.O(n123), 
	.I2(mem_write_en), 
	.I1(n515));
   ND2DHD U829 (.O(n125), 
	.I2(FE_OFN94_mem_write), 
	.I1(n517));
   ND2DHD U831 (.O(n127), 
	.I2(FE_OFN94_mem_write), 
	.I1(n519));
   ND2DHD U833 (.O(n129), 
	.I2(FE_OFN94_mem_write), 
	.I1(n521));
   ND2DHD U835 (.O(n131), 
	.I2(FE_OFN94_mem_write), 
	.I1(n523));
   ND2DHD U837 (.O(n133), 
	.I2(FE_OFN94_mem_write), 
	.I1(n525));
   ND2DHD U839 (.O(n135), 
	.I2(FE_OFN94_mem_write), 
	.I1(n527));
   ND2DHD U841 (.O(n137), 
	.I2(mem_write_en), 
	.I1(n529));
   ND2DHD U843 (.O(n139), 
	.I2(FE_OFN94_mem_write), 
	.I1(n531));
   ND2DHD U845 (.O(n142), 
	.I2(FE_OFN94_mem_write), 
	.I1(n533));
   ND2DHD U847 (.O(n145), 
	.I2(FE_OFN94_mem_write), 
	.I1(n535));
   ND2DHD U849 (.O(n147), 
	.I2(FE_OFN94_mem_write), 
	.I1(n537));
   ND2DHD U851 (.O(n149), 
	.I2(FE_OFN94_mem_write), 
	.I1(n539));
   ND2DHD U853 (.O(n151), 
	.I2(FE_OFN94_mem_write), 
	.I1(n541));
   ND2DHD U855 (.O(n153), 
	.I2(FE_OFN94_mem_write), 
	.I1(n543));
   ND2DHD U857 (.O(n155), 
	.I2(FE_OFN94_mem_write), 
	.I1(n546));
   ND2DHD U859 (.O(n157), 
	.I2(FE_OFN94_mem_write), 
	.I1(n549));
   ND2DHD U861 (.O(n159), 
	.I2(FE_OFN94_mem_write), 
	.I1(n552));
   ND2DHD U863 (.O(n161), 
	.I2(FE_OFN94_mem_write), 
	.I1(n555));
   ND2DHD U865 (.O(n163), 
	.I2(FE_OFN94_mem_write), 
	.I1(n558));
   ND2DHD U867 (.O(n165), 
	.I2(FE_OFN94_mem_write), 
	.I1(n560));
   ND2DHD U869 (.O(n167), 
	.I2(FE_OFN94_mem_write), 
	.I1(n562));
   ND2DHD U871 (.O(n169), 
	.I2(FE_OFN94_mem_write), 
	.I1(n564));
   ND2DHD U873 (.O(n171), 
	.I2(FE_OFN94_mem_write), 
	.I1(n567));
   ND2DHD U875 (.O(n173), 
	.I2(FE_OFN94_mem_write), 
	.I1(n569));
   ND2DHD U877 (.O(n176), 
	.I2(FE_OFN94_mem_write), 
	.I1(n56));
   ND2DHD U879 (.O(n179), 
	.I2(FE_OFN94_mem_write), 
	.I1(n58));
   ND2DHD U881 (.O(n181), 
	.I2(FE_OFN94_mem_write), 
	.I1(n59));
   ND2DHD U883 (.O(n183), 
	.I2(FE_OFN94_mem_write), 
	.I1(n61));
   ND2DHD U885 (.O(n185), 
	.I2(FE_OFN94_mem_write), 
	.I1(n62));
   ND2DHD U887 (.O(n187), 
	.I2(FE_OFN94_mem_write), 
	.I1(n64));
   ND2DHD U889 (.O(n189), 
	.I2(FE_OFN94_mem_write), 
	.I1(n65));
   ND2DHD U891 (.O(n191), 
	.I2(FE_OFN94_mem_write), 
	.I1(n67));
   ND2DHD U893 (.O(n193), 
	.I2(FE_OFN92_mem_write), 
	.I1(n68));
   ND2DHD U895 (.O(n195), 
	.I2(FE_OFN92_mem_write), 
	.I1(n70));
   ND2DHD U897 (.O(n197), 
	.I2(FE_OFN92_mem_write), 
	.I1(n73));
   ND2DHD U899 (.O(n199), 
	.I2(FE_OFN92_mem_write), 
	.I1(n75));
   ND2DHD U901 (.O(n201), 
	.I2(FE_OFN92_mem_write), 
	.I1(n76));
   ND2DHD U903 (.O(n203), 
	.I2(FE_OFN92_mem_write), 
	.I1(n78));
   ND2DHD U905 (.O(n205), 
	.I2(FE_OFN92_mem_write), 
	.I1(n80));
   ND2DHD U907 (.O(n207), 
	.I2(FE_OFN92_mem_write), 
	.I1(n82));
   ND2DHD U909 (.O(n210), 
	.I2(FE_OFN94_mem_write), 
	.I1(n84));
   ND2DHD U911 (.O(n213), 
	.I2(FE_OFN94_mem_write), 
	.I1(n86));
   ND2DHD U913 (.O(n215), 
	.I2(FE_OFN94_mem_write), 
	.I1(n88));
   ND2DHD U915 (.O(n217), 
	.I2(FE_OFN94_mem_write), 
	.I1(n90));
   ND2DHD U917 (.O(n219), 
	.I2(FE_OFN94_mem_write), 
	.I1(n92));
   ND2DHD U919 (.O(n221), 
	.I2(FE_OFN94_mem_write), 
	.I1(n94));
   ND2DHD U921 (.O(n223), 
	.I2(FE_OFN94_mem_write), 
	.I1(n96));
   ND2DHD U923 (.O(n225), 
	.I2(FE_OFN94_mem_write), 
	.I1(n98));
   ND2DHD U925 (.O(n227), 
	.I2(FE_OFN94_mem_write), 
	.I1(n100));
   ND2DHD U927 (.O(n229), 
	.I2(FE_OFN94_mem_write), 
	.I1(n102));
   ND2DHD U929 (.O(n231), 
	.I2(FE_OFN94_mem_write), 
	.I1(n104));
   ND2DHD U931 (.O(n233), 
	.I2(FE_OFN94_mem_write), 
	.I1(n107));
   ND2DHD U933 (.O(n235), 
	.I2(FE_OFN94_mem_write), 
	.I1(n109));
   ND2DHD U935 (.O(n237), 
	.I2(FE_OFN94_mem_write), 
	.I1(n110));
   ND2DHD U937 (.O(n239), 
	.I2(FE_OFN94_mem_write), 
	.I1(n112));
   ND2DHD U939 (.O(n241), 
	.I2(FE_OFN94_mem_write), 
	.I1(n114));
   ND2DHD U941 (.O(n243), 
	.I2(FE_OFN92_mem_write), 
	.I1(n116));
   ND2DHD U943 (.O(n246), 
	.I2(FE_OFN92_mem_write), 
	.I1(n118));
   ND2DHD U945 (.O(n248), 
	.I2(FE_OFN92_mem_write), 
	.I1(n120));
   ND2DHD U947 (.O(n250), 
	.I2(FE_OFN92_mem_write), 
	.I1(n122));
   ND2DHD U949 (.O(n252), 
	.I2(FE_OFN94_mem_write), 
	.I1(n124));
   ND2DHD U951 (.O(n254), 
	.I2(FE_OFN94_mem_write), 
	.I1(n126));
   ND2DHD U953 (.O(n256), 
	.I2(FE_OFN94_mem_write), 
	.I1(n128));
   ND2DHD U955 (.O(n258), 
	.I2(FE_OFN94_mem_write), 
	.I1(n130));
   ND2DHD U957 (.O(n260), 
	.I2(FE_OFN94_mem_write), 
	.I1(n132));
   ND2DHD U959 (.O(n262), 
	.I2(FE_OFN94_mem_write), 
	.I1(n134));
   ND2DHD U961 (.O(n264), 
	.I2(FE_OFN94_mem_write), 
	.I1(n136));
   ND2DHD U963 (.O(n266), 
	.I2(FE_OFN94_mem_write), 
	.I1(n138));
   ND2DHD U965 (.O(n268), 
	.I2(FE_OFN94_mem_write), 
	.I1(n141));
   ND2DHD U967 (.O(n270), 
	.I2(FE_OFN94_mem_write), 
	.I1(n143));
   ND2DHD U969 (.O(n272), 
	.I2(FE_OFN94_mem_write), 
	.I1(n144));
   ND2DHD U971 (.O(n274), 
	.I2(FE_OFN94_mem_write), 
	.I1(n146));
   ND2DHD U973 (.O(n276), 
	.I2(FE_OFN92_mem_write), 
	.I1(n148));
   ND2DHD U975 (.O(n279), 
	.I2(FE_OFN92_mem_write), 
	.I1(n150));
   ND2DHD U977 (.O(n281), 
	.I2(FE_OFN92_mem_write), 
	.I1(n152));
   ND2DHD U979 (.O(n283), 
	.I2(FE_OFN92_mem_write), 
	.I1(n154));
   ND2DHD U981 (.O(n285), 
	.I2(FE_OFN94_mem_write), 
	.I1(n156));
   ND2DHD U983 (.O(n287), 
	.I2(FE_OFN94_mem_write), 
	.I1(n158));
   ND2DHD U985 (.O(n289), 
	.I2(FE_OFN94_mem_write), 
	.I1(n160));
   ND2DHD U987 (.O(n291), 
	.I2(FE_OFN94_mem_write), 
	.I1(n162));
   ND2DHD U989 (.O(n293), 
	.I2(FE_OFN94_mem_write), 
	.I1(n164));
   ND2DHD U991 (.O(n295), 
	.I2(FE_OFN94_mem_write), 
	.I1(n166));
   ND2DHD U993 (.O(n297), 
	.I2(FE_OFN94_mem_write), 
	.I1(n168));
   ND2DHD U995 (.O(n299), 
	.I2(FE_OFN94_mem_write), 
	.I1(n170));
   ND2DHD U997 (.O(n301), 
	.I2(FE_OFN94_mem_write), 
	.I1(n172));
   ND2DHD U999 (.O(n303), 
	.I2(FE_OFN94_mem_write), 
	.I1(n175));
   ND2DHD U1001 (.O(n305), 
	.I2(FE_OFN94_mem_write), 
	.I1(n177));
   ND2DHD U1003 (.O(n307), 
	.I2(FE_OFN94_mem_write), 
	.I1(n178));
   ND2DHD U1005 (.O(n309), 
	.I2(FE_OFN93_mem_write), 
	.I1(n180));
   ND2DHD U1007 (.O(n312), 
	.I2(FE_OFN93_mem_write), 
	.I1(n182));
   ND2DHD U1009 (.O(n314), 
	.I2(FE_OFN93_mem_write), 
	.I1(n184));
   ND2DHD U1011 (.O(n316), 
	.I2(FE_OFN93_mem_write), 
	.I1(n186));
   ND2DHD U1013 (.O(n318), 
	.I2(FE_OFN93_mem_write), 
	.I1(n188));
   ND2DHD U1015 (.O(n320), 
	.I2(FE_OFN93_mem_write), 
	.I1(n190));
   ND2DHD U1017 (.O(n322), 
	.I2(FE_OFN93_mem_write), 
	.I1(n192));
   ND2DHD U1019 (.O(n324), 
	.I2(FE_OFN93_mem_write), 
	.I1(n194));
   ND2DHD U1021 (.O(n326), 
	.I2(FE_OFN93_mem_write), 
	.I1(n196));
   ND2DHD U1023 (.O(n328), 
	.I2(FE_OFN93_mem_write), 
	.I1(n198));
   ND2DHD U1025 (.O(n334), 
	.I2(FE_OFN93_mem_write), 
	.I1(n204));
   ND2DHD U1027 (.O(n338), 
	.I2(FE_OFN93_mem_write), 
	.I1(n209));
   ND2DHD U1029 (.O(n340), 
	.I2(FE_OFN93_mem_write), 
	.I1(n211));
   ND2DHD U1031 (.O(n343), 
	.I2(FE_OFN93_mem_write), 
	.I1(n212));
   ND2DHD U1033 (.O(n346), 
	.I2(FE_OFN93_mem_write), 
	.I1(n214));
   ND2DHD U1035 (.O(n348), 
	.I2(FE_OFN93_mem_write), 
	.I1(n216));
   ND2DHD U1037 (.O(n350), 
	.I2(FE_OFN93_mem_write), 
	.I1(n218));
   ND2DHD U1039 (.O(n352), 
	.I2(mem_write_en), 
	.I1(n220));
   ND2DHD U1041 (.O(n354), 
	.I2(mem_write_en), 
	.I1(n222));
   ND2DHD U1043 (.O(n356), 
	.I2(mem_write_en), 
	.I1(n224));
   ND2DHD U1045 (.O(n358), 
	.I2(mem_write_en), 
	.I1(n226));
   ND2DHD U1047 (.O(n360), 
	.I2(mem_write_en), 
	.I1(n228));
   ND2DHD U1049 (.O(n362), 
	.I2(mem_write_en), 
	.I1(n230));
   ND2DHD U1051 (.O(n364), 
	.I2(mem_write_en), 
	.I1(n232));
   ND2DHD U1053 (.O(n366), 
	.I2(mem_write_en), 
	.I1(n234));
   ND2DHD U1055 (.O(n368), 
	.I2(FE_OFN93_mem_write), 
	.I1(n236));
   ND2DHD U1057 (.O(n370), 
	.I2(FE_OFN93_mem_write), 
	.I1(n238));
   ND2DHD U1059 (.O(n372), 
	.I2(FE_OFN93_mem_write), 
	.I1(n240));
   ND2DHD U1061 (.O(n374), 
	.I2(FE_OFN93_mem_write), 
	.I1(n242));
   ND2DHD U1063 (.O(n376), 
	.I2(FE_OFN93_mem_write), 
	.I1(n244));
   ND2DHD U1065 (.O(n379), 
	.I2(FE_OFN93_mem_write), 
	.I1(n245));
   ND2DHD U1067 (.O(n381), 
	.I2(FE_OFN93_mem_write), 
	.I1(n247));
   ND2DHD U1069 (.O(n383), 
	.I2(FE_OFN93_mem_write), 
	.I1(n249));
   ND2DHD U1071 (.O(n385), 
	.I2(FE_OFN93_mem_write), 
	.I1(n251));
   ND2DHD U1073 (.O(n387), 
	.I2(FE_OFN93_mem_write), 
	.I1(n253));
   ND2DHD U1075 (.O(n389), 
	.I2(FE_OFN93_mem_write), 
	.I1(n255));
   ND2DHD U1077 (.O(n391), 
	.I2(FE_OFN93_mem_write), 
	.I1(n257));
   ND2DHD U1079 (.O(n393), 
	.I2(FE_OFN93_mem_write), 
	.I1(n259));
   ND2DHD U1081 (.O(n395), 
	.I2(FE_OFN93_mem_write), 
	.I1(n261));
   ND2DHD U1083 (.O(n397), 
	.I2(FE_OFN93_mem_write), 
	.I1(n263));
   ND2DHD U1085 (.O(n399), 
	.I2(FE_OFN93_mem_write), 
	.I1(n265));
   ND2DHD U1087 (.O(n401), 
	.I2(FE_OFN93_mem_write), 
	.I1(n267));
   ND2DHD U1089 (.O(n403), 
	.I2(FE_OFN93_mem_write), 
	.I1(n269));
   ND2DHD U1091 (.O(n405), 
	.I2(FE_OFN93_mem_write), 
	.I1(n271));
   ND2DHD U1093 (.O(n407), 
	.I2(FE_OFN93_mem_write), 
	.I1(n273));
   ND2DHD U1095 (.O(n409), 
	.I2(mem_write_en), 
	.I1(n275));
   ND2DHD U1097 (.O(n412), 
	.I2(mem_write_en), 
	.I1(n277));
   ND2DHD U1099 (.O(n414), 
	.I2(mem_write_en), 
	.I1(n278));
   ND2DHD U1101 (.O(n416), 
	.I2(mem_write_en), 
	.I1(n280));
   ND2DHD U1103 (.O(n418), 
	.I2(FE_OFN93_mem_write), 
	.I1(n282));
   ND2DHD U1105 (.O(n420), 
	.I2(FE_OFN93_mem_write), 
	.I1(n284));
   ND2DHD U1107 (.O(n422), 
	.I2(FE_OFN93_mem_write), 
	.I1(n286));
   ND2DHD U1109 (.O(n424), 
	.I2(FE_OFN93_mem_write), 
	.I1(n288));
   ND2DHD U1111 (.O(n426), 
	.I2(FE_OFN93_mem_write), 
	.I1(n290));
   ND2DHD U1113 (.O(n428), 
	.I2(FE_OFN93_mem_write), 
	.I1(n292));
   ND2DHD U1115 (.O(n430), 
	.I2(FE_OFN93_mem_write), 
	.I1(n294));
   ND2DHD U1117 (.O(n432), 
	.I2(FE_OFN93_mem_write), 
	.I1(n296));
   ND2DHD U1119 (.O(n434), 
	.I2(FE_OFN93_mem_write), 
	.I1(n298));
   ND2DHD U1121 (.O(n436), 
	.I2(FE_OFN93_mem_write), 
	.I1(n300));
   ND2DHD U1123 (.O(n438), 
	.I2(FE_OFN93_mem_write), 
	.I1(n302));
   ND2DHD U1125 (.O(n440), 
	.I2(FE_OFN93_mem_write), 
	.I1(n304));
   ND2DHD U1127 (.O(n442), 
	.I2(FE_OFN92_mem_write), 
	.I1(n306));
   ND2DHD U1129 (.O(n445), 
	.I2(FE_OFN92_mem_write), 
	.I1(n308));
   ND2DHD U1131 (.O(n447), 
	.I2(FE_OFN92_mem_write), 
	.I1(n310));
   ND2DHD U1133 (.O(n449), 
	.I2(FE_OFN92_mem_write), 
	.I1(n311));
   ND2DHD U1135 (.O(n451), 
	.I2(FE_OFN92_mem_write), 
	.I1(n313));
   ND2DHD U1137 (.O(n453), 
	.I2(FE_OFN92_mem_write), 
	.I1(n315));
   ND2DHD U1139 (.O(n455), 
	.I2(FE_OFN92_mem_write), 
	.I1(n317));
   ND2DHD U1141 (.O(n457), 
	.I2(FE_OFN92_mem_write), 
	.I1(n319));
   ND2DHD U1143 (.O(n459), 
	.I2(FE_OFN92_mem_write), 
	.I1(n321));
   ND2DHD U1145 (.O(n461), 
	.I2(FE_OFN92_mem_write), 
	.I1(n323));
   ND2DHD U1147 (.O(n463), 
	.I2(FE_OFN92_mem_write), 
	.I1(n325));
   ND2DHD U1149 (.O(n465), 
	.I2(FE_OFN92_mem_write), 
	.I1(n327));
   ND2DHD U1151 (.O(n467), 
	.I2(FE_OFN92_mem_write), 
	.I1(n329));
   ND2DHD U1153 (.O(n469), 
	.I2(FE_OFN92_mem_write), 
	.I1(n331));
   ND2DHD U1155 (.O(n471), 
	.I2(FE_OFN92_mem_write), 
	.I1(n333));
   ND2DHD U1157 (.O(n473), 
	.I2(FE_OFN92_mem_write), 
	.I1(n335));
   ND2DHD U1159 (.O(n476), 
	.I2(FE_OFN92_mem_write), 
	.I1(n337));
   ND2DHD U1161 (.O(n479), 
	.I2(FE_OFN92_mem_write), 
	.I1(n339));
   ND2DHD U1163 (.O(n481), 
	.I2(FE_OFN92_mem_write), 
	.I1(n342));
   ND2DHD U1165 (.O(n483), 
	.I2(FE_OFN92_mem_write), 
	.I1(n344));
   ND2DHD U1167 (.O(n485), 
	.I2(FE_OFN92_mem_write), 
	.I1(n345));
   ND2DHD U1169 (.O(n487), 
	.I2(FE_OFN92_mem_write), 
	.I1(n347));
   ND2DHD U1171 (.O(n489), 
	.I2(FE_OFN92_mem_write), 
	.I1(n349));
   ND2DHD U1173 (.O(n491), 
	.I2(FE_OFN92_mem_write), 
	.I1(n351));
   ND2DHD U1175 (.O(n493), 
	.I2(FE_OFN92_mem_write), 
	.I1(n353));
   ND2DHD U1177 (.O(n495), 
	.I2(FE_OFN92_mem_write), 
	.I1(n355));
   ND2DHD U1179 (.O(n497), 
	.I2(FE_OFN92_mem_write), 
	.I1(n357));
   ND2DHD U1181 (.O(n499), 
	.I2(FE_OFN92_mem_write), 
	.I1(n359));
   ND2DHD U1183 (.O(n501), 
	.I2(FE_OFN92_mem_write), 
	.I1(n361));
   ND2DHD U1185 (.O(n503), 
	.I2(FE_OFN92_mem_write), 
	.I1(n363));
   ND2DHD U1187 (.O(n505), 
	.I2(FE_OFN92_mem_write), 
	.I1(n365));
   ND2DHD U1189 (.O(n507), 
	.I2(FE_OFN92_mem_write), 
	.I1(n367));
   ND2DHD U1191 (.O(n509), 
	.I2(FE_OFN92_mem_write), 
	.I1(n369));
   ND2DHD U1193 (.O(n512), 
	.I2(FE_OFN92_mem_write), 
	.I1(n371));
   ND2DHD U1195 (.O(n514), 
	.I2(FE_OFN92_mem_write), 
	.I1(n373));
   ND2DHD U1197 (.O(n516), 
	.I2(FE_OFN92_mem_write), 
	.I1(n375));
   ND2DHD U1199 (.O(n518), 
	.I2(FE_OFN92_mem_write), 
	.I1(n377));
   ND2DHD U1201 (.O(n520), 
	.I2(FE_OFN92_mem_write), 
	.I1(n378));
   ND2DHD U1203 (.O(n522), 
	.I2(FE_OFN92_mem_write), 
	.I1(n380));
   ND2DHD U1205 (.O(n524), 
	.I2(FE_OFN92_mem_write), 
	.I1(n382));
   ND2DHD U1207 (.O(n526), 
	.I2(FE_OFN93_mem_write), 
	.I1(n384));
   ND2DHD U1209 (.O(n528), 
	.I2(FE_OFN93_mem_write), 
	.I1(n386));
   ND2DHD U1211 (.O(n530), 
	.I2(FE_OFN93_mem_write), 
	.I1(n388));
   ND2DHD U1213 (.O(n532), 
	.I2(FE_OFN93_mem_write), 
	.I1(n390));
   ND2DHD U1215 (.O(n534), 
	.I2(FE_OFN93_mem_write), 
	.I1(n392));
   ND2DHD U1217 (.O(n536), 
	.I2(FE_OFN93_mem_write), 
	.I1(n394));
   ND2DHD U1219 (.O(n538), 
	.I2(FE_OFN93_mem_write), 
	.I1(n396));
   ND2DHD U1221 (.O(n540), 
	.I2(FE_OFN93_mem_write), 
	.I1(n398));
   ND2DHD U1223 (.O(n542), 
	.I2(FE_OFN93_mem_write), 
	.I1(n400));
   ND2DHD U1225 (.O(n547), 
	.I2(FE_OFN93_mem_write), 
	.I1(n402));
   ND2DHD U1227 (.O(n550), 
	.I2(FE_OFN93_mem_write), 
	.I1(n404));
   ND2DHD U1229 (.O(n553), 
	.I2(FE_OFN93_mem_write), 
	.I1(n406));
   ND2DHD U1231 (.O(n556), 
	.I2(FE_OFN93_mem_write), 
	.I1(n408));
   ND2DHD U1233 (.O(n559), 
	.I2(FE_OFN93_mem_write), 
	.I1(n410));
   ND2DHD U1235 (.O(n561), 
	.I2(FE_OFN93_mem_write), 
	.I1(n411));
   ND2DHD U1237 (.O(n563), 
	.I2(FE_OFN93_mem_write), 
	.I1(n413));
   ND2DHD U1239 (.O(n565), 
	.I2(FE_OFN92_mem_write), 
	.I1(n415));
   ND2DHD U1241 (.O(n568), 
	.I2(FE_OFN92_mem_write), 
	.I1(n417));
   ND2DHD U1243 (.O(n570), 
	.I2(FE_OFN92_mem_write), 
	.I1(n419));
   ND2DHD U1245 (.O(n572), 
	.I2(FE_OFN92_mem_write), 
	.I1(n421));
   ND2DHD U1247 (.O(n574), 
	.I2(FE_OFN92_mem_write), 
	.I1(n423));
   ND2DHD U1249 (.O(n577), 
	.I2(FE_OFN92_mem_write), 
	.I1(n425));
   ND2DHD U1251 (.O(n579), 
	.I2(FE_OFN92_mem_write), 
	.I1(n427));
   ND2DHD U1253 (.O(n581), 
	.I2(FE_OFN92_mem_write), 
	.I1(n429));
   ND2DHD U1255 (.O(n330), 
	.I2(FE_OFN93_mem_write), 
	.I1(n200));
   ND2DHD U1257 (.O(n332), 
	.I2(FE_OFN93_mem_write), 
	.I1(n202));
   ND2DHD U1259 (.O(n336), 
	.I2(FE_OFN93_mem_write), 
	.I1(n206));
   ND2DHD U1261 (.O(n8), 
	.I2(n433), 
	.I1(mem_write_en));
   BUFEHD U1267 (.O(n6459), 
	.I(N20));
   BUFHHD U1271 (.O(n6136), 
	.I(N22));
   BUFHHD U1272 (.O(n6038), 
	.I(N24));
   AN2EHD U1671 (.O(n140), 
	.I2(n7443), 
	.I1(n7444));
   AN2EHD U1672 (.O(n551), 
	.I2(n7439), 
	.I1(n7440));
   AN2EHD U1673 (.O(n174), 
	.I2(N24), 
	.I1(n7444));
   AN2EHD U1674 (.O(n554), 
	.I2(N20), 
	.I1(n7440));
   NR2CHD U1675 (.O(n72), 
	.I2(n7444), 
	.I1(N24));
   NR2CHD U1676 (.O(n106), 
	.I2(n7444), 
	.I1(n7443));
   NR2BHD U1677 (.O(n544), 
	.I2(n7442), 
	.I1(N22));
   AN2EHD U1678 (.O(n566), 
	.I2(n7441), 
	.I1(n7442));
   AN2EHD U1679 (.O(n575), 
	.I2(N22), 
	.I1(n7442));
   NR2BHD U1680 (.O(n557), 
	.I2(n7442), 
	.I1(n7441));
   NR2CHD U1681 (.O(n545), 
	.I2(n7440), 
	.I1(N20));
   NR2CHD U1682 (.O(n548), 
	.I2(n7440), 
	.I1(n7439));
   INVDHD U1879 (.O(n7443), 
	.I(N24));
   INVDHD U1880 (.O(n7441), 
	.I(N22));
   INVDHD U1881 (.O(n7439), 
	.I(N20));
   BUFIHD U1882 (.O(n7440), 
	.I(N21));
   BUFHHD U1883 (.O(n7442), 
	.I(N23));
   BUFIHD U1884 (.O(n7444), 
	.I(N25));
   NR2CHD U1951 (.O(n71), 
	.I2(N27), 
	.I1(N26));
   NR2CHD U1952 (.O(n208), 
	.I2(N27), 
	.I1(n7445));
   INVDHD U1953 (.O(n7445), 
	.I(N26));
   AN2EHD U1954 (.O(n341), 
	.I2(n7445), 
	.I1(N27));
   AN2EHD U1955 (.O(n474), 
	.I2(N26), 
	.I1(N27));
   BUFEHD U1956 (.O(n6470), 
	.I(N27));
   BUFEHD U1957 (.O(n6469), 
	.I(N26));
   AN2EHD U1990 (.O(mem_read_data[9]), 
	.I2(N4132), 
	.I1(n6471));
   AN2EHD U1991 (.O(mem_read_data[8]), 
	.I2(n6471), 
	.I1(N4133));
   AN2EHD U1992 (.O(mem_read_data[1]), 
	.I2(n6471), 
	.I1(N4140));
   AN2EHD U1993 (.O(mem_read_data[2]), 
	.I2(n6471), 
	.I1(N4139));
   AN2EHD U1994 (.O(mem_read_data[3]), 
	.I2(n6471), 
	.I1(N4138));
   AN2EHD U1995 (.O(mem_read_data[4]), 
	.I2(n6471), 
	.I1(N4137));
   AN2EHD U1996 (.O(mem_read_data[5]), 
	.I2(n6471), 
	.I1(N4136));
   AN2EHD U1997 (.O(mem_read_data[6]), 
	.I2(n6471), 
	.I1(N4135));
   AN2EHD U1998 (.O(mem_read_data[7]), 
	.I2(n6471), 
	.I1(N4134));
   AN2EHD U1999 (.O(mem_read_data[10]), 
	.I2(n6471), 
	.I1(N4131));
   AN2EHD U2000 (.O(mem_read_data[11]), 
	.I2(n6471), 
	.I1(N4130));
   AN2EHD U2001 (.O(mem_read_data[12]), 
	.I2(n6471), 
	.I1(N4129));
   AN2EHD U2002 (.O(mem_read_data[13]), 
	.I2(n6471), 
	.I1(N4128));
   AN2EHD U2003 (.O(mem_read_data[14]), 
	.I2(n6471), 
	.I1(N4127));
   AN2EHD U2004 (.O(mem_read_data[15]), 
	.I2(n6471), 
	.I1(N4126));
   AN2HHD U2005 (.O(n6), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[0]));
   AN2HHD U2006 (.O(n9), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[1]));
   AN2HHD U2007 (.O(n10), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[2]));
   AN2EHD U2008 (.O(n11), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[3]));
   AN2EHD U2009 (.O(n12), 
	.I2(FE_OFN92_mem_write), 
	.I1(mem_write_data[4]));
   AN2EHD U2010 (.O(n13), 
	.I2(mem_write_en), 
	.I1(mem_write_data[5]));
   AN2HHD U2011 (.O(n14), 
	.I2(mem_write_en), 
	.I1(mem_write_data[6]));
   AN2EHD U2012 (.O(n15), 
	.I2(mem_write_en), 
	.I1(mem_write_data[7]));
   AN2EHD U2013 (.O(n16), 
	.I2(mem_write_en), 
	.I1(mem_write_data[8]));
   AN2HHD U2014 (.O(n17), 
	.I2(mem_write_en), 
	.I1(mem_write_data[9]));
   AN2HHD U2015 (.O(n18), 
	.I2(mem_write_en), 
	.I1(mem_write_data[10]));
   AN2HHD U2016 (.O(n19), 
	.I2(mem_write_en), 
	.I1(mem_write_data[11]));
   AN2EHD U2017 (.O(n20), 
	.I2(mem_write_en), 
	.I1(mem_write_data[12]));
   AN2HHD U2018 (.O(n21), 
	.I2(mem_write_en), 
	.I1(mem_write_data[13]));
   AN2HHD U2019 (.O(n22), 
	.I2(mem_write_en), 
	.I1(mem_write_data[14]));
   AN2HHD U2020 (.O(n23), 
	.I2(mem_write_en), 
	.I1(mem_write_data[15]));
   BUFEHD U2021 (.O(n6471), 
	.I(mem_read));
   AN2EHD U2022 (.O(mem_read_data[0]), 
	.I2(n6471), 
	.I1(N4141));
   AO22CHD U2023 (.O(n598), 
	.B2(n27), 
	.B1(\ram[1][0] ), 
	.A2(n6), 
	.A1(n441));
   AO22CHD U2024 (.O(n599), 
	.B2(n27), 
	.B1(\ram[1][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n441));
   AO22CHD U2025 (.O(n600), 
	.B2(n27), 
	.B1(\ram[1][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n441));
   AO22CHD U2026 (.O(n601), 
	.B2(n27), 
	.B1(\ram[1][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n441));
   AO22CHD U2027 (.O(n602), 
	.B2(n27), 
	.B1(\ram[1][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n441));
   AO22CHD U2028 (.O(n603), 
	.B2(n27), 
	.B1(\ram[1][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n441));
   AO22CHD U2029 (.O(n604), 
	.B2(n27), 
	.B1(\ram[1][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n441));
   AO22CHD U2030 (.O(n605), 
	.B2(n27), 
	.B1(\ram[1][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n441));
   AO22CHD U2031 (.O(n606), 
	.B2(n27), 
	.B1(\ram[1][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n441));
   AO22CHD U2032 (.O(n607), 
	.B2(n27), 
	.B1(\ram[1][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n441));
   AO22CHD U2033 (.O(n608), 
	.B2(n27), 
	.B1(\ram[1][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n441));
   AO22CHD U2034 (.O(n609), 
	.B2(n27), 
	.B1(\ram[1][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n441));
   AO22CHD U2035 (.O(n610), 
	.B2(n27), 
	.B1(\ram[1][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n441));
   AO22CHD U2036 (.O(n611), 
	.B2(n27), 
	.B1(\ram[1][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n441));
   AO22CHD U2037 (.O(n612), 
	.B2(n27), 
	.B1(\ram[1][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n441));
   AO22CHD U2038 (.O(n613), 
	.B2(n27), 
	.B1(\ram[1][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n441));
   AO22CHD U2039 (.O(n614), 
	.B2(n30), 
	.B1(\ram[2][0] ), 
	.A2(n6), 
	.A1(n443));
   AO22CHD U2040 (.O(n615), 
	.B2(n30), 
	.B1(\ram[2][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n443));
   AO22CHD U2041 (.O(n616), 
	.B2(n30), 
	.B1(\ram[2][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n443));
   AO22CHD U2042 (.O(n617), 
	.B2(n30), 
	.B1(\ram[2][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n443));
   AO22CHD U2043 (.O(n618), 
	.B2(n30), 
	.B1(\ram[2][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n443));
   AO22CHD U2044 (.O(n619), 
	.B2(n30), 
	.B1(\ram[2][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n443));
   AO22CHD U2045 (.O(n620), 
	.B2(n30), 
	.B1(\ram[2][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n443));
   AO22CHD U2046 (.O(n621), 
	.B2(n30), 
	.B1(\ram[2][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n443));
   AO22CHD U2047 (.O(n622), 
	.B2(n30), 
	.B1(\ram[2][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n443));
   AO22CHD U2048 (.O(n623), 
	.B2(n30), 
	.B1(\ram[2][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n443));
   AO22CHD U2049 (.O(n624), 
	.B2(n30), 
	.B1(\ram[2][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n443));
   AO22CHD U2050 (.O(n625), 
	.B2(n30), 
	.B1(\ram[2][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n443));
   AO22CHD U2051 (.O(n626), 
	.B2(n30), 
	.B1(\ram[2][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n443));
   AO22CHD U2052 (.O(n627), 
	.B2(n30), 
	.B1(\ram[2][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n443));
   AO22CHD U2053 (.O(n628), 
	.B2(n30), 
	.B1(\ram[2][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n443));
   AO22CHD U2054 (.O(n629), 
	.B2(n30), 
	.B1(\ram[2][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n443));
   AO22CHD U2055 (.O(n630), 
	.B2(n33), 
	.B1(\ram[3][0] ), 
	.A2(n6), 
	.A1(n444));
   AO22CHD U2056 (.O(n631), 
	.B2(n33), 
	.B1(\ram[3][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n444));
   AO22CHD U2057 (.O(n632), 
	.B2(n33), 
	.B1(\ram[3][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n444));
   AO22CHD U2058 (.O(n633), 
	.B2(n33), 
	.B1(\ram[3][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n444));
   AO22CHD U2059 (.O(n634), 
	.B2(n33), 
	.B1(\ram[3][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n444));
   AO22CHD U2060 (.O(n635), 
	.B2(n33), 
	.B1(\ram[3][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n444));
   AO22CHD U2061 (.O(n636), 
	.B2(n33), 
	.B1(\ram[3][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n444));
   AO22CHD U2062 (.O(n637), 
	.B2(n33), 
	.B1(\ram[3][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n444));
   AO22CHD U2063 (.O(n638), 
	.B2(n33), 
	.B1(\ram[3][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n444));
   AO22CHD U2064 (.O(n639), 
	.B2(n33), 
	.B1(\ram[3][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n444));
   AO22CHD U2065 (.O(n640), 
	.B2(n33), 
	.B1(\ram[3][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n444));
   AO22CHD U2066 (.O(n641), 
	.B2(n33), 
	.B1(\ram[3][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n444));
   AO22CHD U2067 (.O(n642), 
	.B2(n33), 
	.B1(\ram[3][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n444));
   AO22CHD U2068 (.O(n643), 
	.B2(n33), 
	.B1(\ram[3][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n444));
   AO22CHD U2069 (.O(n644), 
	.B2(n33), 
	.B1(\ram[3][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n444));
   AO22CHD U2070 (.O(n645), 
	.B2(n33), 
	.B1(\ram[3][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n444));
   AO22CHD U2071 (.O(n646), 
	.B2(n36), 
	.B1(\ram[4][0] ), 
	.A2(n6), 
	.A1(n446));
   AO22CHD U2072 (.O(n647), 
	.B2(n36), 
	.B1(\ram[4][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n446));
   AO22CHD U2073 (.O(n648), 
	.B2(n36), 
	.B1(\ram[4][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n446));
   AO22CHD U2074 (.O(n649), 
	.B2(n36), 
	.B1(\ram[4][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n446));
   AO22CHD U2075 (.O(n650), 
	.B2(n36), 
	.B1(\ram[4][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n446));
   AO22CHD U2076 (.O(n651), 
	.B2(n36), 
	.B1(\ram[4][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n446));
   AO22CHD U2077 (.O(n652), 
	.B2(n36), 
	.B1(\ram[4][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n446));
   AO22CHD U2078 (.O(n653), 
	.B2(n36), 
	.B1(\ram[4][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n446));
   AO22CHD U2079 (.O(n654), 
	.B2(n36), 
	.B1(\ram[4][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n446));
   AO22CHD U2080 (.O(n655), 
	.B2(n36), 
	.B1(\ram[4][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n446));
   AO22CHD U2081 (.O(n656), 
	.B2(n36), 
	.B1(\ram[4][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n446));
   AO22CHD U2082 (.O(n657), 
	.B2(n36), 
	.B1(\ram[4][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n446));
   AO22CHD U2083 (.O(n658), 
	.B2(n36), 
	.B1(\ram[4][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n446));
   AO22CHD U2084 (.O(n659), 
	.B2(n36), 
	.B1(\ram[4][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n446));
   AO22CHD U2085 (.O(n660), 
	.B2(n36), 
	.B1(\ram[4][14] ), 
	.A2(n22), 
	.A1(n446));
   AO22CHD U2086 (.O(n661), 
	.B2(n36), 
	.B1(\ram[4][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n446));
   AO22CHD U2087 (.O(n662), 
	.B2(n39), 
	.B1(\ram[5][0] ), 
	.A2(n6), 
	.A1(n448));
   AO22CHD U2088 (.O(n663), 
	.B2(n39), 
	.B1(\ram[5][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n448));
   AO22CHD U2089 (.O(n664), 
	.B2(n39), 
	.B1(\ram[5][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n448));
   AO22CHD U2090 (.O(n665), 
	.B2(n39), 
	.B1(\ram[5][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n448));
   AO22CHD U2091 (.O(n666), 
	.B2(n39), 
	.B1(\ram[5][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n448));
   AO22CHD U2092 (.O(n667), 
	.B2(n39), 
	.B1(\ram[5][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n448));
   AO22CHD U2093 (.O(n668), 
	.B2(n39), 
	.B1(\ram[5][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n448));
   AO22CHD U2094 (.O(n669), 
	.B2(n39), 
	.B1(\ram[5][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n448));
   AO22CHD U2095 (.O(n670), 
	.B2(n39), 
	.B1(\ram[5][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n448));
   AO22CHD U2096 (.O(n671), 
	.B2(n39), 
	.B1(\ram[5][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n448));
   AO22CHD U2097 (.O(n672), 
	.B2(n39), 
	.B1(\ram[5][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n448));
   AO22CHD U2098 (.O(n673), 
	.B2(n39), 
	.B1(\ram[5][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n448));
   AO22CHD U2099 (.O(n674), 
	.B2(n39), 
	.B1(\ram[5][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n448));
   AO22CHD U2100 (.O(n675), 
	.B2(n39), 
	.B1(\ram[5][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n448));
   AO22CHD U2101 (.O(n676), 
	.B2(n39), 
	.B1(\ram[5][14] ), 
	.A2(n22), 
	.A1(n448));
   AO22CHD U2102 (.O(n677), 
	.B2(n39), 
	.B1(\ram[5][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n448));
   AO22CHD U2103 (.O(n678), 
	.B2(n42), 
	.B1(\ram[6][0] ), 
	.A2(n6), 
	.A1(n450));
   AO22CHD U2104 (.O(n679), 
	.B2(n42), 
	.B1(\ram[6][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n450));
   AO22CHD U2105 (.O(n680), 
	.B2(n42), 
	.B1(\ram[6][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n450));
   AO22CHD U2106 (.O(n681), 
	.B2(n42), 
	.B1(\ram[6][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n450));
   AO22CHD U2107 (.O(n682), 
	.B2(n42), 
	.B1(\ram[6][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n450));
   AO22CHD U2108 (.O(n683), 
	.B2(n42), 
	.B1(\ram[6][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n450));
   AO22CHD U2109 (.O(n684), 
	.B2(n42), 
	.B1(\ram[6][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n450));
   AO22CHD U2110 (.O(n685), 
	.B2(n42), 
	.B1(\ram[6][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n450));
   AO22CHD U2111 (.O(n686), 
	.B2(n42), 
	.B1(\ram[6][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n450));
   AO22CHD U2112 (.O(n687), 
	.B2(n42), 
	.B1(\ram[6][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n450));
   AO22CHD U2113 (.O(n688), 
	.B2(n42), 
	.B1(\ram[6][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n450));
   AO22CHD U2114 (.O(n689), 
	.B2(n42), 
	.B1(\ram[6][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n450));
   AO22CHD U2115 (.O(n690), 
	.B2(n42), 
	.B1(\ram[6][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n450));
   AO22CHD U2116 (.O(n691), 
	.B2(n42), 
	.B1(\ram[6][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n450));
   AO22CHD U2117 (.O(n692), 
	.B2(n42), 
	.B1(\ram[6][14] ), 
	.A2(n22), 
	.A1(n450));
   AO22CHD U2118 (.O(n693), 
	.B2(n42), 
	.B1(\ram[6][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n450));
   AO22CHD U2119 (.O(n694), 
	.B2(n45), 
	.B1(\ram[7][0] ), 
	.A2(n6), 
	.A1(n452));
   AO22CHD U2120 (.O(n695), 
	.B2(n45), 
	.B1(\ram[7][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n452));
   AO22CHD U2121 (.O(n696), 
	.B2(n45), 
	.B1(\ram[7][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n452));
   AO22CHD U2122 (.O(n697), 
	.B2(n45), 
	.B1(\ram[7][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n452));
   AO22CHD U2123 (.O(n698), 
	.B2(n45), 
	.B1(\ram[7][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n452));
   AO22CHD U2124 (.O(n699), 
	.B2(n45), 
	.B1(\ram[7][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n452));
   AO22CHD U2125 (.O(n700), 
	.B2(n45), 
	.B1(\ram[7][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n452));
   AO22CHD U2126 (.O(n701), 
	.B2(n45), 
	.B1(\ram[7][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n452));
   AO22CHD U2127 (.O(n702), 
	.B2(n45), 
	.B1(\ram[7][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n452));
   AO22CHD U2128 (.O(n703), 
	.B2(n45), 
	.B1(\ram[7][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n452));
   AO22CHD U2129 (.O(n704), 
	.B2(n45), 
	.B1(\ram[7][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n452));
   AO22CHD U2130 (.O(n705), 
	.B2(n45), 
	.B1(\ram[7][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n452));
   AO22CHD U2131 (.O(n706), 
	.B2(n45), 
	.B1(\ram[7][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n452));
   AO22CHD U2132 (.O(n707), 
	.B2(n45), 
	.B1(\ram[7][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n452));
   AO22CHD U2133 (.O(n708), 
	.B2(n45), 
	.B1(\ram[7][14] ), 
	.A2(n22), 
	.A1(n452));
   AO22CHD U2134 (.O(n709), 
	.B2(n45), 
	.B1(\ram[7][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n452));
   AO22CHD U2135 (.O(n710), 
	.B2(n48), 
	.B1(\ram[8][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n454));
   AO22CHD U2136 (.O(n711), 
	.B2(n48), 
	.B1(\ram[8][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n454));
   AO22CHD U2137 (.O(n712), 
	.B2(n48), 
	.B1(\ram[8][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n454));
   AO22CHD U2138 (.O(n713), 
	.B2(n48), 
	.B1(\ram[8][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n454));
   AO22CHD U2139 (.O(n714), 
	.B2(n48), 
	.B1(\ram[8][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n454));
   AO22CHD U2140 (.O(n715), 
	.B2(n48), 
	.B1(\ram[8][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n454));
   AO22CHD U2141 (.O(n716), 
	.B2(n48), 
	.B1(\ram[8][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n454));
   AO22CHD U2142 (.O(n717), 
	.B2(n48), 
	.B1(\ram[8][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n454));
   AO22CHD U2143 (.O(n718), 
	.B2(n48), 
	.B1(\ram[8][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n454));
   AO22CHD U2144 (.O(n719), 
	.B2(n48), 
	.B1(\ram[8][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n454));
   AO22CHD U2145 (.O(n720), 
	.B2(n48), 
	.B1(\ram[8][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n454));
   AO22CHD U2146 (.O(n721), 
	.B2(n48), 
	.B1(\ram[8][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n454));
   AO22CHD U2147 (.O(n722), 
	.B2(n48), 
	.B1(\ram[8][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n454));
   AO22CHD U2148 (.O(n723), 
	.B2(n48), 
	.B1(\ram[8][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n454));
   AO22CHD U2149 (.O(n724), 
	.B2(n48), 
	.B1(\ram[8][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n454));
   AO22CHD U2150 (.O(n725), 
	.B2(n48), 
	.B1(\ram[8][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n454));
   AO22CHD U2151 (.O(n726), 
	.B2(n51), 
	.B1(\ram[9][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n456));
   AO22CHD U2152 (.O(n727), 
	.B2(n51), 
	.B1(FE_PHN2364_ram_9__1_), 
	.A2(FE_OFN46_n9), 
	.A1(n456));
   AO22CHD U2153 (.O(n728), 
	.B2(n51), 
	.B1(\ram[9][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n456));
   AO22CHD U2154 (.O(n729), 
	.B2(n51), 
	.B1(\ram[9][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n456));
   AO22CHD U2155 (.O(n730), 
	.B2(n51), 
	.B1(\ram[9][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n456));
   AO22CHD U2156 (.O(n731), 
	.B2(n51), 
	.B1(\ram[9][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n456));
   AO22CHD U2157 (.O(n732), 
	.B2(n51), 
	.B1(\ram[9][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n456));
   AO22CHD U2158 (.O(n733), 
	.B2(n51), 
	.B1(\ram[9][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n456));
   AO22CHD U2159 (.O(n734), 
	.B2(n51), 
	.B1(\ram[9][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n456));
   AO22CHD U2160 (.O(n735), 
	.B2(n51), 
	.B1(\ram[9][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n456));
   AO22CHD U2161 (.O(n736), 
	.B2(n51), 
	.B1(\ram[9][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n456));
   AO22CHD U2162 (.O(n737), 
	.B2(n51), 
	.B1(\ram[9][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n456));
   AO22CHD U2163 (.O(n738), 
	.B2(n51), 
	.B1(\ram[9][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n456));
   AO22CHD U2164 (.O(n739), 
	.B2(n51), 
	.B1(\ram[9][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n456));
   AO22CHD U2165 (.O(n740), 
	.B2(n51), 
	.B1(\ram[9][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n456));
   AO22CHD U2166 (.O(n741), 
	.B2(n51), 
	.B1(\ram[9][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n456));
   AO22CHD U2167 (.O(n742), 
	.B2(n54), 
	.B1(\ram[10][0] ), 
	.A2(n6), 
	.A1(n458));
   AO22CHD U2168 (.O(n743), 
	.B2(n54), 
	.B1(\ram[10][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n458));
   AO22CHD U2169 (.O(n744), 
	.B2(n54), 
	.B1(\ram[10][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n458));
   AO22CHD U2170 (.O(n745), 
	.B2(n54), 
	.B1(\ram[10][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n458));
   AO22CHD U2171 (.O(n746), 
	.B2(n54), 
	.B1(\ram[10][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n458));
   AO22CHD U2172 (.O(n747), 
	.B2(n54), 
	.B1(\ram[10][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n458));
   AO22CHD U2173 (.O(n748), 
	.B2(n54), 
	.B1(\ram[10][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n458));
   AO22CHD U2174 (.O(n749), 
	.B2(n54), 
	.B1(\ram[10][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n458));
   AO22CHD U2175 (.O(n750), 
	.B2(n54), 
	.B1(\ram[10][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n458));
   AO22CHD U2176 (.O(n751), 
	.B2(n54), 
	.B1(\ram[10][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n458));
   AO22CHD U2177 (.O(n752), 
	.B2(n54), 
	.B1(\ram[10][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n458));
   AO22CHD U2178 (.O(n753), 
	.B2(n54), 
	.B1(\ram[10][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n458));
   AO22CHD U2179 (.O(n754), 
	.B2(n54), 
	.B1(\ram[10][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n458));
   AO22CHD U2180 (.O(n755), 
	.B2(n54), 
	.B1(\ram[10][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n458));
   AO22CHD U2181 (.O(n756), 
	.B2(n54), 
	.B1(\ram[10][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n458));
   AO22CHD U2182 (.O(n757), 
	.B2(n54), 
	.B1(\ram[10][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n458));
   AO22CHD U2183 (.O(n758), 
	.B2(n57), 
	.B1(\ram[11][0] ), 
	.A2(n6), 
	.A1(n460));
   AO22CHD U2184 (.O(n759), 
	.B2(n57), 
	.B1(\ram[11][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n460));
   AO22CHD U2185 (.O(n760), 
	.B2(n57), 
	.B1(\ram[11][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n460));
   AO22CHD U2186 (.O(n761), 
	.B2(n57), 
	.B1(\ram[11][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n460));
   AO22CHD U2187 (.O(n762), 
	.B2(n57), 
	.B1(\ram[11][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n460));
   AO22CHD U2188 (.O(n763), 
	.B2(n57), 
	.B1(\ram[11][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n460));
   AO22CHD U2189 (.O(n764), 
	.B2(n57), 
	.B1(\ram[11][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n460));
   AO22CHD U2190 (.O(n765), 
	.B2(n57), 
	.B1(\ram[11][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n460));
   AO22CHD U2191 (.O(n766), 
	.B2(n57), 
	.B1(\ram[11][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n460));
   AO22CHD U2192 (.O(n767), 
	.B2(n57), 
	.B1(\ram[11][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n460));
   AO22CHD U2193 (.O(n768), 
	.B2(n57), 
	.B1(\ram[11][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n460));
   AO22CHD U2194 (.O(n769), 
	.B2(n57), 
	.B1(\ram[11][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n460));
   AO22CHD U2195 (.O(n770), 
	.B2(n57), 
	.B1(\ram[11][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n460));
   AO22CHD U2196 (.O(n771), 
	.B2(n57), 
	.B1(\ram[11][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n460));
   AO22CHD U2197 (.O(n772), 
	.B2(n57), 
	.B1(\ram[11][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n460));
   AO22CHD U2198 (.O(n773), 
	.B2(n57), 
	.B1(\ram[11][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n460));
   AO22CHD U2199 (.O(n774), 
	.B2(n60), 
	.B1(\ram[12][0] ), 
	.A2(n6), 
	.A1(n462));
   AO22CHD U2200 (.O(n775), 
	.B2(n60), 
	.B1(\ram[12][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n462));
   AO22CHD U2201 (.O(n776), 
	.B2(n60), 
	.B1(\ram[12][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n462));
   AO22CHD U2202 (.O(n777), 
	.B2(n60), 
	.B1(\ram[12][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n462));
   AO22CHD U2203 (.O(n778), 
	.B2(n60), 
	.B1(\ram[12][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n462));
   AO22CHD U2204 (.O(n779), 
	.B2(n60), 
	.B1(\ram[12][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n462));
   AO22CHD U2205 (.O(n780), 
	.B2(n60), 
	.B1(\ram[12][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n462));
   AO22CHD U2206 (.O(n781), 
	.B2(n60), 
	.B1(\ram[12][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n462));
   AO22CHD U2207 (.O(n782), 
	.B2(n60), 
	.B1(\ram[12][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n462));
   AO22CHD U2208 (.O(n783), 
	.B2(n60), 
	.B1(\ram[12][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n462));
   AO22CHD U2209 (.O(n784), 
	.B2(n60), 
	.B1(\ram[12][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n462));
   AO22CHD U2210 (.O(n785), 
	.B2(n60), 
	.B1(\ram[12][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n462));
   AO22CHD U2211 (.O(n786), 
	.B2(n60), 
	.B1(\ram[12][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n462));
   AO22CHD U2212 (.O(n787), 
	.B2(n60), 
	.B1(\ram[12][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n462));
   AO22CHD U2213 (.O(n788), 
	.B2(n60), 
	.B1(\ram[12][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n462));
   AO22CHD U2214 (.O(n789), 
	.B2(n60), 
	.B1(\ram[12][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n462));
   AO22CHD U2215 (.O(n790), 
	.B2(n63), 
	.B1(\ram[13][0] ), 
	.A2(n6), 
	.A1(n464));
   AO22CHD U2216 (.O(n791), 
	.B2(n63), 
	.B1(\ram[13][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n464));
   AO22CHD U2217 (.O(n792), 
	.B2(n63), 
	.B1(\ram[13][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n464));
   AO22CHD U2218 (.O(n793), 
	.B2(n63), 
	.B1(\ram[13][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n464));
   AO22CHD U2219 (.O(n794), 
	.B2(n63), 
	.B1(\ram[13][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n464));
   AO22CHD U2220 (.O(n795), 
	.B2(n63), 
	.B1(\ram[13][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n464));
   AO22CHD U2221 (.O(n796), 
	.B2(n63), 
	.B1(\ram[13][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n464));
   AO22CHD U2222 (.O(n797), 
	.B2(n63), 
	.B1(\ram[13][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n464));
   AO22CHD U2223 (.O(n798), 
	.B2(n63), 
	.B1(\ram[13][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n464));
   AO22CHD U2224 (.O(n799), 
	.B2(n63), 
	.B1(\ram[13][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n464));
   AO22CHD U2225 (.O(n800), 
	.B2(n63), 
	.B1(\ram[13][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n464));
   AO22CHD U2226 (.O(n801), 
	.B2(n63), 
	.B1(\ram[13][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n464));
   AO22CHD U2227 (.O(n802), 
	.B2(n63), 
	.B1(\ram[13][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n464));
   AO22CHD U2228 (.O(n803), 
	.B2(n63), 
	.B1(\ram[13][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n464));
   AO22CHD U2229 (.O(n804), 
	.B2(n63), 
	.B1(\ram[13][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n464));
   AO22CHD U2230 (.O(n805), 
	.B2(n63), 
	.B1(\ram[13][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n464));
   AO22CHD U2231 (.O(n806), 
	.B2(n66), 
	.B1(\ram[14][0] ), 
	.A2(n6), 
	.A1(n466));
   AO22CHD U2232 (.O(n807), 
	.B2(n66), 
	.B1(\ram[14][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n466));
   AO22CHD U2233 (.O(n808), 
	.B2(n66), 
	.B1(\ram[14][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n466));
   AO22CHD U2234 (.O(n809), 
	.B2(n66), 
	.B1(\ram[14][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n466));
   AO22CHD U2235 (.O(n810), 
	.B2(n66), 
	.B1(\ram[14][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n466));
   AO22CHD U2236 (.O(n811), 
	.B2(n66), 
	.B1(\ram[14][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n466));
   AO22CHD U2237 (.O(n812), 
	.B2(n66), 
	.B1(\ram[14][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n466));
   AO22CHD U2238 (.O(n813), 
	.B2(n66), 
	.B1(\ram[14][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n466));
   AO22CHD U2239 (.O(n814), 
	.B2(n66), 
	.B1(\ram[14][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n466));
   AO22CHD U2240 (.O(n815), 
	.B2(n66), 
	.B1(\ram[14][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n466));
   AO22CHD U2241 (.O(n816), 
	.B2(n66), 
	.B1(\ram[14][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n466));
   AO22CHD U2242 (.O(n817), 
	.B2(n66), 
	.B1(\ram[14][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n466));
   AO22CHD U2243 (.O(n818), 
	.B2(n66), 
	.B1(\ram[14][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n466));
   AO22CHD U2244 (.O(n819), 
	.B2(n66), 
	.B1(\ram[14][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n466));
   AO22CHD U2245 (.O(n820), 
	.B2(n66), 
	.B1(\ram[14][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n466));
   AO22CHD U2246 (.O(n821), 
	.B2(n66), 
	.B1(\ram[14][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n466));
   AO22CHD U2247 (.O(n822), 
	.B2(n69), 
	.B1(\ram[15][0] ), 
	.A2(n6), 
	.A1(n468));
   AO22CHD U2248 (.O(n823), 
	.B2(n69), 
	.B1(\ram[15][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n468));
   AO22CHD U2249 (.O(n824), 
	.B2(n69), 
	.B1(\ram[15][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n468));
   AO22CHD U2250 (.O(n825), 
	.B2(n69), 
	.B1(\ram[15][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n468));
   AO22CHD U2251 (.O(n826), 
	.B2(n69), 
	.B1(\ram[15][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n468));
   AO22CHD U2252 (.O(n827), 
	.B2(n69), 
	.B1(\ram[15][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n468));
   AO22CHD U2253 (.O(n828), 
	.B2(n69), 
	.B1(\ram[15][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n468));
   AO22CHD U2254 (.O(n829), 
	.B2(n69), 
	.B1(\ram[15][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n468));
   AO22CHD U2255 (.O(n830), 
	.B2(n69), 
	.B1(\ram[15][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n468));
   AO22CHD U2256 (.O(n831), 
	.B2(n69), 
	.B1(\ram[15][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n468));
   AO22CHD U2257 (.O(n832), 
	.B2(n69), 
	.B1(\ram[15][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n468));
   AO22CHD U2258 (.O(n833), 
	.B2(n69), 
	.B1(\ram[15][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n468));
   AO22CHD U2259 (.O(n834), 
	.B2(n69), 
	.B1(\ram[15][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n468));
   AO22CHD U2260 (.O(n835), 
	.B2(n69), 
	.B1(\ram[15][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n468));
   AO22CHD U2261 (.O(n836), 
	.B2(n69), 
	.B1(\ram[15][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n468));
   AO22CHD U2262 (.O(n837), 
	.B2(n69), 
	.B1(\ram[15][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n468));
   AO22CHD U2263 (.O(n838), 
	.B2(n74), 
	.B1(\ram[16][0] ), 
	.A2(n6), 
	.A1(n470));
   AO22CHD U2264 (.O(n839), 
	.B2(n74), 
	.B1(\ram[16][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n470));
   AO22CHD U2265 (.O(n840), 
	.B2(n74), 
	.B1(\ram[16][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n470));
   AO22CHD U2266 (.O(n841), 
	.B2(n74), 
	.B1(\ram[16][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n470));
   AO22CHD U2267 (.O(n842), 
	.B2(n74), 
	.B1(\ram[16][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n470));
   AO22CHD U2268 (.O(n843), 
	.B2(n74), 
	.B1(\ram[16][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n470));
   AO22CHD U2269 (.O(n844), 
	.B2(n74), 
	.B1(\ram[16][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n470));
   AO22CHD U2270 (.O(n845), 
	.B2(n74), 
	.B1(\ram[16][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n470));
   AO22CHD U2271 (.O(n846), 
	.B2(n74), 
	.B1(\ram[16][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n470));
   AO22CHD U2272 (.O(n847), 
	.B2(n74), 
	.B1(\ram[16][9] ), 
	.A2(n17), 
	.A1(n470));
   AO22CHD U2273 (.O(n848), 
	.B2(n74), 
	.B1(\ram[16][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n470));
   AO22CHD U2274 (.O(n849), 
	.B2(n74), 
	.B1(\ram[16][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n470));
   AO22CHD U2275 (.O(n850), 
	.B2(n74), 
	.B1(\ram[16][12] ), 
	.A2(n20), 
	.A1(n470));
   AO22CHD U2276 (.O(n851), 
	.B2(n74), 
	.B1(\ram[16][13] ), 
	.A2(n21), 
	.A1(n470));
   AO22CHD U2277 (.O(n852), 
	.B2(n74), 
	.B1(\ram[16][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n470));
   AO22CHD U2278 (.O(n853), 
	.B2(n74), 
	.B1(\ram[16][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n470));
   AO22CHD U2279 (.O(n854), 
	.B2(n77), 
	.B1(\ram[17][0] ), 
	.A2(n6), 
	.A1(n472));
   AO22CHD U2280 (.O(n855), 
	.B2(n77), 
	.B1(\ram[17][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n472));
   AO22CHD U2281 (.O(n856), 
	.B2(n77), 
	.B1(\ram[17][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n472));
   AO22CHD U2282 (.O(n857), 
	.B2(n77), 
	.B1(\ram[17][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n472));
   AO22CHD U2283 (.O(n858), 
	.B2(n77), 
	.B1(\ram[17][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n472));
   AO22CHD U2284 (.O(n859), 
	.B2(n77), 
	.B1(\ram[17][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n472));
   AO22CHD U2285 (.O(n860), 
	.B2(n77), 
	.B1(\ram[17][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n472));
   AO22CHD U2286 (.O(n861), 
	.B2(n77), 
	.B1(\ram[17][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n472));
   AO22CHD U2287 (.O(n862), 
	.B2(n77), 
	.B1(\ram[17][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n472));
   AO22CHD U2288 (.O(n863), 
	.B2(n77), 
	.B1(\ram[17][9] ), 
	.A2(n17), 
	.A1(n472));
   AO22CHD U2289 (.O(n864), 
	.B2(n77), 
	.B1(\ram[17][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n472));
   AO22CHD U2290 (.O(n865), 
	.B2(n77), 
	.B1(\ram[17][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n472));
   AO22CHD U2291 (.O(n866), 
	.B2(n77), 
	.B1(\ram[17][12] ), 
	.A2(n20), 
	.A1(n472));
   AO22CHD U2292 (.O(n867), 
	.B2(n77), 
	.B1(\ram[17][13] ), 
	.A2(n21), 
	.A1(n472));
   AO22CHD U2293 (.O(n868), 
	.B2(n77), 
	.B1(FE_PHN4092_ram_17__14_), 
	.A2(FE_OFN88_n22), 
	.A1(n472));
   AO22CHD U2294 (.O(n869), 
	.B2(n77), 
	.B1(\ram[17][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n472));
   AO22CHD U2295 (.O(n870), 
	.B2(n79), 
	.B1(\ram[18][0] ), 
	.A2(n6), 
	.A1(n475));
   AO22CHD U2296 (.O(n871), 
	.B2(n79), 
	.B1(\ram[18][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n475));
   AO22CHD U2297 (.O(n872), 
	.B2(n79), 
	.B1(\ram[18][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n475));
   AO22CHD U2298 (.O(n873), 
	.B2(n79), 
	.B1(\ram[18][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n475));
   AO22CHD U2299 (.O(n874), 
	.B2(n79), 
	.B1(\ram[18][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n475));
   AO22CHD U2300 (.O(n875), 
	.B2(n79), 
	.B1(\ram[18][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n475));
   AO22CHD U2301 (.O(n876), 
	.B2(n79), 
	.B1(\ram[18][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n475));
   AO22CHD U2302 (.O(n877), 
	.B2(n79), 
	.B1(\ram[18][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n475));
   AO22CHD U2303 (.O(n878), 
	.B2(n79), 
	.B1(\ram[18][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n475));
   AO22CHD U2304 (.O(n879), 
	.B2(n79), 
	.B1(\ram[18][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n475));
   AO22CHD U2305 (.O(n880), 
	.B2(n79), 
	.B1(\ram[18][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n475));
   AO22CHD U2306 (.O(n881), 
	.B2(n79), 
	.B1(\ram[18][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n475));
   AO22CHD U2307 (.O(n882), 
	.B2(n79), 
	.B1(\ram[18][12] ), 
	.A2(n20), 
	.A1(n475));
   AO22CHD U2308 (.O(n883), 
	.B2(n79), 
	.B1(\ram[18][13] ), 
	.A2(n21), 
	.A1(n475));
   AO22CHD U2309 (.O(n884), 
	.B2(n79), 
	.B1(\ram[18][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n475));
   AO22CHD U2310 (.O(n885), 
	.B2(n79), 
	.B1(\ram[18][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n475));
   AO22CHD U2311 (.O(n886), 
	.B2(n81), 
	.B1(\ram[19][0] ), 
	.A2(n6), 
	.A1(n477));
   AO22CHD U2312 (.O(n887), 
	.B2(n81), 
	.B1(\ram[19][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n477));
   AO22CHD U2313 (.O(n888), 
	.B2(n81), 
	.B1(\ram[19][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n477));
   AO22CHD U2314 (.O(n889), 
	.B2(n81), 
	.B1(\ram[19][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n477));
   AO22CHD U2315 (.O(n890), 
	.B2(n81), 
	.B1(\ram[19][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n477));
   AO22CHD U2316 (.O(n891), 
	.B2(n81), 
	.B1(\ram[19][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n477));
   AO22CHD U2317 (.O(n892), 
	.B2(n81), 
	.B1(\ram[19][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n477));
   AO22CHD U2318 (.O(n893), 
	.B2(n81), 
	.B1(\ram[19][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n477));
   AO22CHD U2319 (.O(n894), 
	.B2(n81), 
	.B1(\ram[19][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n477));
   AO22CHD U2320 (.O(n895), 
	.B2(n81), 
	.B1(\ram[19][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n477));
   AO22CHD U2321 (.O(n896), 
	.B2(n81), 
	.B1(\ram[19][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n477));
   AO22CHD U2322 (.O(n897), 
	.B2(n81), 
	.B1(\ram[19][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n477));
   AO22CHD U2323 (.O(n898), 
	.B2(n81), 
	.B1(\ram[19][12] ), 
	.A2(n20), 
	.A1(n477));
   AO22CHD U2324 (.O(n899), 
	.B2(n81), 
	.B1(\ram[19][13] ), 
	.A2(n21), 
	.A1(n477));
   AO22CHD U2325 (.O(n900), 
	.B2(n81), 
	.B1(\ram[19][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n477));
   AO22CHD U2326 (.O(n901), 
	.B2(n81), 
	.B1(\ram[19][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n477));
   AO22CHD U2327 (.O(n902), 
	.B2(n83), 
	.B1(\ram[20][0] ), 
	.A2(n6), 
	.A1(n478));
   AO22CHD U2328 (.O(n903), 
	.B2(n83), 
	.B1(\ram[20][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n478));
   AO22CHD U2329 (.O(n904), 
	.B2(n83), 
	.B1(\ram[20][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n478));
   AO22CHD U2330 (.O(n905), 
	.B2(n83), 
	.B1(\ram[20][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n478));
   AO22CHD U2331 (.O(n906), 
	.B2(n83), 
	.B1(\ram[20][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n478));
   AO22CHD U2332 (.O(n907), 
	.B2(n83), 
	.B1(\ram[20][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n478));
   AO22CHD U2333 (.O(n908), 
	.B2(n83), 
	.B1(\ram[20][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n478));
   AO22CHD U2334 (.O(n909), 
	.B2(n83), 
	.B1(\ram[20][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n478));
   AO22CHD U2335 (.O(n910), 
	.B2(n83), 
	.B1(\ram[20][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n478));
   AO22CHD U2336 (.O(n911), 
	.B2(n83), 
	.B1(\ram[20][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n478));
   AO22CHD U2337 (.O(n912), 
	.B2(n83), 
	.B1(FE_PHN4459_ram_20__10_), 
	.A2(FE_OFN73_n18), 
	.A1(n478));
   AO22CHD U2338 (.O(n913), 
	.B2(n83), 
	.B1(\ram[20][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n478));
   AO22CHD U2339 (.O(n914), 
	.B2(n83), 
	.B1(\ram[20][12] ), 
	.A2(n20), 
	.A1(n478));
   AO22CHD U2340 (.O(n915), 
	.B2(n83), 
	.B1(\ram[20][13] ), 
	.A2(n21), 
	.A1(n478));
   AO22CHD U2341 (.O(n916), 
	.B2(n83), 
	.B1(\ram[20][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n478));
   AO22CHD U2342 (.O(n917), 
	.B2(n83), 
	.B1(\ram[20][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n478));
   AO22CHD U2343 (.O(n918), 
	.B2(n85), 
	.B1(\ram[21][0] ), 
	.A2(n6), 
	.A1(n480));
   AO22CHD U2344 (.O(n919), 
	.B2(n85), 
	.B1(\ram[21][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n480));
   AO22CHD U2345 (.O(n920), 
	.B2(n85), 
	.B1(\ram[21][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n480));
   AO22CHD U2346 (.O(n921), 
	.B2(n85), 
	.B1(\ram[21][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n480));
   AO22CHD U2347 (.O(n922), 
	.B2(n85), 
	.B1(\ram[21][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n480));
   AO22CHD U2348 (.O(n923), 
	.B2(n85), 
	.B1(\ram[21][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n480));
   AO22CHD U2349 (.O(n924), 
	.B2(n85), 
	.B1(\ram[21][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n480));
   AO22CHD U2350 (.O(n925), 
	.B2(n85), 
	.B1(\ram[21][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n480));
   AO22CHD U2351 (.O(n926), 
	.B2(n85), 
	.B1(\ram[21][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n480));
   AO22CHD U2352 (.O(n927), 
	.B2(n85), 
	.B1(\ram[21][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n480));
   AO22CHD U2353 (.O(n928), 
	.B2(n85), 
	.B1(\ram[21][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n480));
   AO22CHD U2354 (.O(n929), 
	.B2(n85), 
	.B1(\ram[21][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n480));
   AO22CHD U2355 (.O(n930), 
	.B2(n85), 
	.B1(\ram[21][12] ), 
	.A2(n20), 
	.A1(n480));
   AO22CHD U2356 (.O(n931), 
	.B2(n85), 
	.B1(\ram[21][13] ), 
	.A2(n21), 
	.A1(n480));
   AO22CHD U2357 (.O(n932), 
	.B2(n85), 
	.B1(\ram[21][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n480));
   AO22CHD U2358 (.O(n933), 
	.B2(n85), 
	.B1(\ram[21][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n480));
   AO22CHD U2359 (.O(n934), 
	.B2(n87), 
	.B1(\ram[22][0] ), 
	.A2(n6), 
	.A1(n482));
   AO22CHD U2360 (.O(n935), 
	.B2(n87), 
	.B1(\ram[22][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n482));
   AO22CHD U2361 (.O(n936), 
	.B2(n87), 
	.B1(\ram[22][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n482));
   AO22CHD U2362 (.O(n937), 
	.B2(n87), 
	.B1(\ram[22][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n482));
   AO22CHD U2363 (.O(n938), 
	.B2(n87), 
	.B1(\ram[22][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n482));
   AO22CHD U2364 (.O(n939), 
	.B2(n87), 
	.B1(\ram[22][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n482));
   AO22CHD U2365 (.O(n940), 
	.B2(n87), 
	.B1(\ram[22][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n482));
   AO22CHD U2366 (.O(n941), 
	.B2(n87), 
	.B1(\ram[22][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n482));
   AO22CHD U2367 (.O(n942), 
	.B2(n87), 
	.B1(\ram[22][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n482));
   AO22CHD U2368 (.O(n943), 
	.B2(n87), 
	.B1(\ram[22][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n482));
   AO22CHD U2369 (.O(n944), 
	.B2(n87), 
	.B1(\ram[22][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n482));
   AO22CHD U2370 (.O(n945), 
	.B2(n87), 
	.B1(\ram[22][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n482));
   AO22CHD U2371 (.O(n946), 
	.B2(n87), 
	.B1(\ram[22][12] ), 
	.A2(n20), 
	.A1(n482));
   AO22CHD U2372 (.O(n947), 
	.B2(n87), 
	.B1(\ram[22][13] ), 
	.A2(n21), 
	.A1(n482));
   AO22CHD U2373 (.O(n948), 
	.B2(n87), 
	.B1(\ram[22][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n482));
   AO22CHD U2374 (.O(n949), 
	.B2(n87), 
	.B1(\ram[22][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n482));
   AO22CHD U2375 (.O(n950), 
	.B2(n89), 
	.B1(\ram[23][0] ), 
	.A2(n6), 
	.A1(n484));
   AO22CHD U2376 (.O(n951), 
	.B2(n89), 
	.B1(\ram[23][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n484));
   AO22CHD U2377 (.O(n952), 
	.B2(n89), 
	.B1(\ram[23][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n484));
   AO22CHD U2378 (.O(n953), 
	.B2(n89), 
	.B1(\ram[23][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n484));
   AO22CHD U2379 (.O(n954), 
	.B2(n89), 
	.B1(\ram[23][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n484));
   AO22CHD U2380 (.O(n955), 
	.B2(n89), 
	.B1(\ram[23][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n484));
   AO22CHD U2381 (.O(n956), 
	.B2(n89), 
	.B1(\ram[23][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n484));
   AO22CHD U2382 (.O(n957), 
	.B2(n89), 
	.B1(\ram[23][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n484));
   AO22CHD U2383 (.O(n958), 
	.B2(n89), 
	.B1(\ram[23][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n484));
   AO22CHD U2384 (.O(n959), 
	.B2(n89), 
	.B1(\ram[23][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n484));
   AO22CHD U2385 (.O(n960), 
	.B2(n89), 
	.B1(\ram[23][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n484));
   AO22CHD U2386 (.O(n961), 
	.B2(n89), 
	.B1(\ram[23][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n484));
   AO22CHD U2387 (.O(n962), 
	.B2(n89), 
	.B1(\ram[23][12] ), 
	.A2(n20), 
	.A1(n484));
   AO22CHD U2388 (.O(n963), 
	.B2(n89), 
	.B1(\ram[23][13] ), 
	.A2(n21), 
	.A1(n484));
   AO22CHD U2389 (.O(n964), 
	.B2(n89), 
	.B1(\ram[23][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n484));
   AO22CHD U2390 (.O(n965), 
	.B2(n89), 
	.B1(\ram[23][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n484));
   AO22CHD U2391 (.O(n966), 
	.B2(n91), 
	.B1(\ram[24][0] ), 
	.A2(n6), 
	.A1(n486));
   AO22CHD U2392 (.O(n967), 
	.B2(n91), 
	.B1(\ram[24][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n486));
   AO22CHD U2393 (.O(n968), 
	.B2(n91), 
	.B1(\ram[24][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n486));
   AO22CHD U2394 (.O(n969), 
	.B2(n91), 
	.B1(\ram[24][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n486));
   AO22CHD U2395 (.O(n970), 
	.B2(n91), 
	.B1(\ram[24][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n486));
   AO22CHD U2396 (.O(n971), 
	.B2(n91), 
	.B1(\ram[24][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n486));
   AO22CHD U2397 (.O(n972), 
	.B2(n91), 
	.B1(\ram[24][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n486));
   AO22CHD U2398 (.O(n973), 
	.B2(n91), 
	.B1(\ram[24][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n486));
   AO22CHD U2399 (.O(FE_PHN7451_n974), 
	.B2(n91), 
	.B1(\ram[24][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n486));
   AO22CHD U2400 (.O(n975), 
	.B2(n91), 
	.B1(\ram[24][9] ), 
	.A2(n17), 
	.A1(n486));
   AO22CHD U2401 (.O(n976), 
	.B2(n91), 
	.B1(\ram[24][10] ), 
	.A2(n18), 
	.A1(n486));
   AO22CHD U2402 (.O(n977), 
	.B2(n91), 
	.B1(\ram[24][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n486));
   AO22CHD U2403 (.O(n978), 
	.B2(n91), 
	.B1(\ram[24][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n486));
   AO22CHD U2404 (.O(n979), 
	.B2(n91), 
	.B1(\ram[24][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n486));
   AO22CHD U2405 (.O(n980), 
	.B2(n91), 
	.B1(\ram[24][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n486));
   AO22CHD U2406 (.O(n981), 
	.B2(n91), 
	.B1(\ram[24][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n486));
   AO22CHD U2407 (.O(n982), 
	.B2(n93), 
	.B1(\ram[25][0] ), 
	.A2(n6), 
	.A1(n488));
   AO22CHD U2408 (.O(n983), 
	.B2(n93), 
	.B1(\ram[25][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n488));
   AO22CHD U2409 (.O(n984), 
	.B2(n93), 
	.B1(\ram[25][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n488));
   AO22CHD U2410 (.O(n985), 
	.B2(n93), 
	.B1(\ram[25][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n488));
   AO22CHD U2411 (.O(n986), 
	.B2(n93), 
	.B1(\ram[25][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n488));
   AO22CHD U2412 (.O(n987), 
	.B2(n93), 
	.B1(\ram[25][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n488));
   AO22CHD U2413 (.O(n988), 
	.B2(n93), 
	.B1(\ram[25][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n488));
   AO22CHD U2414 (.O(n989), 
	.B2(n93), 
	.B1(\ram[25][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n488));
   AO22CHD U2415 (.O(n990), 
	.B2(n93), 
	.B1(\ram[25][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n488));
   AO22CHD U2416 (.O(n991), 
	.B2(n93), 
	.B1(\ram[25][9] ), 
	.A2(n17), 
	.A1(n488));
   AO22CHD U2417 (.O(n992), 
	.B2(n93), 
	.B1(\ram[25][10] ), 
	.A2(n18), 
	.A1(n488));
   AO22CHD U2418 (.O(n993), 
	.B2(n93), 
	.B1(\ram[25][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n488));
   AO22CHD U2419 (.O(n994), 
	.B2(n93), 
	.B1(\ram[25][12] ), 
	.A2(n20), 
	.A1(n488));
   AO22CHD U2420 (.O(n995), 
	.B2(n93), 
	.B1(\ram[25][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n488));
   AO22CHD U2421 (.O(n996), 
	.B2(n93), 
	.B1(\ram[25][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n488));
   AO22CHD U2422 (.O(n997), 
	.B2(n93), 
	.B1(\ram[25][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n488));
   AO22CHD U2423 (.O(n998), 
	.B2(n95), 
	.B1(\ram[26][0] ), 
	.A2(n6), 
	.A1(n490));
   AO22CHD U2424 (.O(n999), 
	.B2(n95), 
	.B1(\ram[26][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n490));
   AO22CHD U2425 (.O(n1000), 
	.B2(n95), 
	.B1(\ram[26][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n490));
   AO22CHD U2426 (.O(n1001), 
	.B2(n95), 
	.B1(\ram[26][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n490));
   AO22CHD U2427 (.O(n1002), 
	.B2(n95), 
	.B1(\ram[26][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n490));
   AO22CHD U2428 (.O(n1003), 
	.B2(n95), 
	.B1(\ram[26][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n490));
   AO22CHD U2429 (.O(n1004), 
	.B2(n95), 
	.B1(\ram[26][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n490));
   AO22CHD U2430 (.O(n1005), 
	.B2(n95), 
	.B1(\ram[26][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n490));
   AO22CHD U2431 (.O(n1006), 
	.B2(n95), 
	.B1(\ram[26][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n490));
   AO22CHD U2432 (.O(n1007), 
	.B2(n95), 
	.B1(\ram[26][9] ), 
	.A2(n17), 
	.A1(n490));
   AO22CHD U2433 (.O(n1008), 
	.B2(n95), 
	.B1(\ram[26][10] ), 
	.A2(n18), 
	.A1(n490));
   AO22CHD U2434 (.O(n1009), 
	.B2(n95), 
	.B1(\ram[26][11] ), 
	.A2(n19), 
	.A1(n490));
   AO22CHD U2435 (.O(n1010), 
	.B2(n95), 
	.B1(\ram[26][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n490));
   AO22CHD U2436 (.O(n1011), 
	.B2(n95), 
	.B1(\ram[26][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n490));
   AO22CHD U2437 (.O(n1012), 
	.B2(n95), 
	.B1(\ram[26][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n490));
   AO22CHD U2438 (.O(FE_PHN7495_n1013), 
	.B2(n95), 
	.B1(\ram[26][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n490));
   AO22CHD U2439 (.O(FE_PHN7449_n1014), 
	.B2(n97), 
	.B1(\ram[27][0] ), 
	.A2(n6), 
	.A1(n492));
   AO22CHD U2440 (.O(n1015), 
	.B2(n97), 
	.B1(\ram[27][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n492));
   AO22CHD U2441 (.O(n1016), 
	.B2(n97), 
	.B1(\ram[27][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n492));
   AO22CHD U2442 (.O(n1017), 
	.B2(n97), 
	.B1(\ram[27][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n492));
   AO22CHD U2443 (.O(n1018), 
	.B2(n97), 
	.B1(\ram[27][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n492));
   AO22CHD U2444 (.O(n1019), 
	.B2(n97), 
	.B1(\ram[27][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n492));
   AO22CHD U2445 (.O(n1020), 
	.B2(n97), 
	.B1(\ram[27][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n492));
   AO22CHD U2446 (.O(n1021), 
	.B2(n97), 
	.B1(\ram[27][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n492));
   AO22CHD U2447 (.O(n1022), 
	.B2(n97), 
	.B1(\ram[27][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n492));
   AO22CHD U2448 (.O(n1023), 
	.B2(n97), 
	.B1(\ram[27][9] ), 
	.A2(n17), 
	.A1(n492));
   AO22CHD U2449 (.O(n1024), 
	.B2(n97), 
	.B1(\ram[27][10] ), 
	.A2(n18), 
	.A1(n492));
   AO22CHD U2450 (.O(n1025), 
	.B2(n97), 
	.B1(\ram[27][11] ), 
	.A2(n19), 
	.A1(n492));
   AO22CHD U2451 (.O(n1026), 
	.B2(n97), 
	.B1(\ram[27][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n492));
   AO22CHD U2452 (.O(n1027), 
	.B2(n97), 
	.B1(\ram[27][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n492));
   AO22CHD U2453 (.O(n1028), 
	.B2(n97), 
	.B1(\ram[27][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n492));
   AO22CHD U2454 (.O(n1029), 
	.B2(n97), 
	.B1(\ram[27][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n492));
   AO22CHD U2455 (.O(n1030), 
	.B2(n99), 
	.B1(\ram[28][0] ), 
	.A2(n6), 
	.A1(n494));
   AO22CHD U2456 (.O(n1031), 
	.B2(n99), 
	.B1(\ram[28][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n494));
   AO22CHD U2457 (.O(n1032), 
	.B2(n99), 
	.B1(\ram[28][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n494));
   AO22CHD U2458 (.O(n1033), 
	.B2(n99), 
	.B1(\ram[28][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n494));
   AO22CHD U2459 (.O(n1034), 
	.B2(n99), 
	.B1(\ram[28][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n494));
   AO22CHD U2460 (.O(n1035), 
	.B2(n99), 
	.B1(\ram[28][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n494));
   AO22CHD U2461 (.O(n1036), 
	.B2(n99), 
	.B1(\ram[28][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n494));
   AO22CHD U2462 (.O(n1037), 
	.B2(n99), 
	.B1(\ram[28][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n494));
   AO22CHD U2463 (.O(n1038), 
	.B2(n99), 
	.B1(\ram[28][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n494));
   AO22CHD U2464 (.O(n1039), 
	.B2(n99), 
	.B1(\ram[28][9] ), 
	.A2(n17), 
	.A1(n494));
   AO22CHD U2465 (.O(n1040), 
	.B2(n99), 
	.B1(\ram[28][10] ), 
	.A2(n18), 
	.A1(n494));
   AO22CHD U2466 (.O(n1041), 
	.B2(n99), 
	.B1(\ram[28][11] ), 
	.A2(n19), 
	.A1(n494));
   AO22CHD U2467 (.O(n1042), 
	.B2(n99), 
	.B1(\ram[28][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n494));
   AO22CHD U2468 (.O(n1043), 
	.B2(n99), 
	.B1(\ram[28][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n494));
   AO22CHD U2469 (.O(n1044), 
	.B2(n99), 
	.B1(\ram[28][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n494));
   AO22CHD U2470 (.O(n1045), 
	.B2(n99), 
	.B1(\ram[28][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n494));
   AO22CHD U2471 (.O(n1046), 
	.B2(n101), 
	.B1(\ram[29][0] ), 
	.A2(n6), 
	.A1(n496));
   AO22CHD U2472 (.O(n1047), 
	.B2(n101), 
	.B1(\ram[29][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n496));
   AO22CHD U2473 (.O(n1048), 
	.B2(n101), 
	.B1(\ram[29][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n496));
   AO22CHD U2474 (.O(n1049), 
	.B2(n101), 
	.B1(\ram[29][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n496));
   AO22CHD U2475 (.O(n1050), 
	.B2(n101), 
	.B1(\ram[29][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n496));
   AO22CHD U2476 (.O(n1051), 
	.B2(n101), 
	.B1(\ram[29][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n496));
   AO22CHD U2477 (.O(n1052), 
	.B2(n101), 
	.B1(\ram[29][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n496));
   AO22CHD U2478 (.O(n1053), 
	.B2(n101), 
	.B1(\ram[29][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n496));
   AO22CHD U2479 (.O(n1054), 
	.B2(n101), 
	.B1(\ram[29][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n496));
   AO22CHD U2480 (.O(n1055), 
	.B2(n101), 
	.B1(\ram[29][9] ), 
	.A2(n17), 
	.A1(n496));
   AO22CHD U2481 (.O(n1056), 
	.B2(n101), 
	.B1(\ram[29][10] ), 
	.A2(n18), 
	.A1(n496));
   AO22CHD U2482 (.O(n1057), 
	.B2(n101), 
	.B1(\ram[29][11] ), 
	.A2(n19), 
	.A1(n496));
   AO22CHD U2483 (.O(n1058), 
	.B2(n101), 
	.B1(\ram[29][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n496));
   AO22CHD U2484 (.O(n1059), 
	.B2(n101), 
	.B1(\ram[29][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n496));
   AO22CHD U2485 (.O(n1060), 
	.B2(n101), 
	.B1(FE_PHN516_ram_29__14_), 
	.A2(FE_OFN88_n22), 
	.A1(n496));
   AO22CHD U2486 (.O(n1061), 
	.B2(n101), 
	.B1(\ram[29][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n496));
   AO22CHD U2487 (.O(n1062), 
	.B2(n103), 
	.B1(\ram[30][0] ), 
	.A2(n6), 
	.A1(n498));
   AO22CHD U2488 (.O(n1063), 
	.B2(n103), 
	.B1(\ram[30][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n498));
   AO22CHD U2489 (.O(n1064), 
	.B2(n103), 
	.B1(\ram[30][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n498));
   AO22CHD U2490 (.O(n1065), 
	.B2(n103), 
	.B1(\ram[30][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n498));
   AO22CHD U2491 (.O(n1066), 
	.B2(n103), 
	.B1(\ram[30][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n498));
   AO22CHD U2492 (.O(n1067), 
	.B2(n103), 
	.B1(\ram[30][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n498));
   AO22CHD U2493 (.O(n1068), 
	.B2(n103), 
	.B1(\ram[30][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n498));
   AO22CHD U2494 (.O(n1069), 
	.B2(n103), 
	.B1(\ram[30][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n498));
   AO22CHD U2495 (.O(n1070), 
	.B2(n103), 
	.B1(\ram[30][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n498));
   AO22CHD U2496 (.O(n1071), 
	.B2(n103), 
	.B1(\ram[30][9] ), 
	.A2(n17), 
	.A1(n498));
   AO22CHD U2497 (.O(n1072), 
	.B2(n103), 
	.B1(\ram[30][10] ), 
	.A2(n18), 
	.A1(n498));
   AO22CHD U2498 (.O(n1073), 
	.B2(n103), 
	.B1(\ram[30][11] ), 
	.A2(n19), 
	.A1(n498));
   AO22CHD U2499 (.O(n1074), 
	.B2(n103), 
	.B1(\ram[30][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n498));
   AO22CHD U2500 (.O(n1075), 
	.B2(n103), 
	.B1(\ram[30][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n498));
   AO22CHD U2501 (.O(n1076), 
	.B2(n103), 
	.B1(\ram[30][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n498));
   AO22CHD U2502 (.O(n1077), 
	.B2(n103), 
	.B1(\ram[30][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n498));
   AO22CHD U2503 (.O(n1078), 
	.B2(n105), 
	.B1(\ram[31][0] ), 
	.A2(n6), 
	.A1(n500));
   AO22CHD U2504 (.O(n1079), 
	.B2(n105), 
	.B1(\ram[31][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n500));
   AO22CHD U2505 (.O(n1080), 
	.B2(n105), 
	.B1(FE_PHN5410_ram_31__2_), 
	.A2(FE_OFN47_n10), 
	.A1(n500));
   AO22CHD U2506 (.O(n1081), 
	.B2(n105), 
	.B1(\ram[31][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n500));
   AO22CHD U2507 (.O(n1082), 
	.B2(n105), 
	.B1(\ram[31][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n500));
   AO22CHD U2508 (.O(n1083), 
	.B2(n105), 
	.B1(\ram[31][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n500));
   AO22CHD U2509 (.O(n1084), 
	.B2(n105), 
	.B1(\ram[31][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n500));
   AO22CHD U2510 (.O(n1085), 
	.B2(n105), 
	.B1(\ram[31][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n500));
   AO22CHD U2511 (.O(n1086), 
	.B2(n105), 
	.B1(\ram[31][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n500));
   AO22CHD U2512 (.O(n1087), 
	.B2(n105), 
	.B1(\ram[31][9] ), 
	.A2(n17), 
	.A1(n500));
   AO22CHD U2513 (.O(n1088), 
	.B2(n105), 
	.B1(\ram[31][10] ), 
	.A2(n18), 
	.A1(n500));
   AO22CHD U2514 (.O(n1089), 
	.B2(n105), 
	.B1(\ram[31][11] ), 
	.A2(n19), 
	.A1(n500));
   AO22CHD U2515 (.O(n1090), 
	.B2(n105), 
	.B1(\ram[31][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n500));
   AO22CHD U2516 (.O(n1091), 
	.B2(n105), 
	.B1(\ram[31][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n500));
   AO22CHD U2517 (.O(n1092), 
	.B2(n105), 
	.B1(\ram[31][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n500));
   AO22CHD U2518 (.O(n1093), 
	.B2(n105), 
	.B1(\ram[31][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n500));
   AO22CHD U2519 (.O(n1094), 
	.B2(n108), 
	.B1(\ram[32][0] ), 
	.A2(n6), 
	.A1(n502));
   AO22CHD U2520 (.O(n1095), 
	.B2(n108), 
	.B1(\ram[32][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n502));
   AO22CHD U2521 (.O(n1096), 
	.B2(n108), 
	.B1(\ram[32][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n502));
   AO22CHD U2522 (.O(n1097), 
	.B2(n108), 
	.B1(\ram[32][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n502));
   AO22CHD U2523 (.O(n1098), 
	.B2(n108), 
	.B1(\ram[32][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n502));
   AO22CHD U2524 (.O(n1099), 
	.B2(n108), 
	.B1(\ram[32][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n502));
   AO22CHD U2525 (.O(n1100), 
	.B2(n108), 
	.B1(\ram[32][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n502));
   AO22CHD U2526 (.O(n1101), 
	.B2(n108), 
	.B1(\ram[32][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n502));
   AO22CHD U2527 (.O(n1102), 
	.B2(n108), 
	.B1(\ram[32][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n502));
   AO22CHD U2528 (.O(n1103), 
	.B2(n108), 
	.B1(\ram[32][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n502));
   AO22CHD U2529 (.O(n1104), 
	.B2(n108), 
	.B1(\ram[32][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n502));
   AO22CHD U2530 (.O(n1105), 
	.B2(n108), 
	.B1(\ram[32][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n502));
   AO22CHD U2531 (.O(n1106), 
	.B2(n108), 
	.B1(\ram[32][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n502));
   AO22CHD U2532 (.O(n1107), 
	.B2(n108), 
	.B1(\ram[32][13] ), 
	.A2(n21), 
	.A1(n502));
   AO22CHD U2533 (.O(n1108), 
	.B2(n108), 
	.B1(\ram[32][14] ), 
	.A2(n22), 
	.A1(n502));
   AO22CHD U2534 (.O(n1109), 
	.B2(n108), 
	.B1(\ram[32][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n502));
   AO22CHD U2535 (.O(n1110), 
	.B2(n111), 
	.B1(\ram[33][0] ), 
	.A2(n6), 
	.A1(n504));
   AO22CHD U2536 (.O(n1111), 
	.B2(n111), 
	.B1(\ram[33][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n504));
   AO22CHD U2537 (.O(n1112), 
	.B2(n111), 
	.B1(\ram[33][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n504));
   AO22CHD U2538 (.O(n1113), 
	.B2(n111), 
	.B1(\ram[33][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n504));
   AO22CHD U2539 (.O(n1114), 
	.B2(n111), 
	.B1(\ram[33][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n504));
   AO22CHD U2540 (.O(n1115), 
	.B2(n111), 
	.B1(\ram[33][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n504));
   AO22CHD U2541 (.O(n1116), 
	.B2(n111), 
	.B1(\ram[33][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n504));
   AO22CHD U2542 (.O(n1117), 
	.B2(n111), 
	.B1(\ram[33][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n504));
   AO22CHD U2543 (.O(n1118), 
	.B2(n111), 
	.B1(\ram[33][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n504));
   AO22CHD U2544 (.O(n1119), 
	.B2(n111), 
	.B1(FE_PHN2658_ram_33__9_), 
	.A2(FE_OFN70_n17), 
	.A1(n504));
   AO22CHD U2545 (.O(n1120), 
	.B2(n111), 
	.B1(\ram[33][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n504));
   AO22CHD U2546 (.O(n1121), 
	.B2(n111), 
	.B1(\ram[33][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n504));
   AO22CHD U2547 (.O(n1122), 
	.B2(n111), 
	.B1(\ram[33][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n504));
   AO22CHD U2548 (.O(n1123), 
	.B2(n111), 
	.B1(\ram[33][13] ), 
	.A2(n21), 
	.A1(n504));
   AO22CHD U2549 (.O(n1124), 
	.B2(n111), 
	.B1(\ram[33][14] ), 
	.A2(n22), 
	.A1(n504));
   AO22CHD U2550 (.O(n1125), 
	.B2(n111), 
	.B1(\ram[33][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n504));
   AO22CHD U2551 (.O(n1126), 
	.B2(n113), 
	.B1(\ram[34][0] ), 
	.A2(n6), 
	.A1(n506));
   AO22CHD U2552 (.O(n1127), 
	.B2(n113), 
	.B1(\ram[34][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n506));
   AO22CHD U2553 (.O(n1128), 
	.B2(n113), 
	.B1(\ram[34][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n506));
   AO22CHD U2554 (.O(n1129), 
	.B2(n113), 
	.B1(\ram[34][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n506));
   AO22CHD U2555 (.O(n1130), 
	.B2(n113), 
	.B1(\ram[34][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n506));
   AO22CHD U2556 (.O(n1131), 
	.B2(n113), 
	.B1(\ram[34][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n506));
   AO22CHD U2557 (.O(n1132), 
	.B2(n113), 
	.B1(\ram[34][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n506));
   AO22CHD U2558 (.O(n1133), 
	.B2(n113), 
	.B1(\ram[34][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n506));
   AO22CHD U2559 (.O(n1134), 
	.B2(n113), 
	.B1(\ram[34][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n506));
   AO22CHD U2560 (.O(n1135), 
	.B2(n113), 
	.B1(\ram[34][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n506));
   AO22CHD U2561 (.O(n1136), 
	.B2(n113), 
	.B1(\ram[34][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n506));
   AO22CHD U2562 (.O(n1137), 
	.B2(n113), 
	.B1(\ram[34][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n506));
   AO22CHD U2563 (.O(n1138), 
	.B2(n113), 
	.B1(\ram[34][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n506));
   AO22CHD U2564 (.O(n1139), 
	.B2(n113), 
	.B1(\ram[34][13] ), 
	.A2(n21), 
	.A1(n506));
   AO22CHD U2565 (.O(n1140), 
	.B2(n113), 
	.B1(\ram[34][14] ), 
	.A2(n22), 
	.A1(n506));
   AO22CHD U2566 (.O(n1141), 
	.B2(n113), 
	.B1(\ram[34][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n506));
   AO22CHD U2567 (.O(n1142), 
	.B2(n115), 
	.B1(\ram[35][0] ), 
	.A2(n6), 
	.A1(n508));
   AO22CHD U2568 (.O(n1143), 
	.B2(n115), 
	.B1(\ram[35][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n508));
   AO22CHD U2569 (.O(n1144), 
	.B2(n115), 
	.B1(\ram[35][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n508));
   AO22CHD U2570 (.O(n1145), 
	.B2(n115), 
	.B1(\ram[35][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n508));
   AO22CHD U2571 (.O(n1146), 
	.B2(n115), 
	.B1(\ram[35][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n508));
   AO22CHD U2572 (.O(n1147), 
	.B2(n115), 
	.B1(\ram[35][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n508));
   AO22CHD U2573 (.O(n1148), 
	.B2(n115), 
	.B1(\ram[35][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n508));
   AO22CHD U2574 (.O(n1149), 
	.B2(n115), 
	.B1(\ram[35][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n508));
   AO22CHD U2575 (.O(n1150), 
	.B2(n115), 
	.B1(\ram[35][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n508));
   AO22CHD U2576 (.O(n1151), 
	.B2(n115), 
	.B1(\ram[35][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n508));
   AO22CHD U2577 (.O(n1152), 
	.B2(n115), 
	.B1(\ram[35][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n508));
   AO22CHD U2578 (.O(n1153), 
	.B2(n115), 
	.B1(\ram[35][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n508));
   AO22CHD U2579 (.O(n1154), 
	.B2(n115), 
	.B1(\ram[35][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n508));
   AO22CHD U2580 (.O(n1155), 
	.B2(n115), 
	.B1(\ram[35][13] ), 
	.A2(n21), 
	.A1(n508));
   AO22CHD U2581 (.O(n1156), 
	.B2(n115), 
	.B1(\ram[35][14] ), 
	.A2(n22), 
	.A1(n508));
   AO22CHD U2582 (.O(n1157), 
	.B2(n115), 
	.B1(\ram[35][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n508));
   AO22CHD U2583 (.O(n1158), 
	.B2(n117), 
	.B1(\ram[36][0] ), 
	.A2(n6), 
	.A1(n510));
   AO22CHD U2584 (.O(n1159), 
	.B2(n117), 
	.B1(\ram[36][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n510));
   AO22CHD U2585 (.O(n1160), 
	.B2(n117), 
	.B1(\ram[36][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n510));
   AO22CHD U2586 (.O(n1161), 
	.B2(n117), 
	.B1(\ram[36][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n510));
   AO22CHD U2587 (.O(n1162), 
	.B2(n117), 
	.B1(\ram[36][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n510));
   AO22CHD U2588 (.O(n1163), 
	.B2(n117), 
	.B1(\ram[36][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n510));
   AO22CHD U2589 (.O(n1164), 
	.B2(n117), 
	.B1(\ram[36][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n510));
   AO22CHD U2590 (.O(n1165), 
	.B2(n117), 
	.B1(\ram[36][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n510));
   AO22CHD U2591 (.O(n1166), 
	.B2(n117), 
	.B1(\ram[36][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n510));
   AO22CHD U2592 (.O(n1167), 
	.B2(n117), 
	.B1(\ram[36][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n510));
   AO22CHD U2593 (.O(n1168), 
	.B2(n117), 
	.B1(\ram[36][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n510));
   AO22CHD U2594 (.O(n1169), 
	.B2(n117), 
	.B1(\ram[36][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n510));
   AO22CHD U2595 (.O(n1170), 
	.B2(n117), 
	.B1(\ram[36][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n510));
   AO22CHD U2596 (.O(n1171), 
	.B2(n117), 
	.B1(\ram[36][13] ), 
	.A2(n21), 
	.A1(n510));
   AO22CHD U2597 (.O(n1172), 
	.B2(n117), 
	.B1(\ram[36][14] ), 
	.A2(n22), 
	.A1(n510));
   AO22CHD U2598 (.O(n1173), 
	.B2(n117), 
	.B1(\ram[36][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n510));
   AO22CHD U2599 (.O(n1174), 
	.B2(n119), 
	.B1(\ram[37][0] ), 
	.A2(n6), 
	.A1(n511));
   AO22CHD U2600 (.O(n1175), 
	.B2(n119), 
	.B1(\ram[37][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n511));
   AO22CHD U2601 (.O(n1176), 
	.B2(n119), 
	.B1(\ram[37][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n511));
   AO22CHD U2602 (.O(n1177), 
	.B2(n119), 
	.B1(\ram[37][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n511));
   AO22CHD U2603 (.O(n1178), 
	.B2(n119), 
	.B1(\ram[37][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n511));
   AO22CHD U2604 (.O(n1179), 
	.B2(n119), 
	.B1(\ram[37][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n511));
   AO22CHD U2605 (.O(n1180), 
	.B2(n119), 
	.B1(\ram[37][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n511));
   AO22CHD U2606 (.O(n1181), 
	.B2(n119), 
	.B1(\ram[37][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n511));
   AO22CHD U2607 (.O(n1182), 
	.B2(n119), 
	.B1(\ram[37][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n511));
   AO22CHD U2608 (.O(n1183), 
	.B2(n119), 
	.B1(\ram[37][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n511));
   AO22CHD U2609 (.O(n1184), 
	.B2(n119), 
	.B1(\ram[37][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n511));
   AO22CHD U2610 (.O(n1185), 
	.B2(n119), 
	.B1(\ram[37][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n511));
   AO22CHD U2611 (.O(n1186), 
	.B2(n119), 
	.B1(\ram[37][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n511));
   AO22CHD U2612 (.O(n1187), 
	.B2(n119), 
	.B1(\ram[37][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n511));
   AO22CHD U2613 (.O(n1188), 
	.B2(n119), 
	.B1(\ram[37][14] ), 
	.A2(n22), 
	.A1(n511));
   AO22CHD U2614 (.O(n1189), 
	.B2(n119), 
	.B1(\ram[37][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n511));
   AO22CHD U2615 (.O(n1190), 
	.B2(n121), 
	.B1(\ram[38][0] ), 
	.A2(n6), 
	.A1(n513));
   AO22CHD U2616 (.O(n1191), 
	.B2(n121), 
	.B1(\ram[38][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n513));
   AO22CHD U2617 (.O(n1192), 
	.B2(n121), 
	.B1(\ram[38][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n513));
   AO22CHD U2618 (.O(n1193), 
	.B2(n121), 
	.B1(\ram[38][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n513));
   AO22CHD U2619 (.O(n1194), 
	.B2(n121), 
	.B1(\ram[38][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n513));
   AO22CHD U2620 (.O(n1195), 
	.B2(n121), 
	.B1(\ram[38][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n513));
   AO22CHD U2621 (.O(n1196), 
	.B2(n121), 
	.B1(\ram[38][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n513));
   AO22CHD U2622 (.O(n1197), 
	.B2(n121), 
	.B1(\ram[38][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n513));
   AO22CHD U2623 (.O(n1198), 
	.B2(n121), 
	.B1(\ram[38][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n513));
   AO22CHD U2624 (.O(n1199), 
	.B2(n121), 
	.B1(\ram[38][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n513));
   AO22CHD U2625 (.O(n1200), 
	.B2(n121), 
	.B1(\ram[38][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n513));
   AO22CHD U2626 (.O(n1201), 
	.B2(n121), 
	.B1(\ram[38][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n513));
   AO22CHD U2627 (.O(n1202), 
	.B2(n121), 
	.B1(\ram[38][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n513));
   AO22CHD U2628 (.O(n1203), 
	.B2(n121), 
	.B1(\ram[38][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n513));
   AO22CHD U2629 (.O(n1204), 
	.B2(n121), 
	.B1(\ram[38][14] ), 
	.A2(n22), 
	.A1(n513));
   AO22CHD U2630 (.O(n1205), 
	.B2(n121), 
	.B1(\ram[38][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n513));
   AO22CHD U2631 (.O(n1206), 
	.B2(n123), 
	.B1(\ram[39][0] ), 
	.A2(n6), 
	.A1(n515));
   AO22CHD U2632 (.O(n1207), 
	.B2(n123), 
	.B1(\ram[39][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n515));
   AO22CHD U2633 (.O(n1208), 
	.B2(n123), 
	.B1(\ram[39][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n515));
   AO22CHD U2634 (.O(n1209), 
	.B2(n123), 
	.B1(\ram[39][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n515));
   AO22CHD U2635 (.O(n1210), 
	.B2(n123), 
	.B1(\ram[39][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n515));
   AO22CHD U2636 (.O(n1211), 
	.B2(n123), 
	.B1(\ram[39][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n515));
   AO22CHD U2637 (.O(n1212), 
	.B2(n123), 
	.B1(\ram[39][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n515));
   AO22CHD U2638 (.O(n1213), 
	.B2(n123), 
	.B1(\ram[39][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n515));
   AO22CHD U2639 (.O(n1214), 
	.B2(n123), 
	.B1(\ram[39][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n515));
   AO22CHD U2640 (.O(n1215), 
	.B2(n123), 
	.B1(\ram[39][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n515));
   AO22CHD U2641 (.O(n1216), 
	.B2(n123), 
	.B1(\ram[39][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n515));
   AO22CHD U2642 (.O(n1217), 
	.B2(n123), 
	.B1(\ram[39][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n515));
   AO22CHD U2643 (.O(n1218), 
	.B2(n123), 
	.B1(\ram[39][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n515));
   AO22CHD U2644 (.O(n1219), 
	.B2(n123), 
	.B1(\ram[39][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n515));
   AO22CHD U2645 (.O(n1220), 
	.B2(n123), 
	.B1(\ram[39][14] ), 
	.A2(n22), 
	.A1(n515));
   AO22CHD U2646 (.O(n1221), 
	.B2(n123), 
	.B1(\ram[39][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n515));
   AO22CHD U2647 (.O(n1222), 
	.B2(n125), 
	.B1(\ram[40][0] ), 
	.A2(n6), 
	.A1(n517));
   AO22CHD U2648 (.O(n1223), 
	.B2(n125), 
	.B1(\ram[40][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n517));
   AO22CHD U2649 (.O(n1224), 
	.B2(n125), 
	.B1(\ram[40][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n517));
   AO22CHD U2650 (.O(n1225), 
	.B2(n125), 
	.B1(\ram[40][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n517));
   AO22CHD U2651 (.O(n1226), 
	.B2(n125), 
	.B1(\ram[40][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n517));
   AO22CHD U2652 (.O(n1227), 
	.B2(n125), 
	.B1(\ram[40][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n517));
   AO22CHD U2653 (.O(n1228), 
	.B2(n125), 
	.B1(\ram[40][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n517));
   AO22CHD U2654 (.O(n1229), 
	.B2(n125), 
	.B1(\ram[40][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n517));
   AO22CHD U2655 (.O(n1230), 
	.B2(n125), 
	.B1(\ram[40][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n517));
   AO22CHD U2656 (.O(n1231), 
	.B2(n125), 
	.B1(\ram[40][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n517));
   AO22CHD U2657 (.O(n1232), 
	.B2(n125), 
	.B1(\ram[40][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n517));
   AO22CHD U2658 (.O(n1233), 
	.B2(n125), 
	.B1(\ram[40][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n517));
   AO22CHD U2659 (.O(n1234), 
	.B2(n125), 
	.B1(\ram[40][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n517));
   AO22CHD U2660 (.O(n1235), 
	.B2(n125), 
	.B1(\ram[40][13] ), 
	.A2(n21), 
	.A1(n517));
   AO22CHD U2661 (.O(n1236), 
	.B2(n125), 
	.B1(\ram[40][14] ), 
	.A2(n22), 
	.A1(n517));
   AO22CHD U2662 (.O(n1237), 
	.B2(n125), 
	.B1(\ram[40][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n517));
   AO22CHD U2663 (.O(n1238), 
	.B2(n127), 
	.B1(\ram[41][0] ), 
	.A2(n6), 
	.A1(n519));
   AO22CHD U2664 (.O(n1239), 
	.B2(n127), 
	.B1(\ram[41][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n519));
   AO22CHD U2665 (.O(n1240), 
	.B2(n127), 
	.B1(\ram[41][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n519));
   AO22CHD U2666 (.O(n1241), 
	.B2(n127), 
	.B1(\ram[41][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n519));
   AO22CHD U2667 (.O(n1242), 
	.B2(n127), 
	.B1(\ram[41][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n519));
   AO22CHD U2668 (.O(n1243), 
	.B2(n127), 
	.B1(\ram[41][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n519));
   AO22CHD U2669 (.O(n1244), 
	.B2(n127), 
	.B1(\ram[41][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n519));
   AO22CHD U2670 (.O(n1245), 
	.B2(n127), 
	.B1(\ram[41][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n519));
   AO22CHD U2671 (.O(n1246), 
	.B2(n127), 
	.B1(\ram[41][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n519));
   AO22CHD U2672 (.O(n1247), 
	.B2(n127), 
	.B1(\ram[41][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n519));
   AO22CHD U2673 (.O(n1248), 
	.B2(n127), 
	.B1(\ram[41][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n519));
   AO22CHD U2674 (.O(n1249), 
	.B2(n127), 
	.B1(\ram[41][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n519));
   AO22CHD U2675 (.O(n1250), 
	.B2(n127), 
	.B1(\ram[41][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n519));
   AO22CHD U2676 (.O(n1251), 
	.B2(n127), 
	.B1(\ram[41][13] ), 
	.A2(n21), 
	.A1(n519));
   AO22CHD U2677 (.O(n1252), 
	.B2(n127), 
	.B1(\ram[41][14] ), 
	.A2(n22), 
	.A1(n519));
   AO22CHD U2678 (.O(n1253), 
	.B2(n127), 
	.B1(\ram[41][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n519));
   AO22CHD U2679 (.O(n1254), 
	.B2(n129), 
	.B1(\ram[42][0] ), 
	.A2(n6), 
	.A1(n521));
   AO22CHD U2680 (.O(n1255), 
	.B2(n129), 
	.B1(\ram[42][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n521));
   AO22CHD U2681 (.O(n1256), 
	.B2(n129), 
	.B1(\ram[42][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n521));
   AO22CHD U2682 (.O(n1257), 
	.B2(n129), 
	.B1(\ram[42][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n521));
   AO22CHD U2683 (.O(n1258), 
	.B2(n129), 
	.B1(\ram[42][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n521));
   AO22CHD U2684 (.O(n1259), 
	.B2(n129), 
	.B1(\ram[42][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n521));
   AO22CHD U2685 (.O(n1260), 
	.B2(n129), 
	.B1(\ram[42][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n521));
   AO22CHD U2686 (.O(n1261), 
	.B2(n129), 
	.B1(\ram[42][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n521));
   AO22CHD U2687 (.O(n1262), 
	.B2(n129), 
	.B1(\ram[42][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n521));
   AO22CHD U2688 (.O(n1263), 
	.B2(n129), 
	.B1(\ram[42][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n521));
   AO22CHD U2689 (.O(n1264), 
	.B2(n129), 
	.B1(\ram[42][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n521));
   AO22CHD U2690 (.O(n1265), 
	.B2(n129), 
	.B1(\ram[42][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n521));
   AO22CHD U2691 (.O(n1266), 
	.B2(n129), 
	.B1(\ram[42][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n521));
   AO22CHD U2692 (.O(n1267), 
	.B2(n129), 
	.B1(\ram[42][13] ), 
	.A2(n21), 
	.A1(n521));
   AO22CHD U2693 (.O(n1268), 
	.B2(n129), 
	.B1(\ram[42][14] ), 
	.A2(n22), 
	.A1(n521));
   AO22CHD U2694 (.O(n1269), 
	.B2(n129), 
	.B1(\ram[42][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n521));
   AO22CHD U2695 (.O(n1270), 
	.B2(n131), 
	.B1(\ram[43][0] ), 
	.A2(n6), 
	.A1(n523));
   AO22CHD U2696 (.O(n1271), 
	.B2(n131), 
	.B1(\ram[43][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n523));
   AO22CHD U2697 (.O(n1272), 
	.B2(n131), 
	.B1(\ram[43][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n523));
   AO22CHD U2698 (.O(n1273), 
	.B2(n131), 
	.B1(\ram[43][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n523));
   AO22CHD U2699 (.O(n1274), 
	.B2(n131), 
	.B1(\ram[43][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n523));
   AO22CHD U2700 (.O(n1275), 
	.B2(n131), 
	.B1(\ram[43][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n523));
   AO22CHD U2701 (.O(n1276), 
	.B2(n131), 
	.B1(\ram[43][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n523));
   AO22CHD U2702 (.O(n1277), 
	.B2(n131), 
	.B1(\ram[43][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n523));
   AO22CHD U2703 (.O(n1278), 
	.B2(n131), 
	.B1(\ram[43][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n523));
   AO22CHD U2704 (.O(n1279), 
	.B2(n131), 
	.B1(\ram[43][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n523));
   AO22CHD U2705 (.O(n1280), 
	.B2(n131), 
	.B1(\ram[43][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n523));
   AO22CHD U2706 (.O(n1281), 
	.B2(n131), 
	.B1(\ram[43][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n523));
   AO22CHD U2707 (.O(n1282), 
	.B2(n131), 
	.B1(\ram[43][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n523));
   AO22CHD U2708 (.O(n1283), 
	.B2(n131), 
	.B1(\ram[43][13] ), 
	.A2(n21), 
	.A1(n523));
   AO22CHD U2709 (.O(n1284), 
	.B2(n131), 
	.B1(\ram[43][14] ), 
	.A2(n22), 
	.A1(n523));
   AO22CHD U2710 (.O(n1285), 
	.B2(n131), 
	.B1(\ram[43][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n523));
   AO22CHD U2711 (.O(n1286), 
	.B2(n133), 
	.B1(\ram[44][0] ), 
	.A2(n6), 
	.A1(n525));
   AO22CHD U2712 (.O(n1287), 
	.B2(n133), 
	.B1(\ram[44][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n525));
   AO22CHD U2713 (.O(n1288), 
	.B2(n133), 
	.B1(\ram[44][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n525));
   AO22CHD U2714 (.O(n1289), 
	.B2(n133), 
	.B1(\ram[44][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n525));
   AO22CHD U2715 (.O(n1290), 
	.B2(n133), 
	.B1(\ram[44][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n525));
   AO22CHD U2716 (.O(n1291), 
	.B2(n133), 
	.B1(\ram[44][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n525));
   AO22CHD U2717 (.O(n1292), 
	.B2(n133), 
	.B1(\ram[44][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n525));
   AO22CHD U2718 (.O(n1293), 
	.B2(n133), 
	.B1(\ram[44][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n525));
   AO22CHD U2719 (.O(n1294), 
	.B2(n133), 
	.B1(\ram[44][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n525));
   AO22CHD U2720 (.O(n1295), 
	.B2(n133), 
	.B1(\ram[44][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n525));
   AO22CHD U2721 (.O(n1296), 
	.B2(n133), 
	.B1(\ram[44][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n525));
   AO22CHD U2722 (.O(n1297), 
	.B2(n133), 
	.B1(\ram[44][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n525));
   AO22CHD U2723 (.O(n1298), 
	.B2(n133), 
	.B1(\ram[44][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n525));
   AO22CHD U2724 (.O(n1299), 
	.B2(n133), 
	.B1(\ram[44][13] ), 
	.A2(n21), 
	.A1(n525));
   AO22CHD U2725 (.O(n1300), 
	.B2(n133), 
	.B1(\ram[44][14] ), 
	.A2(n22), 
	.A1(n525));
   AO22CHD U2726 (.O(n1301), 
	.B2(n133), 
	.B1(\ram[44][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n525));
   AO22CHD U2727 (.O(n1302), 
	.B2(n135), 
	.B1(FE_PHN2598_ram_45__0_), 
	.A2(n6), 
	.A1(n527));
   AO22CHD U2728 (.O(n1303), 
	.B2(n135), 
	.B1(\ram[45][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n527));
   AO22CHD U2729 (.O(n1304), 
	.B2(n135), 
	.B1(\ram[45][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n527));
   AO22CHD U2730 (.O(n1305), 
	.B2(n135), 
	.B1(\ram[45][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n527));
   AO22CHD U2731 (.O(n1306), 
	.B2(n135), 
	.B1(\ram[45][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n527));
   AO22CHD U2732 (.O(n1307), 
	.B2(n135), 
	.B1(\ram[45][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n527));
   AO22CHD U2733 (.O(n1308), 
	.B2(n135), 
	.B1(\ram[45][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n527));
   AO22CHD U2734 (.O(n1309), 
	.B2(n135), 
	.B1(\ram[45][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n527));
   AO22CHD U2735 (.O(n1310), 
	.B2(n135), 
	.B1(FE_PHN2288_ram_45__8_), 
	.A2(FE_OFN66_n16), 
	.A1(n527));
   AO22CHD U2736 (.O(n1311), 
	.B2(n135), 
	.B1(\ram[45][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n527));
   AO22CHD U2737 (.O(n1312), 
	.B2(n135), 
	.B1(\ram[45][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n527));
   AO22CHD U2738 (.O(n1313), 
	.B2(n135), 
	.B1(FE_PHN2802_ram_45__11_), 
	.A2(FE_OFN76_n19), 
	.A1(n527));
   AO22CHD U2739 (.O(n1314), 
	.B2(n135), 
	.B1(\ram[45][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n527));
   AO22CHD U2740 (.O(n1315), 
	.B2(n135), 
	.B1(\ram[45][13] ), 
	.A2(n21), 
	.A1(n527));
   AO22CHD U2741 (.O(n1316), 
	.B2(n135), 
	.B1(FE_PHN2494_ram_45__14_), 
	.A2(n22), 
	.A1(n527));
   AO22CHD U2742 (.O(n1317), 
	.B2(n135), 
	.B1(\ram[45][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n527));
   AO22CHD U2743 (.O(n1318), 
	.B2(n137), 
	.B1(\ram[46][0] ), 
	.A2(n6), 
	.A1(n529));
   AO22CHD U2744 (.O(n1319), 
	.B2(n137), 
	.B1(\ram[46][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n529));
   AO22CHD U2745 (.O(n1320), 
	.B2(n137), 
	.B1(FE_PHN2979_ram_46__2_), 
	.A2(FE_OFN49_n10), 
	.A1(n529));
   AO22CHD U2746 (.O(n1321), 
	.B2(n137), 
	.B1(\ram[46][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n529));
   AO22CHD U2747 (.O(n1322), 
	.B2(n137), 
	.B1(\ram[46][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n529));
   AO22CHD U2748 (.O(n1323), 
	.B2(n137), 
	.B1(\ram[46][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n529));
   AO22CHD U2749 (.O(n1324), 
	.B2(n137), 
	.B1(\ram[46][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n529));
   AO22CHD U2750 (.O(n1325), 
	.B2(n137), 
	.B1(\ram[46][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n529));
   AO22CHD U2751 (.O(n1326), 
	.B2(n137), 
	.B1(\ram[46][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n529));
   AO22CHD U2752 (.O(n1327), 
	.B2(n137), 
	.B1(\ram[46][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n529));
   AO22CHD U2753 (.O(n1328), 
	.B2(n137), 
	.B1(\ram[46][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n529));
   AO22CHD U2754 (.O(n1329), 
	.B2(n137), 
	.B1(\ram[46][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n529));
   AO22CHD U2755 (.O(n1330), 
	.B2(n137), 
	.B1(\ram[46][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n529));
   AO22CHD U2756 (.O(n1331), 
	.B2(n137), 
	.B1(\ram[46][13] ), 
	.A2(n21), 
	.A1(n529));
   AO22CHD U2757 (.O(n1332), 
	.B2(n137), 
	.B1(\ram[46][14] ), 
	.A2(n22), 
	.A1(n529));
   AO22CHD U2758 (.O(n1333), 
	.B2(n137), 
	.B1(\ram[46][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n529));
   AO22CHD U2759 (.O(n1334), 
	.B2(n139), 
	.B1(\ram[47][0] ), 
	.A2(n6), 
	.A1(n531));
   AO22CHD U2760 (.O(n1335), 
	.B2(n139), 
	.B1(\ram[47][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n531));
   AO22CHD U2761 (.O(n1336), 
	.B2(n139), 
	.B1(\ram[47][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n531));
   AO22CHD U2762 (.O(n1337), 
	.B2(n139), 
	.B1(\ram[47][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n531));
   AO22CHD U2763 (.O(n1338), 
	.B2(n139), 
	.B1(\ram[47][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n531));
   AO22CHD U2764 (.O(n1339), 
	.B2(n139), 
	.B1(\ram[47][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n531));
   AO22CHD U2765 (.O(n1340), 
	.B2(n139), 
	.B1(\ram[47][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n531));
   AO22CHD U2766 (.O(n1341), 
	.B2(n139), 
	.B1(\ram[47][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n531));
   AO22CHD U2767 (.O(n1342), 
	.B2(n139), 
	.B1(\ram[47][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n531));
   AO22CHD U2768 (.O(n1343), 
	.B2(n139), 
	.B1(\ram[47][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n531));
   AO22CHD U2769 (.O(n1344), 
	.B2(n139), 
	.B1(\ram[47][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n531));
   AO22CHD U2770 (.O(n1345), 
	.B2(n139), 
	.B1(\ram[47][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n531));
   AO22CHD U2771 (.O(n1346), 
	.B2(n139), 
	.B1(\ram[47][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n531));
   AO22CHD U2772 (.O(n1347), 
	.B2(n139), 
	.B1(\ram[47][13] ), 
	.A2(n21), 
	.A1(n531));
   AO22CHD U2773 (.O(n1348), 
	.B2(n139), 
	.B1(\ram[47][14] ), 
	.A2(n22), 
	.A1(n531));
   AO22CHD U2774 (.O(n1349), 
	.B2(n139), 
	.B1(\ram[47][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n531));
   AO22CHD U2775 (.O(n1350), 
	.B2(n142), 
	.B1(\ram[48][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n533));
   AO22CHD U2776 (.O(n1351), 
	.B2(n142), 
	.B1(\ram[48][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n533));
   AO22CHD U2777 (.O(n1352), 
	.B2(n142), 
	.B1(\ram[48][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n533));
   AO22CHD U2778 (.O(n1353), 
	.B2(n142), 
	.B1(\ram[48][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n533));
   AO22CHD U2779 (.O(n1354), 
	.B2(n142), 
	.B1(\ram[48][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n533));
   AO22CHD U2780 (.O(n1355), 
	.B2(n142), 
	.B1(\ram[48][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n533));
   AO22CHD U2781 (.O(n1356), 
	.B2(n142), 
	.B1(\ram[48][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n533));
   AO22CHD U2782 (.O(n1357), 
	.B2(n142), 
	.B1(\ram[48][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n533));
   AO22CHD U2783 (.O(n1358), 
	.B2(n142), 
	.B1(\ram[48][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n533));
   AO22CHD U2784 (.O(n1359), 
	.B2(n142), 
	.B1(\ram[48][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n533));
   AO22CHD U2785 (.O(n1360), 
	.B2(n142), 
	.B1(\ram[48][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n533));
   AO22CHD U2786 (.O(n1361), 
	.B2(n142), 
	.B1(\ram[48][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n533));
   AO22CHD U2787 (.O(n1362), 
	.B2(n142), 
	.B1(\ram[48][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n533));
   AO22CHD U2788 (.O(n1363), 
	.B2(n142), 
	.B1(\ram[48][13] ), 
	.A2(n21), 
	.A1(n533));
   AO22CHD U2789 (.O(n1364), 
	.B2(n142), 
	.B1(\ram[48][14] ), 
	.A2(n22), 
	.A1(n533));
   AO22CHD U2790 (.O(n1365), 
	.B2(n142), 
	.B1(\ram[48][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n533));
   AO22CHD U2791 (.O(n1366), 
	.B2(n145), 
	.B1(\ram[49][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n535));
   AO22CHD U2792 (.O(n1367), 
	.B2(n145), 
	.B1(\ram[49][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n535));
   AO22CHD U2793 (.O(n1368), 
	.B2(n145), 
	.B1(\ram[49][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n535));
   AO22CHD U2794 (.O(n1369), 
	.B2(n145), 
	.B1(\ram[49][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n535));
   AO22CHD U2795 (.O(n1370), 
	.B2(n145), 
	.B1(\ram[49][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n535));
   AO22CHD U2796 (.O(n1371), 
	.B2(n145), 
	.B1(\ram[49][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n535));
   AO22CHD U2797 (.O(n1372), 
	.B2(n145), 
	.B1(\ram[49][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n535));
   AO22CHD U2798 (.O(n1373), 
	.B2(n145), 
	.B1(\ram[49][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n535));
   AO22CHD U2799 (.O(n1374), 
	.B2(n145), 
	.B1(\ram[49][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n535));
   AO22CHD U2800 (.O(n1375), 
	.B2(n145), 
	.B1(\ram[49][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n535));
   AO22CHD U2801 (.O(n1376), 
	.B2(n145), 
	.B1(\ram[49][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n535));
   AO22CHD U2802 (.O(n1377), 
	.B2(n145), 
	.B1(\ram[49][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n535));
   AO22CHD U2803 (.O(n1378), 
	.B2(n145), 
	.B1(\ram[49][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n535));
   AO22CHD U2804 (.O(n1379), 
	.B2(n145), 
	.B1(\ram[49][13] ), 
	.A2(n21), 
	.A1(n535));
   AO22CHD U2805 (.O(n1380), 
	.B2(n145), 
	.B1(\ram[49][14] ), 
	.A2(n22), 
	.A1(n535));
   AO22CHD U2806 (.O(n1381), 
	.B2(n145), 
	.B1(\ram[49][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n535));
   AO22CHD U2807 (.O(n1382), 
	.B2(n147), 
	.B1(\ram[50][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n537));
   AO22CHD U2808 (.O(n1383), 
	.B2(n147), 
	.B1(\ram[50][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n537));
   AO22CHD U2809 (.O(n1384), 
	.B2(n147), 
	.B1(\ram[50][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n537));
   AO22CHD U2810 (.O(n1385), 
	.B2(n147), 
	.B1(\ram[50][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n537));
   AO22CHD U2811 (.O(n1386), 
	.B2(n147), 
	.B1(\ram[50][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n537));
   AO22CHD U2812 (.O(n1387), 
	.B2(n147), 
	.B1(\ram[50][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n537));
   AO22CHD U2813 (.O(n1388), 
	.B2(n147), 
	.B1(\ram[50][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n537));
   AO22CHD U2814 (.O(n1389), 
	.B2(n147), 
	.B1(\ram[50][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n537));
   AO22CHD U2815 (.O(n1390), 
	.B2(n147), 
	.B1(\ram[50][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n537));
   AO22CHD U2816 (.O(n1391), 
	.B2(n147), 
	.B1(\ram[50][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n537));
   AO22CHD U2817 (.O(n1392), 
	.B2(n147), 
	.B1(\ram[50][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n537));
   AO22CHD U2818 (.O(n1393), 
	.B2(n147), 
	.B1(\ram[50][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n537));
   AO22CHD U2819 (.O(n1394), 
	.B2(n147), 
	.B1(\ram[50][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n537));
   AO22CHD U2820 (.O(n1395), 
	.B2(n147), 
	.B1(\ram[50][13] ), 
	.A2(n21), 
	.A1(n537));
   AO22CHD U2821 (.O(n1396), 
	.B2(n147), 
	.B1(\ram[50][14] ), 
	.A2(n22), 
	.A1(n537));
   AO22CHD U2822 (.O(n1397), 
	.B2(n147), 
	.B1(\ram[50][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n537));
   AO22CHD U2823 (.O(n1398), 
	.B2(n149), 
	.B1(\ram[51][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n539));
   AO22CHD U2824 (.O(n1399), 
	.B2(n149), 
	.B1(\ram[51][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n539));
   AO22CHD U2825 (.O(n1400), 
	.B2(n149), 
	.B1(\ram[51][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n539));
   AO22CHD U2826 (.O(n1401), 
	.B2(n149), 
	.B1(\ram[51][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n539));
   AO22CHD U2827 (.O(n1402), 
	.B2(n149), 
	.B1(\ram[51][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n539));
   AO22CHD U2828 (.O(n1403), 
	.B2(n149), 
	.B1(\ram[51][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n539));
   AO22CHD U2829 (.O(n1404), 
	.B2(n149), 
	.B1(\ram[51][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n539));
   AO22CHD U2830 (.O(n1405), 
	.B2(n149), 
	.B1(\ram[51][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n539));
   AO22CHD U2831 (.O(n1406), 
	.B2(n149), 
	.B1(\ram[51][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n539));
   AO22CHD U2832 (.O(n1407), 
	.B2(n149), 
	.B1(\ram[51][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n539));
   AO22CHD U2833 (.O(n1408), 
	.B2(n149), 
	.B1(\ram[51][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n539));
   AO22CHD U2834 (.O(n1409), 
	.B2(n149), 
	.B1(\ram[51][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n539));
   AO22CHD U2835 (.O(n1410), 
	.B2(n149), 
	.B1(\ram[51][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n539));
   AO22CHD U2836 (.O(n1411), 
	.B2(n149), 
	.B1(\ram[51][13] ), 
	.A2(n21), 
	.A1(n539));
   AO22CHD U2837 (.O(n1412), 
	.B2(n149), 
	.B1(\ram[51][14] ), 
	.A2(n22), 
	.A1(n539));
   AO22CHD U2838 (.O(n1413), 
	.B2(n149), 
	.B1(\ram[51][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n539));
   AO22CHD U2839 (.O(n1414), 
	.B2(n151), 
	.B1(\ram[52][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n541));
   AO22CHD U2840 (.O(n1415), 
	.B2(n151), 
	.B1(\ram[52][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n541));
   AO22CHD U2841 (.O(n1416), 
	.B2(n151), 
	.B1(\ram[52][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n541));
   AO22CHD U2842 (.O(n1417), 
	.B2(n151), 
	.B1(\ram[52][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n541));
   AO22CHD U2843 (.O(n1418), 
	.B2(n151), 
	.B1(\ram[52][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n541));
   AO22CHD U2844 (.O(n1419), 
	.B2(n151), 
	.B1(\ram[52][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n541));
   AO22CHD U2845 (.O(n1420), 
	.B2(n151), 
	.B1(\ram[52][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n541));
   AO22CHD U2846 (.O(n1421), 
	.B2(n151), 
	.B1(\ram[52][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n541));
   AO22CHD U2847 (.O(n1422), 
	.B2(n151), 
	.B1(\ram[52][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n541));
   AO22CHD U2848 (.O(n1423), 
	.B2(n151), 
	.B1(\ram[52][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n541));
   AO22CHD U2849 (.O(n1424), 
	.B2(n151), 
	.B1(\ram[52][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n541));
   AO22CHD U2850 (.O(n1425), 
	.B2(n151), 
	.B1(\ram[52][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n541));
   AO22CHD U2851 (.O(n1426), 
	.B2(n151), 
	.B1(\ram[52][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n541));
   AO22CHD U2852 (.O(n1427), 
	.B2(n151), 
	.B1(\ram[52][13] ), 
	.A2(n21), 
	.A1(n541));
   AO22CHD U2853 (.O(n1428), 
	.B2(n151), 
	.B1(\ram[52][14] ), 
	.A2(n22), 
	.A1(n541));
   AO22CHD U2854 (.O(n1429), 
	.B2(n151), 
	.B1(FE_PHN3073_ram_52__15_), 
	.A2(FE_OFN89_n23), 
	.A1(n541));
   AO22CHD U2855 (.O(n1430), 
	.B2(n153), 
	.B1(\ram[53][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n543));
   AO22CHD U2856 (.O(n1431), 
	.B2(n153), 
	.B1(\ram[53][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n543));
   AO22CHD U2857 (.O(n1432), 
	.B2(n153), 
	.B1(\ram[53][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n543));
   AO22CHD U2858 (.O(n1433), 
	.B2(n153), 
	.B1(\ram[53][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n543));
   AO22CHD U2859 (.O(n1434), 
	.B2(n153), 
	.B1(\ram[53][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n543));
   AO22CHD U2860 (.O(n1435), 
	.B2(n153), 
	.B1(\ram[53][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n543));
   AO22CHD U2861 (.O(n1436), 
	.B2(n153), 
	.B1(\ram[53][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n543));
   AO22CHD U2862 (.O(n1437), 
	.B2(n153), 
	.B1(\ram[53][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n543));
   AO22CHD U2863 (.O(n1438), 
	.B2(n153), 
	.B1(\ram[53][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n543));
   AO22CHD U2864 (.O(n1439), 
	.B2(n153), 
	.B1(\ram[53][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n543));
   AO22CHD U2865 (.O(n1440), 
	.B2(n153), 
	.B1(\ram[53][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n543));
   AO22CHD U2866 (.O(n1441), 
	.B2(n153), 
	.B1(\ram[53][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n543));
   AO22CHD U2867 (.O(n1442), 
	.B2(n153), 
	.B1(\ram[53][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n543));
   AO22CHD U2868 (.O(n1443), 
	.B2(n153), 
	.B1(\ram[53][13] ), 
	.A2(n21), 
	.A1(n543));
   AO22CHD U2869 (.O(n1444), 
	.B2(n153), 
	.B1(\ram[53][14] ), 
	.A2(n22), 
	.A1(n543));
   AO22CHD U2870 (.O(n1445), 
	.B2(n153), 
	.B1(\ram[53][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n543));
   AO22CHD U2871 (.O(n1446), 
	.B2(n155), 
	.B1(\ram[54][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n546));
   AO22CHD U2872 (.O(n1447), 
	.B2(n155), 
	.B1(\ram[54][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n546));
   AO22CHD U2873 (.O(n1448), 
	.B2(n155), 
	.B1(\ram[54][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n546));
   AO22CHD U2874 (.O(n1449), 
	.B2(n155), 
	.B1(\ram[54][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n546));
   AO22CHD U2875 (.O(n1450), 
	.B2(n155), 
	.B1(\ram[54][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n546));
   AO22CHD U2876 (.O(n1451), 
	.B2(n155), 
	.B1(\ram[54][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n546));
   AO22CHD U2877 (.O(n1452), 
	.B2(n155), 
	.B1(\ram[54][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n546));
   AO22CHD U2878 (.O(n1453), 
	.B2(n155), 
	.B1(\ram[54][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n546));
   AO22CHD U2879 (.O(n1454), 
	.B2(n155), 
	.B1(\ram[54][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n546));
   AO22CHD U2880 (.O(n1455), 
	.B2(n155), 
	.B1(\ram[54][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n546));
   AO22CHD U2881 (.O(n1456), 
	.B2(n155), 
	.B1(\ram[54][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n546));
   AO22CHD U2882 (.O(n1457), 
	.B2(n155), 
	.B1(\ram[54][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n546));
   AO22CHD U2883 (.O(n1458), 
	.B2(n155), 
	.B1(\ram[54][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n546));
   AO22CHD U2884 (.O(n1459), 
	.B2(n155), 
	.B1(\ram[54][13] ), 
	.A2(n21), 
	.A1(n546));
   AO22CHD U2885 (.O(n1460), 
	.B2(n155), 
	.B1(\ram[54][14] ), 
	.A2(n22), 
	.A1(n546));
   AO22CHD U2886 (.O(n1461), 
	.B2(n155), 
	.B1(\ram[54][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n546));
   AO22CHD U2887 (.O(n1462), 
	.B2(n157), 
	.B1(\ram[55][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n549));
   AO22CHD U2888 (.O(n1463), 
	.B2(n157), 
	.B1(\ram[55][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n549));
   AO22CHD U2889 (.O(n1464), 
	.B2(n157), 
	.B1(\ram[55][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n549));
   AO22CHD U2890 (.O(n1465), 
	.B2(n157), 
	.B1(\ram[55][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n549));
   AO22CHD U2891 (.O(n1466), 
	.B2(n157), 
	.B1(\ram[55][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n549));
   AO22CHD U2892 (.O(n1467), 
	.B2(n157), 
	.B1(\ram[55][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n549));
   AO22CHD U2893 (.O(n1468), 
	.B2(n157), 
	.B1(\ram[55][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n549));
   AO22CHD U2894 (.O(n1469), 
	.B2(n157), 
	.B1(\ram[55][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n549));
   AO22CHD U2895 (.O(n1470), 
	.B2(n157), 
	.B1(\ram[55][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n549));
   AO22CHD U2896 (.O(n1471), 
	.B2(n157), 
	.B1(\ram[55][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n549));
   AO22CHD U2897 (.O(n1472), 
	.B2(n157), 
	.B1(\ram[55][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n549));
   AO22CHD U2898 (.O(n1473), 
	.B2(n157), 
	.B1(\ram[55][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n549));
   AO22CHD U2899 (.O(n1474), 
	.B2(n157), 
	.B1(\ram[55][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n549));
   AO22CHD U2900 (.O(n1475), 
	.B2(n157), 
	.B1(\ram[55][13] ), 
	.A2(n21), 
	.A1(n549));
   AO22CHD U2901 (.O(n1476), 
	.B2(n157), 
	.B1(\ram[55][14] ), 
	.A2(n22), 
	.A1(n549));
   AO22CHD U2902 (.O(n1477), 
	.B2(n157), 
	.B1(\ram[55][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n549));
   AO22CHD U2903 (.O(n1478), 
	.B2(n159), 
	.B1(\ram[56][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n552));
   AO22CHD U2904 (.O(n1479), 
	.B2(n159), 
	.B1(\ram[56][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n552));
   AO22CHD U2905 (.O(n1480), 
	.B2(n159), 
	.B1(\ram[56][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n552));
   AO22CHD U2906 (.O(n1481), 
	.B2(n159), 
	.B1(\ram[56][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n552));
   AO22CHD U2907 (.O(n1482), 
	.B2(n159), 
	.B1(\ram[56][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n552));
   AO22CHD U2908 (.O(n1483), 
	.B2(n159), 
	.B1(\ram[56][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n552));
   AO22CHD U2909 (.O(n1484), 
	.B2(n159), 
	.B1(\ram[56][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n552));
   AO22CHD U2910 (.O(n1485), 
	.B2(n159), 
	.B1(\ram[56][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n552));
   AO22CHD U2911 (.O(n1486), 
	.B2(n159), 
	.B1(\ram[56][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n552));
   AO22CHD U2912 (.O(n1487), 
	.B2(n159), 
	.B1(\ram[56][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n552));
   AO22CHD U2913 (.O(n1488), 
	.B2(n159), 
	.B1(\ram[56][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n552));
   AO22CHD U2914 (.O(n1489), 
	.B2(n159), 
	.B1(\ram[56][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n552));
   AO22CHD U2915 (.O(n1490), 
	.B2(n159), 
	.B1(\ram[56][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n552));
   AO22CHD U2916 (.O(n1491), 
	.B2(n159), 
	.B1(\ram[56][13] ), 
	.A2(n21), 
	.A1(n552));
   AO22CHD U2917 (.O(n1492), 
	.B2(n159), 
	.B1(\ram[56][14] ), 
	.A2(n22), 
	.A1(n552));
   AO22CHD U2918 (.O(n1493), 
	.B2(n159), 
	.B1(\ram[56][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n552));
   AO22CHD U2919 (.O(n1494), 
	.B2(n161), 
	.B1(\ram[57][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n555));
   AO22CHD U2920 (.O(n1495), 
	.B2(n161), 
	.B1(\ram[57][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n555));
   AO22CHD U2921 (.O(n1496), 
	.B2(n161), 
	.B1(\ram[57][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n555));
   AO22CHD U2922 (.O(n1497), 
	.B2(n161), 
	.B1(\ram[57][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n555));
   AO22CHD U2923 (.O(n1498), 
	.B2(n161), 
	.B1(\ram[57][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n555));
   AO22CHD U2924 (.O(n1499), 
	.B2(n161), 
	.B1(\ram[57][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n555));
   AO22CHD U2925 (.O(n1500), 
	.B2(n161), 
	.B1(\ram[57][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n555));
   AO22CHD U2926 (.O(n1501), 
	.B2(n161), 
	.B1(\ram[57][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n555));
   AO22CHD U2927 (.O(n1502), 
	.B2(n161), 
	.B1(\ram[57][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n555));
   AO22CHD U2928 (.O(n1503), 
	.B2(n161), 
	.B1(\ram[57][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n555));
   AO22CHD U2929 (.O(n1504), 
	.B2(n161), 
	.B1(\ram[57][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n555));
   AO22CHD U2930 (.O(n1505), 
	.B2(n161), 
	.B1(\ram[57][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n555));
   AO22CHD U2931 (.O(n1506), 
	.B2(n161), 
	.B1(\ram[57][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n555));
   AO22CHD U2932 (.O(n1507), 
	.B2(n161), 
	.B1(\ram[57][13] ), 
	.A2(n21), 
	.A1(n555));
   AO22CHD U2933 (.O(n1508), 
	.B2(n161), 
	.B1(\ram[57][14] ), 
	.A2(n22), 
	.A1(n555));
   AO22CHD U2934 (.O(n1509), 
	.B2(n161), 
	.B1(\ram[57][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n555));
   AO22CHD U2935 (.O(n1510), 
	.B2(n163), 
	.B1(\ram[58][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n558));
   AO22CHD U2936 (.O(n1511), 
	.B2(n163), 
	.B1(\ram[58][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n558));
   AO22CHD U2937 (.O(n1512), 
	.B2(n163), 
	.B1(\ram[58][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n558));
   AO22CHD U2938 (.O(n1513), 
	.B2(n163), 
	.B1(\ram[58][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n558));
   AO22CHD U2939 (.O(n1514), 
	.B2(n163), 
	.B1(\ram[58][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n558));
   AO22CHD U2940 (.O(n1515), 
	.B2(n163), 
	.B1(\ram[58][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n558));
   AO22CHD U2941 (.O(n1516), 
	.B2(n163), 
	.B1(\ram[58][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n558));
   AO22CHD U2942 (.O(n1517), 
	.B2(n163), 
	.B1(\ram[58][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n558));
   AO22CHD U2943 (.O(n1518), 
	.B2(n163), 
	.B1(\ram[58][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n558));
   AO22CHD U2944 (.O(n1519), 
	.B2(n163), 
	.B1(\ram[58][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n558));
   AO22CHD U2945 (.O(n1520), 
	.B2(n163), 
	.B1(\ram[58][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n558));
   AO22CHD U2946 (.O(n1521), 
	.B2(n163), 
	.B1(\ram[58][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n558));
   AO22CHD U2947 (.O(n1522), 
	.B2(n163), 
	.B1(\ram[58][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n558));
   AO22CHD U2948 (.O(n1523), 
	.B2(n163), 
	.B1(\ram[58][13] ), 
	.A2(n21), 
	.A1(n558));
   AO22CHD U2949 (.O(n1524), 
	.B2(n163), 
	.B1(\ram[58][14] ), 
	.A2(n22), 
	.A1(n558));
   AO22CHD U2950 (.O(n1525), 
	.B2(n163), 
	.B1(\ram[58][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n558));
   AO22CHD U2951 (.O(n1526), 
	.B2(n165), 
	.B1(\ram[59][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n560));
   AO22CHD U2952 (.O(n1527), 
	.B2(n165), 
	.B1(\ram[59][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n560));
   AO22CHD U2953 (.O(n1528), 
	.B2(n165), 
	.B1(\ram[59][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n560));
   AO22CHD U2954 (.O(n1529), 
	.B2(n165), 
	.B1(\ram[59][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n560));
   AO22CHD U2955 (.O(n1530), 
	.B2(n165), 
	.B1(\ram[59][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n560));
   AO22CHD U2956 (.O(n1531), 
	.B2(n165), 
	.B1(\ram[59][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n560));
   AO22CHD U2957 (.O(n1532), 
	.B2(n165), 
	.B1(\ram[59][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n560));
   AO22CHD U2958 (.O(n1533), 
	.B2(n165), 
	.B1(\ram[59][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n560));
   AO22CHD U2959 (.O(n1534), 
	.B2(n165), 
	.B1(\ram[59][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n560));
   AO22CHD U2960 (.O(n1535), 
	.B2(n165), 
	.B1(\ram[59][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n560));
   AO22CHD U2961 (.O(n1536), 
	.B2(n165), 
	.B1(\ram[59][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n560));
   AO22CHD U2962 (.O(n1537), 
	.B2(n165), 
	.B1(\ram[59][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n560));
   AO22CHD U2963 (.O(n1538), 
	.B2(n165), 
	.B1(\ram[59][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n560));
   AO22CHD U2964 (.O(n1539), 
	.B2(n165), 
	.B1(\ram[59][13] ), 
	.A2(n21), 
	.A1(n560));
   AO22CHD U2965 (.O(n1540), 
	.B2(n165), 
	.B1(\ram[59][14] ), 
	.A2(n22), 
	.A1(n560));
   AO22CHD U2966 (.O(n1541), 
	.B2(n165), 
	.B1(\ram[59][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n560));
   AO22CHD U2967 (.O(n1542), 
	.B2(n167), 
	.B1(\ram[60][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n562));
   AO22CHD U2968 (.O(n1543), 
	.B2(n167), 
	.B1(\ram[60][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n562));
   AO22CHD U2969 (.O(n1544), 
	.B2(n167), 
	.B1(\ram[60][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n562));
   AO22CHD U2970 (.O(n1545), 
	.B2(n167), 
	.B1(\ram[60][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n562));
   AO22CHD U2971 (.O(n1546), 
	.B2(n167), 
	.B1(\ram[60][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n562));
   AO22CHD U2972 (.O(n1547), 
	.B2(n167), 
	.B1(\ram[60][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n562));
   AO22CHD U2973 (.O(n1548), 
	.B2(n167), 
	.B1(\ram[60][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n562));
   AO22CHD U2974 (.O(n1549), 
	.B2(n167), 
	.B1(\ram[60][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n562));
   AO22CHD U2975 (.O(n1550), 
	.B2(n167), 
	.B1(\ram[60][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n562));
   AO22CHD U2976 (.O(n1551), 
	.B2(n167), 
	.B1(\ram[60][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n562));
   AO22CHD U2977 (.O(n1552), 
	.B2(n167), 
	.B1(\ram[60][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n562));
   AO22CHD U2978 (.O(n1553), 
	.B2(n167), 
	.B1(\ram[60][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n562));
   AO22CHD U2979 (.O(n1554), 
	.B2(n167), 
	.B1(\ram[60][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n562));
   AO22CHD U2980 (.O(n1555), 
	.B2(n167), 
	.B1(\ram[60][13] ), 
	.A2(n21), 
	.A1(n562));
   AO22CHD U2981 (.O(n1556), 
	.B2(n167), 
	.B1(\ram[60][14] ), 
	.A2(n22), 
	.A1(n562));
   AO22CHD U2982 (.O(n1557), 
	.B2(n167), 
	.B1(\ram[60][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n562));
   AO22CHD U2983 (.O(n1558), 
	.B2(n169), 
	.B1(\ram[61][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n564));
   AO22CHD U2984 (.O(n1559), 
	.B2(n169), 
	.B1(\ram[61][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n564));
   AO22CHD U2985 (.O(n1560), 
	.B2(n169), 
	.B1(\ram[61][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n564));
   AO22CHD U2986 (.O(n1561), 
	.B2(n169), 
	.B1(\ram[61][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n564));
   AO22CHD U2987 (.O(n1562), 
	.B2(n169), 
	.B1(\ram[61][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n564));
   AO22CHD U2988 (.O(n1563), 
	.B2(n169), 
	.B1(\ram[61][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n564));
   AO22CHD U2989 (.O(n1564), 
	.B2(n169), 
	.B1(\ram[61][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n564));
   AO22CHD U2990 (.O(n1565), 
	.B2(n169), 
	.B1(\ram[61][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n564));
   AO22CHD U2991 (.O(n1566), 
	.B2(n169), 
	.B1(\ram[61][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n564));
   AO22CHD U2992 (.O(n1567), 
	.B2(n169), 
	.B1(\ram[61][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n564));
   AO22CHD U2993 (.O(n1568), 
	.B2(n169), 
	.B1(\ram[61][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n564));
   AO22CHD U2994 (.O(n1569), 
	.B2(n169), 
	.B1(\ram[61][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n564));
   AO22CHD U2995 (.O(n1570), 
	.B2(n169), 
	.B1(\ram[61][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n564));
   AO22CHD U2996 (.O(n1571), 
	.B2(n169), 
	.B1(FE_PHN1778_ram_61__13_), 
	.A2(n21), 
	.A1(n564));
   AO22CHD U2997 (.O(n1572), 
	.B2(n169), 
	.B1(\ram[61][14] ), 
	.A2(n22), 
	.A1(n564));
   AO22CHD U2998 (.O(n1573), 
	.B2(n169), 
	.B1(\ram[61][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n564));
   AO22CHD U2999 (.O(n1574), 
	.B2(n171), 
	.B1(\ram[62][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n567));
   AO22CHD U3000 (.O(n1575), 
	.B2(n171), 
	.B1(\ram[62][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n567));
   AO22CHD U3001 (.O(n1576), 
	.B2(n171), 
	.B1(\ram[62][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n567));
   AO22CHD U3002 (.O(n1577), 
	.B2(n171), 
	.B1(\ram[62][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n567));
   AO22CHD U3003 (.O(n1578), 
	.B2(n171), 
	.B1(\ram[62][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n567));
   AO22CHD U3004 (.O(n1579), 
	.B2(n171), 
	.B1(\ram[62][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n567));
   AO22CHD U3005 (.O(n1580), 
	.B2(n171), 
	.B1(\ram[62][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n567));
   AO22CHD U3006 (.O(n1581), 
	.B2(n171), 
	.B1(\ram[62][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n567));
   AO22CHD U3007 (.O(n1582), 
	.B2(n171), 
	.B1(\ram[62][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n567));
   AO22CHD U3008 (.O(n1583), 
	.B2(n171), 
	.B1(\ram[62][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n567));
   AO22CHD U3009 (.O(n1584), 
	.B2(n171), 
	.B1(\ram[62][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n567));
   AO22CHD U3010 (.O(n1585), 
	.B2(n171), 
	.B1(\ram[62][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n567));
   AO22CHD U3011 (.O(n1586), 
	.B2(n171), 
	.B1(\ram[62][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n567));
   AO22CHD U3012 (.O(n1587), 
	.B2(n171), 
	.B1(\ram[62][13] ), 
	.A2(n21), 
	.A1(n567));
   AO22CHD U3013 (.O(n1588), 
	.B2(n171), 
	.B1(\ram[62][14] ), 
	.A2(n22), 
	.A1(n567));
   AO22CHD U3014 (.O(n1589), 
	.B2(n171), 
	.B1(\ram[62][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n567));
   AO22CHD U3015 (.O(n1590), 
	.B2(n173), 
	.B1(\ram[63][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n569));
   AO22CHD U3016 (.O(n1591), 
	.B2(n173), 
	.B1(\ram[63][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n569));
   AO22CHD U3017 (.O(n1592), 
	.B2(n173), 
	.B1(\ram[63][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n569));
   AO22CHD U3018 (.O(n1593), 
	.B2(n173), 
	.B1(\ram[63][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n569));
   AO22CHD U3019 (.O(n1594), 
	.B2(n173), 
	.B1(\ram[63][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n569));
   AO22CHD U3020 (.O(n1595), 
	.B2(n173), 
	.B1(FE_PHN1781_ram_63__5_), 
	.A2(FE_OFN58_n13), 
	.A1(n569));
   AO22CHD U3021 (.O(n1596), 
	.B2(n173), 
	.B1(\ram[63][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n569));
   AO22CHD U3022 (.O(n1597), 
	.B2(n173), 
	.B1(\ram[63][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n569));
   AO22CHD U3023 (.O(n1598), 
	.B2(n173), 
	.B1(\ram[63][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n569));
   AO22CHD U3024 (.O(n1599), 
	.B2(n173), 
	.B1(\ram[63][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n569));
   AO22CHD U3025 (.O(n1600), 
	.B2(n173), 
	.B1(\ram[63][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n569));
   AO22CHD U3026 (.O(n1601), 
	.B2(n173), 
	.B1(\ram[63][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n569));
   AO22CHD U3027 (.O(n1602), 
	.B2(n173), 
	.B1(\ram[63][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n569));
   AO22CHD U3028 (.O(n1603), 
	.B2(n173), 
	.B1(\ram[63][13] ), 
	.A2(n21), 
	.A1(n569));
   AO22CHD U3029 (.O(n1604), 
	.B2(n173), 
	.B1(\ram[63][14] ), 
	.A2(n22), 
	.A1(n569));
   AO22CHD U3030 (.O(n1605), 
	.B2(n173), 
	.B1(\ram[63][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n569));
   AO22CHD U3031 (.O(n1606), 
	.B2(n176), 
	.B1(\ram[64][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n56));
   AO22CHD U3032 (.O(n1607), 
	.B2(n176), 
	.B1(\ram[64][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n56));
   AO22CHD U3033 (.O(n1608), 
	.B2(n176), 
	.B1(\ram[64][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n56));
   AO22CHD U3034 (.O(n1609), 
	.B2(n176), 
	.B1(\ram[64][3] ), 
	.A2(n11), 
	.A1(n56));
   AO22CHD U3035 (.O(n1610), 
	.B2(n176), 
	.B1(\ram[64][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n56));
   AO22CHD U3036 (.O(n1611), 
	.B2(n176), 
	.B1(\ram[64][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n56));
   AO22CHD U3037 (.O(n1612), 
	.B2(n176), 
	.B1(\ram[64][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n56));
   AO22CHD U3038 (.O(n1613), 
	.B2(n176), 
	.B1(\ram[64][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n56));
   AO22CHD U3039 (.O(n1614), 
	.B2(n176), 
	.B1(\ram[64][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n56));
   AO22CHD U3040 (.O(n1615), 
	.B2(n176), 
	.B1(\ram[64][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n56));
   AO22CHD U3041 (.O(n1616), 
	.B2(n176), 
	.B1(\ram[64][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n56));
   AO22CHD U3042 (.O(n1617), 
	.B2(n176), 
	.B1(\ram[64][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n56));
   AO22CHD U3043 (.O(n1618), 
	.B2(n176), 
	.B1(\ram[64][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n56));
   AO22CHD U3044 (.O(n1619), 
	.B2(n176), 
	.B1(\ram[64][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n56));
   AO22CHD U3045 (.O(n1620), 
	.B2(n176), 
	.B1(\ram[64][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n56));
   AO22CHD U3046 (.O(n1621), 
	.B2(n176), 
	.B1(\ram[64][15] ), 
	.A2(n23), 
	.A1(n56));
   AO22CHD U3047 (.O(n1622), 
	.B2(n179), 
	.B1(\ram[65][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n58));
   AO22CHD U3048 (.O(n1623), 
	.B2(n179), 
	.B1(\ram[65][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n58));
   AO22CHD U3049 (.O(n1624), 
	.B2(n179), 
	.B1(\ram[65][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n58));
   AO22CHD U3050 (.O(n1625), 
	.B2(n179), 
	.B1(\ram[65][3] ), 
	.A2(n11), 
	.A1(n58));
   AO22CHD U3051 (.O(n1626), 
	.B2(n179), 
	.B1(\ram[65][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n58));
   AO22CHD U3052 (.O(n1627), 
	.B2(n179), 
	.B1(\ram[65][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n58));
   AO22CHD U3053 (.O(n1628), 
	.B2(n179), 
	.B1(\ram[65][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n58));
   AO22CHD U3054 (.O(n1629), 
	.B2(n179), 
	.B1(\ram[65][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n58));
   AO22CHD U3055 (.O(n1630), 
	.B2(n179), 
	.B1(FE_PHN1321_ram_65__8_), 
	.A2(FE_OFN67_n16), 
	.A1(n58));
   AO22CHD U3056 (.O(n1631), 
	.B2(n179), 
	.B1(\ram[65][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n58));
   AO22CHD U3057 (.O(n1632), 
	.B2(n179), 
	.B1(\ram[65][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n58));
   AO22CHD U3058 (.O(n1633), 
	.B2(n179), 
	.B1(\ram[65][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n58));
   AO22CHD U3059 (.O(n1634), 
	.B2(n179), 
	.B1(\ram[65][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n58));
   AO22CHD U3060 (.O(n1635), 
	.B2(n179), 
	.B1(\ram[65][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n58));
   AO22CHD U3061 (.O(n1636), 
	.B2(n179), 
	.B1(\ram[65][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n58));
   AO22CHD U3062 (.O(n1637), 
	.B2(n179), 
	.B1(\ram[65][15] ), 
	.A2(n23), 
	.A1(n58));
   AO22CHD U3063 (.O(n1638), 
	.B2(n181), 
	.B1(\ram[66][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n59));
   AO22CHD U3064 (.O(n1639), 
	.B2(n181), 
	.B1(\ram[66][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n59));
   AO22CHD U3065 (.O(n1640), 
	.B2(n181), 
	.B1(\ram[66][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n59));
   AO22CHD U3066 (.O(n1641), 
	.B2(n181), 
	.B1(\ram[66][3] ), 
	.A2(n11), 
	.A1(n59));
   AO22CHD U3067 (.O(n1642), 
	.B2(n181), 
	.B1(\ram[66][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n59));
   AO22CHD U3068 (.O(n1643), 
	.B2(n181), 
	.B1(\ram[66][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n59));
   AO22CHD U3069 (.O(n1644), 
	.B2(n181), 
	.B1(\ram[66][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n59));
   AO22CHD U3070 (.O(n1645), 
	.B2(n181), 
	.B1(\ram[66][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n59));
   AO22CHD U3071 (.O(n1646), 
	.B2(n181), 
	.B1(\ram[66][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n59));
   AO22CHD U3072 (.O(n1647), 
	.B2(n181), 
	.B1(\ram[66][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n59));
   AO22CHD U3073 (.O(n1648), 
	.B2(n181), 
	.B1(\ram[66][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n59));
   AO22CHD U3074 (.O(n1649), 
	.B2(n181), 
	.B1(\ram[66][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n59));
   AO22CHD U3075 (.O(n1650), 
	.B2(n181), 
	.B1(\ram[66][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n59));
   AO22CHD U3076 (.O(n1651), 
	.B2(n181), 
	.B1(\ram[66][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n59));
   AO22CHD U3077 (.O(n1652), 
	.B2(n181), 
	.B1(\ram[66][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n59));
   AO22CHD U3078 (.O(n1653), 
	.B2(n181), 
	.B1(\ram[66][15] ), 
	.A2(n23), 
	.A1(n59));
   AO22CHD U3079 (.O(n1654), 
	.B2(n183), 
	.B1(\ram[67][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n61));
   AO22CHD U3080 (.O(n1655), 
	.B2(n183), 
	.B1(\ram[67][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n61));
   AO22CHD U3081 (.O(n1656), 
	.B2(n183), 
	.B1(\ram[67][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n61));
   AO22CHD U3082 (.O(n1657), 
	.B2(n183), 
	.B1(\ram[67][3] ), 
	.A2(n11), 
	.A1(n61));
   AO22CHD U3083 (.O(n1658), 
	.B2(n183), 
	.B1(\ram[67][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n61));
   AO22CHD U3084 (.O(n1659), 
	.B2(n183), 
	.B1(\ram[67][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n61));
   AO22CHD U3085 (.O(n1660), 
	.B2(n183), 
	.B1(\ram[67][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n61));
   AO22CHD U3086 (.O(n1661), 
	.B2(n183), 
	.B1(\ram[67][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n61));
   AO22CHD U3087 (.O(n1662), 
	.B2(n183), 
	.B1(\ram[67][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n61));
   AO22CHD U3088 (.O(n1663), 
	.B2(n183), 
	.B1(FE_PHN2326_ram_67__9_), 
	.A2(FE_OFN71_n17), 
	.A1(n61));
   AO22CHD U3089 (.O(n1664), 
	.B2(n183), 
	.B1(\ram[67][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n61));
   AO22CHD U3090 (.O(n1665), 
	.B2(n183), 
	.B1(\ram[67][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n61));
   AO22CHD U3091 (.O(n1666), 
	.B2(n183), 
	.B1(\ram[67][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n61));
   AO22CHD U3092 (.O(n1667), 
	.B2(n183), 
	.B1(\ram[67][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n61));
   AO22CHD U3093 (.O(n1668), 
	.B2(n183), 
	.B1(\ram[67][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n61));
   AO22CHD U3094 (.O(n1669), 
	.B2(n183), 
	.B1(\ram[67][15] ), 
	.A2(n23), 
	.A1(n61));
   AO22CHD U3095 (.O(n1670), 
	.B2(n185), 
	.B1(\ram[68][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n62));
   AO22CHD U3096 (.O(n1671), 
	.B2(n185), 
	.B1(\ram[68][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n62));
   AO22CHD U3097 (.O(n1672), 
	.B2(n185), 
	.B1(\ram[68][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n62));
   AO22CHD U3098 (.O(n1673), 
	.B2(n185), 
	.B1(\ram[68][3] ), 
	.A2(n11), 
	.A1(n62));
   AO22CHD U3099 (.O(n1674), 
	.B2(n185), 
	.B1(\ram[68][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n62));
   AO22CHD U3100 (.O(n1675), 
	.B2(n185), 
	.B1(\ram[68][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n62));
   AO22CHD U3101 (.O(n1676), 
	.B2(n185), 
	.B1(\ram[68][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n62));
   AO22CHD U3102 (.O(n1677), 
	.B2(n185), 
	.B1(\ram[68][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n62));
   AO22CHD U3103 (.O(n1678), 
	.B2(n185), 
	.B1(\ram[68][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n62));
   AO22CHD U3104 (.O(n1679), 
	.B2(n185), 
	.B1(\ram[68][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n62));
   AO22CHD U3105 (.O(n1680), 
	.B2(n185), 
	.B1(\ram[68][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n62));
   AO22CHD U3106 (.O(n1681), 
	.B2(n185), 
	.B1(\ram[68][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n62));
   AO22CHD U3107 (.O(n1682), 
	.B2(n185), 
	.B1(\ram[68][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n62));
   AO22CHD U3108 (.O(n1683), 
	.B2(n185), 
	.B1(\ram[68][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n62));
   AO22CHD U3109 (.O(n1684), 
	.B2(n185), 
	.B1(\ram[68][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n62));
   AO22CHD U3110 (.O(n1685), 
	.B2(n185), 
	.B1(\ram[68][15] ), 
	.A2(n23), 
	.A1(n62));
   AO22CHD U3111 (.O(n1686), 
	.B2(n187), 
	.B1(\ram[69][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n64));
   AO22CHD U3112 (.O(n1687), 
	.B2(n187), 
	.B1(\ram[69][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n64));
   AO22CHD U3113 (.O(n1688), 
	.B2(n187), 
	.B1(\ram[69][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n64));
   AO22CHD U3114 (.O(n1689), 
	.B2(n187), 
	.B1(\ram[69][3] ), 
	.A2(n11), 
	.A1(n64));
   AO22CHD U3115 (.O(n1690), 
	.B2(n187), 
	.B1(\ram[69][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n64));
   AO22CHD U3116 (.O(n1691), 
	.B2(n187), 
	.B1(\ram[69][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n64));
   AO22CHD U3117 (.O(n1692), 
	.B2(n187), 
	.B1(\ram[69][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n64));
   AO22CHD U3118 (.O(n1693), 
	.B2(n187), 
	.B1(\ram[69][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n64));
   AO22CHD U3119 (.O(n1694), 
	.B2(n187), 
	.B1(\ram[69][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n64));
   AO22CHD U3120 (.O(n1695), 
	.B2(n187), 
	.B1(\ram[69][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n64));
   AO22CHD U3121 (.O(n1696), 
	.B2(n187), 
	.B1(\ram[69][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n64));
   AO22CHD U3122 (.O(n1697), 
	.B2(n187), 
	.B1(\ram[69][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n64));
   AO22CHD U3123 (.O(n1698), 
	.B2(n187), 
	.B1(\ram[69][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n64));
   AO22CHD U3124 (.O(n1699), 
	.B2(n187), 
	.B1(\ram[69][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n64));
   AO22CHD U3125 (.O(n1700), 
	.B2(n187), 
	.B1(\ram[69][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n64));
   AO22CHD U3126 (.O(n1701), 
	.B2(n187), 
	.B1(\ram[69][15] ), 
	.A2(n23), 
	.A1(n64));
   AO22CHD U3127 (.O(n1702), 
	.B2(n189), 
	.B1(\ram[70][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n65));
   AO22CHD U3128 (.O(n1703), 
	.B2(n189), 
	.B1(\ram[70][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n65));
   AO22CHD U3129 (.O(n1704), 
	.B2(n189), 
	.B1(\ram[70][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n65));
   AO22CHD U3130 (.O(n1705), 
	.B2(n189), 
	.B1(\ram[70][3] ), 
	.A2(n11), 
	.A1(n65));
   AO22CHD U3131 (.O(n1706), 
	.B2(n189), 
	.B1(\ram[70][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n65));
   AO22CHD U3132 (.O(n1707), 
	.B2(n189), 
	.B1(\ram[70][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n65));
   AO22CHD U3133 (.O(n1708), 
	.B2(n189), 
	.B1(\ram[70][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n65));
   AO22CHD U3134 (.O(n1709), 
	.B2(n189), 
	.B1(\ram[70][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n65));
   AO22CHD U3135 (.O(n1710), 
	.B2(n189), 
	.B1(\ram[70][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n65));
   AO22CHD U3136 (.O(n1711), 
	.B2(n189), 
	.B1(\ram[70][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n65));
   AO22CHD U3137 (.O(n1712), 
	.B2(n189), 
	.B1(\ram[70][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n65));
   AO22CHD U3138 (.O(n1713), 
	.B2(n189), 
	.B1(\ram[70][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n65));
   AO22CHD U3139 (.O(n1714), 
	.B2(n189), 
	.B1(\ram[70][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n65));
   AO22CHD U3140 (.O(n1715), 
	.B2(n189), 
	.B1(\ram[70][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n65));
   AO22CHD U3141 (.O(n1716), 
	.B2(n189), 
	.B1(\ram[70][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n65));
   AO22CHD U3142 (.O(n1717), 
	.B2(n189), 
	.B1(\ram[70][15] ), 
	.A2(n23), 
	.A1(n65));
   AO22CHD U3143 (.O(n1718), 
	.B2(n191), 
	.B1(\ram[71][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n67));
   AO22CHD U3144 (.O(n1719), 
	.B2(n191), 
	.B1(\ram[71][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n67));
   AO22CHD U3145 (.O(n1720), 
	.B2(n191), 
	.B1(\ram[71][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n67));
   AO22CHD U3146 (.O(n1721), 
	.B2(n191), 
	.B1(\ram[71][3] ), 
	.A2(n11), 
	.A1(n67));
   AO22CHD U3147 (.O(n1722), 
	.B2(n191), 
	.B1(\ram[71][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n67));
   AO22CHD U3148 (.O(n1723), 
	.B2(n191), 
	.B1(\ram[71][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n67));
   AO22CHD U3149 (.O(n1724), 
	.B2(n191), 
	.B1(\ram[71][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n67));
   AO22CHD U3150 (.O(n1725), 
	.B2(n191), 
	.B1(\ram[71][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n67));
   AO22CHD U3151 (.O(n1726), 
	.B2(n191), 
	.B1(\ram[71][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n67));
   AO22CHD U3152 (.O(n1727), 
	.B2(n191), 
	.B1(\ram[71][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n67));
   AO22CHD U3153 (.O(n1728), 
	.B2(n191), 
	.B1(\ram[71][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n67));
   AO22CHD U3154 (.O(n1729), 
	.B2(n191), 
	.B1(\ram[71][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n67));
   AO22CHD U3155 (.O(n1730), 
	.B2(n191), 
	.B1(\ram[71][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n67));
   AO22CHD U3156 (.O(n1731), 
	.B2(n191), 
	.B1(\ram[71][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n67));
   AO22CHD U3157 (.O(n1732), 
	.B2(n191), 
	.B1(\ram[71][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n67));
   AO22CHD U3158 (.O(n1733), 
	.B2(n191), 
	.B1(\ram[71][15] ), 
	.A2(n23), 
	.A1(n67));
   AO22CHD U3159 (.O(n1734), 
	.B2(n193), 
	.B1(\ram[72][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n68));
   AO22CHD U3160 (.O(n1735), 
	.B2(n193), 
	.B1(\ram[72][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n68));
   AO22CHD U3161 (.O(n1736), 
	.B2(n193), 
	.B1(\ram[72][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n68));
   AO22CHD U3162 (.O(n1737), 
	.B2(n193), 
	.B1(\ram[72][3] ), 
	.A2(n11), 
	.A1(n68));
   AO22CHD U3163 (.O(n1738), 
	.B2(n193), 
	.B1(\ram[72][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n68));
   AO22CHD U3164 (.O(n1739), 
	.B2(n193), 
	.B1(\ram[72][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n68));
   AO22CHD U3165 (.O(n1740), 
	.B2(n193), 
	.B1(\ram[72][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n68));
   AO22CHD U3166 (.O(n1741), 
	.B2(n193), 
	.B1(\ram[72][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n68));
   AO22CHD U3167 (.O(n1742), 
	.B2(n193), 
	.B1(\ram[72][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n68));
   AO22CHD U3168 (.O(n1743), 
	.B2(n193), 
	.B1(\ram[72][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n68));
   AO22CHD U3169 (.O(n1744), 
	.B2(n193), 
	.B1(\ram[72][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n68));
   AO22CHD U3170 (.O(n1745), 
	.B2(n193), 
	.B1(\ram[72][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n68));
   AO22CHD U3171 (.O(n1746), 
	.B2(n193), 
	.B1(\ram[72][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n68));
   AO22CHD U3172 (.O(n1747), 
	.B2(n193), 
	.B1(\ram[72][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n68));
   AO22CHD U3173 (.O(n1748), 
	.B2(n193), 
	.B1(\ram[72][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n68));
   AO22CHD U3174 (.O(n1749), 
	.B2(n193), 
	.B1(\ram[72][15] ), 
	.A2(n23), 
	.A1(n68));
   AO22CHD U3175 (.O(n1750), 
	.B2(n195), 
	.B1(\ram[73][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n70));
   AO22CHD U3176 (.O(n1751), 
	.B2(n195), 
	.B1(\ram[73][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n70));
   AO22CHD U3177 (.O(n1752), 
	.B2(n195), 
	.B1(\ram[73][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n70));
   AO22CHD U3178 (.O(n1753), 
	.B2(n195), 
	.B1(\ram[73][3] ), 
	.A2(n11), 
	.A1(n70));
   AO22CHD U3179 (.O(n1754), 
	.B2(n195), 
	.B1(\ram[73][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n70));
   AO22CHD U3180 (.O(n1755), 
	.B2(n195), 
	.B1(\ram[73][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n70));
   AO22CHD U3181 (.O(n1756), 
	.B2(n195), 
	.B1(\ram[73][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n70));
   AO22CHD U3182 (.O(n1757), 
	.B2(n195), 
	.B1(\ram[73][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n70));
   AO22CHD U3183 (.O(n1758), 
	.B2(n195), 
	.B1(\ram[73][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n70));
   AO22CHD U3184 (.O(n1759), 
	.B2(n195), 
	.B1(\ram[73][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n70));
   AO22CHD U3185 (.O(n1760), 
	.B2(n195), 
	.B1(\ram[73][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n70));
   AO22CHD U3186 (.O(n1761), 
	.B2(n195), 
	.B1(\ram[73][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n70));
   AO22CHD U3187 (.O(n1762), 
	.B2(n195), 
	.B1(\ram[73][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n70));
   AO22CHD U3188 (.O(n1763), 
	.B2(n195), 
	.B1(\ram[73][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n70));
   AO22CHD U3189 (.O(n1764), 
	.B2(n195), 
	.B1(\ram[73][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n70));
   AO22CHD U3190 (.O(n1765), 
	.B2(n195), 
	.B1(\ram[73][15] ), 
	.A2(n23), 
	.A1(n70));
   AO22CHD U3191 (.O(n1766), 
	.B2(n197), 
	.B1(\ram[74][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n73));
   AO22CHD U3192 (.O(n1767), 
	.B2(n197), 
	.B1(\ram[74][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n73));
   AO22CHD U3193 (.O(n1768), 
	.B2(n197), 
	.B1(\ram[74][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n73));
   AO22CHD U3194 (.O(n1769), 
	.B2(n197), 
	.B1(\ram[74][3] ), 
	.A2(n11), 
	.A1(n73));
   AO22CHD U3195 (.O(n1770), 
	.B2(n197), 
	.B1(\ram[74][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n73));
   AO22CHD U3196 (.O(n1771), 
	.B2(n197), 
	.B1(\ram[74][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n73));
   AO22CHD U3197 (.O(n1772), 
	.B2(n197), 
	.B1(\ram[74][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n73));
   AO22CHD U3198 (.O(n1773), 
	.B2(n197), 
	.B1(\ram[74][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n73));
   AO22CHD U3199 (.O(n1774), 
	.B2(n197), 
	.B1(\ram[74][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n73));
   AO22CHD U3200 (.O(n1775), 
	.B2(n197), 
	.B1(\ram[74][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n73));
   AO22CHD U3201 (.O(n1776), 
	.B2(n197), 
	.B1(\ram[74][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n73));
   AO22CHD U3202 (.O(n1777), 
	.B2(n197), 
	.B1(\ram[74][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n73));
   AO22CHD U3203 (.O(n1778), 
	.B2(n197), 
	.B1(\ram[74][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n73));
   AO22CHD U3204 (.O(n1779), 
	.B2(n197), 
	.B1(\ram[74][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n73));
   AO22CHD U3205 (.O(n1780), 
	.B2(n197), 
	.B1(\ram[74][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n73));
   AO22CHD U3206 (.O(n1781), 
	.B2(n197), 
	.B1(\ram[74][15] ), 
	.A2(n23), 
	.A1(n73));
   AO22CHD U3207 (.O(n1782), 
	.B2(n199), 
	.B1(\ram[75][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n75));
   AO22CHD U3208 (.O(n1783), 
	.B2(n199), 
	.B1(\ram[75][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n75));
   AO22CHD U3209 (.O(n1784), 
	.B2(n199), 
	.B1(\ram[75][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n75));
   AO22CHD U3210 (.O(n1785), 
	.B2(n199), 
	.B1(\ram[75][3] ), 
	.A2(n11), 
	.A1(n75));
   AO22CHD U3211 (.O(n1786), 
	.B2(n199), 
	.B1(\ram[75][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n75));
   AO22CHD U3212 (.O(n1787), 
	.B2(n199), 
	.B1(\ram[75][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n75));
   AO22CHD U3213 (.O(n1788), 
	.B2(n199), 
	.B1(\ram[75][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n75));
   AO22CHD U3214 (.O(n1789), 
	.B2(n199), 
	.B1(\ram[75][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n75));
   AO22CHD U3215 (.O(n1790), 
	.B2(n199), 
	.B1(\ram[75][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n75));
   AO22CHD U3216 (.O(n1791), 
	.B2(n199), 
	.B1(\ram[75][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n75));
   AO22CHD U3217 (.O(n1792), 
	.B2(n199), 
	.B1(\ram[75][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n75));
   AO22CHD U3218 (.O(n1793), 
	.B2(n199), 
	.B1(\ram[75][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n75));
   AO22CHD U3219 (.O(n1794), 
	.B2(n199), 
	.B1(\ram[75][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n75));
   AO22CHD U3220 (.O(n1795), 
	.B2(n199), 
	.B1(\ram[75][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n75));
   AO22CHD U3221 (.O(n1796), 
	.B2(n199), 
	.B1(\ram[75][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n75));
   AO22CHD U3222 (.O(n1797), 
	.B2(n199), 
	.B1(\ram[75][15] ), 
	.A2(n23), 
	.A1(n75));
   AO22CHD U3223 (.O(n1798), 
	.B2(n201), 
	.B1(\ram[76][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n76));
   AO22CHD U3224 (.O(n1799), 
	.B2(n201), 
	.B1(\ram[76][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n76));
   AO22CHD U3225 (.O(n1800), 
	.B2(n201), 
	.B1(\ram[76][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n76));
   AO22CHD U3226 (.O(n1801), 
	.B2(n201), 
	.B1(\ram[76][3] ), 
	.A2(n11), 
	.A1(n76));
   AO22CHD U3227 (.O(n1802), 
	.B2(n201), 
	.B1(\ram[76][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n76));
   AO22CHD U3228 (.O(n1803), 
	.B2(n201), 
	.B1(\ram[76][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n76));
   AO22CHD U3229 (.O(n1804), 
	.B2(n201), 
	.B1(\ram[76][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n76));
   AO22CHD U3230 (.O(n1805), 
	.B2(n201), 
	.B1(\ram[76][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n76));
   AO22CHD U3231 (.O(n1806), 
	.B2(n201), 
	.B1(\ram[76][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n76));
   AO22CHD U3232 (.O(n1807), 
	.B2(n201), 
	.B1(\ram[76][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n76));
   AO22CHD U3233 (.O(n1808), 
	.B2(n201), 
	.B1(\ram[76][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n76));
   AO22CHD U3234 (.O(n1809), 
	.B2(n201), 
	.B1(\ram[76][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n76));
   AO22CHD U3235 (.O(n1810), 
	.B2(n201), 
	.B1(\ram[76][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n76));
   AO22CHD U3236 (.O(n1811), 
	.B2(n201), 
	.B1(\ram[76][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n76));
   AO22CHD U3237 (.O(n1812), 
	.B2(n201), 
	.B1(\ram[76][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n76));
   AO22CHD U3238 (.O(n1813), 
	.B2(n201), 
	.B1(\ram[76][15] ), 
	.A2(n23), 
	.A1(n76));
   AO22CHD U3239 (.O(n1814), 
	.B2(n203), 
	.B1(\ram[77][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n78));
   AO22CHD U3240 (.O(n1815), 
	.B2(n203), 
	.B1(\ram[77][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n78));
   AO22CHD U3241 (.O(n1816), 
	.B2(n203), 
	.B1(\ram[77][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n78));
   AO22CHD U3242 (.O(n1817), 
	.B2(n203), 
	.B1(\ram[77][3] ), 
	.A2(n11), 
	.A1(n78));
   AO22CHD U3243 (.O(n1818), 
	.B2(n203), 
	.B1(\ram[77][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n78));
   AO22CHD U3244 (.O(n1819), 
	.B2(n203), 
	.B1(\ram[77][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n78));
   AO22CHD U3245 (.O(n1820), 
	.B2(n203), 
	.B1(\ram[77][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n78));
   AO22CHD U3246 (.O(n1821), 
	.B2(n203), 
	.B1(\ram[77][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n78));
   AO22CHD U3247 (.O(n1822), 
	.B2(n203), 
	.B1(\ram[77][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n78));
   AO22CHD U3248 (.O(n1823), 
	.B2(n203), 
	.B1(\ram[77][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n78));
   AO22CHD U3249 (.O(n1824), 
	.B2(n203), 
	.B1(\ram[77][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n78));
   AO22CHD U3250 (.O(n1825), 
	.B2(n203), 
	.B1(\ram[77][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n78));
   AO22CHD U3251 (.O(n1826), 
	.B2(n203), 
	.B1(\ram[77][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n78));
   AO22CHD U3252 (.O(n1827), 
	.B2(n203), 
	.B1(\ram[77][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n78));
   AO22CHD U3253 (.O(n1828), 
	.B2(n203), 
	.B1(\ram[77][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n78));
   AO22CHD U3254 (.O(n1829), 
	.B2(n203), 
	.B1(\ram[77][15] ), 
	.A2(n23), 
	.A1(n78));
   AO22CHD U3255 (.O(n1830), 
	.B2(n205), 
	.B1(\ram[78][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n80));
   AO22CHD U3256 (.O(n1831), 
	.B2(n205), 
	.B1(\ram[78][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n80));
   AO22CHD U3257 (.O(n1832), 
	.B2(n205), 
	.B1(\ram[78][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n80));
   AO22CHD U3258 (.O(n1833), 
	.B2(n205), 
	.B1(\ram[78][3] ), 
	.A2(n11), 
	.A1(n80));
   AO22CHD U3259 (.O(n1834), 
	.B2(n205), 
	.B1(\ram[78][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n80));
   AO22CHD U3260 (.O(n1835), 
	.B2(n205), 
	.B1(\ram[78][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n80));
   AO22CHD U3261 (.O(n1836), 
	.B2(n205), 
	.B1(\ram[78][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n80));
   AO22CHD U3262 (.O(n1837), 
	.B2(n205), 
	.B1(\ram[78][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n80));
   AO22CHD U3263 (.O(n1838), 
	.B2(n205), 
	.B1(FE_PHN2851_ram_78__8_), 
	.A2(FE_OFN67_n16), 
	.A1(n80));
   AO22CHD U3264 (.O(n1839), 
	.B2(n205), 
	.B1(\ram[78][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n80));
   AO22CHD U3265 (.O(n1840), 
	.B2(n205), 
	.B1(\ram[78][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n80));
   AO22CHD U3266 (.O(n1841), 
	.B2(n205), 
	.B1(\ram[78][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n80));
   AO22CHD U3267 (.O(n1842), 
	.B2(n205), 
	.B1(\ram[78][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n80));
   AO22CHD U3268 (.O(n1843), 
	.B2(n205), 
	.B1(\ram[78][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n80));
   AO22CHD U3269 (.O(n1844), 
	.B2(n205), 
	.B1(\ram[78][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n80));
   AO22CHD U3270 (.O(n1845), 
	.B2(n205), 
	.B1(\ram[78][15] ), 
	.A2(n23), 
	.A1(n80));
   AO22CHD U3271 (.O(n1846), 
	.B2(n207), 
	.B1(\ram[79][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n82));
   AO22CHD U3272 (.O(n1847), 
	.B2(n207), 
	.B1(\ram[79][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n82));
   AO22CHD U3273 (.O(n1848), 
	.B2(n207), 
	.B1(\ram[79][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n82));
   AO22CHD U3274 (.O(n1849), 
	.B2(n207), 
	.B1(\ram[79][3] ), 
	.A2(n11), 
	.A1(n82));
   AO22CHD U3275 (.O(n1850), 
	.B2(n207), 
	.B1(\ram[79][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n82));
   AO22CHD U3276 (.O(n1851), 
	.B2(n207), 
	.B1(\ram[79][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n82));
   AO22CHD U3277 (.O(n1852), 
	.B2(n207), 
	.B1(\ram[79][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n82));
   AO22CHD U3278 (.O(n1853), 
	.B2(n207), 
	.B1(\ram[79][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n82));
   AO22CHD U3279 (.O(n1854), 
	.B2(n207), 
	.B1(\ram[79][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n82));
   AO22CHD U3280 (.O(n1855), 
	.B2(n207), 
	.B1(\ram[79][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n82));
   AO22CHD U3281 (.O(n1856), 
	.B2(n207), 
	.B1(\ram[79][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n82));
   AO22CHD U3282 (.O(n1857), 
	.B2(n207), 
	.B1(\ram[79][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n82));
   AO22CHD U3283 (.O(n1858), 
	.B2(n207), 
	.B1(\ram[79][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n82));
   AO22CHD U3284 (.O(n1859), 
	.B2(n207), 
	.B1(\ram[79][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n82));
   AO22CHD U3285 (.O(n1860), 
	.B2(n207), 
	.B1(\ram[79][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n82));
   AO22CHD U3286 (.O(n1861), 
	.B2(n207), 
	.B1(\ram[79][15] ), 
	.A2(n23), 
	.A1(n82));
   AO22CHD U3287 (.O(n1862), 
	.B2(n210), 
	.B1(\ram[80][0] ), 
	.A2(n6), 
	.A1(n84));
   AO22CHD U3288 (.O(n1863), 
	.B2(n210), 
	.B1(\ram[80][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n84));
   AO22CHD U3289 (.O(n1864), 
	.B2(n210), 
	.B1(\ram[80][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n84));
   AO22CHD U3290 (.O(n1865), 
	.B2(n210), 
	.B1(\ram[80][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n84));
   AO22CHD U3291 (.O(n1866), 
	.B2(n210), 
	.B1(\ram[80][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n84));
   AO22CHD U3292 (.O(n1867), 
	.B2(n210), 
	.B1(\ram[80][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n84));
   AO22CHD U3293 (.O(n1868), 
	.B2(n210), 
	.B1(\ram[80][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n84));
   AO22CHD U3294 (.O(n1869), 
	.B2(n210), 
	.B1(\ram[80][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n84));
   AO22CHD U3295 (.O(n1870), 
	.B2(n210), 
	.B1(\ram[80][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n84));
   AO22CHD U3296 (.O(n1871), 
	.B2(n210), 
	.B1(\ram[80][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n84));
   AO22CHD U3297 (.O(n1872), 
	.B2(n210), 
	.B1(\ram[80][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n84));
   AO22CHD U3298 (.O(n1873), 
	.B2(n210), 
	.B1(\ram[80][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n84));
   AO22CHD U3299 (.O(n1874), 
	.B2(n210), 
	.B1(\ram[80][12] ), 
	.A2(n20), 
	.A1(n84));
   AO22CHD U3300 (.O(n1875), 
	.B2(n210), 
	.B1(\ram[80][13] ), 
	.A2(n21), 
	.A1(n84));
   AO22CHD U3301 (.O(n1876), 
	.B2(n210), 
	.B1(\ram[80][14] ), 
	.A2(n22), 
	.A1(n84));
   AO22CHD U3302 (.O(n1877), 
	.B2(n210), 
	.B1(\ram[80][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n84));
   AO22CHD U3303 (.O(n1878), 
	.B2(n213), 
	.B1(\ram[81][0] ), 
	.A2(n6), 
	.A1(n86));
   AO22CHD U3304 (.O(n1879), 
	.B2(n213), 
	.B1(FE_PHN2454_ram_81__1_), 
	.A2(FE_OFN44_n9), 
	.A1(n86));
   AO22CHD U3305 (.O(n1880), 
	.B2(n213), 
	.B1(\ram[81][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n86));
   AO22CHD U3306 (.O(n1881), 
	.B2(n213), 
	.B1(\ram[81][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n86));
   AO22CHD U3307 (.O(n1882), 
	.B2(n213), 
	.B1(\ram[81][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n86));
   AO22CHD U3308 (.O(n1883), 
	.B2(n213), 
	.B1(\ram[81][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n86));
   AO22CHD U3309 (.O(n1884), 
	.B2(n213), 
	.B1(\ram[81][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n86));
   AO22CHD U3310 (.O(n1885), 
	.B2(n213), 
	.B1(\ram[81][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n86));
   AO22CHD U3311 (.O(n1886), 
	.B2(n213), 
	.B1(\ram[81][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n86));
   AO22CHD U3312 (.O(n1887), 
	.B2(n213), 
	.B1(\ram[81][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n86));
   AO22CHD U3313 (.O(n1888), 
	.B2(n213), 
	.B1(\ram[81][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n86));
   AO22CHD U3314 (.O(n1889), 
	.B2(n213), 
	.B1(\ram[81][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n86));
   AO22CHD U3315 (.O(n1890), 
	.B2(n213), 
	.B1(\ram[81][12] ), 
	.A2(n20), 
	.A1(n86));
   AO22CHD U3316 (.O(n1891), 
	.B2(n213), 
	.B1(FE_PHN1318_ram_81__13_), 
	.A2(n21), 
	.A1(n86));
   AO22CHD U3317 (.O(n1892), 
	.B2(n213), 
	.B1(\ram[81][14] ), 
	.A2(n22), 
	.A1(n86));
   AO22CHD U3318 (.O(n1893), 
	.B2(n213), 
	.B1(\ram[81][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n86));
   AO22CHD U3319 (.O(n1894), 
	.B2(n215), 
	.B1(\ram[82][0] ), 
	.A2(n6), 
	.A1(n88));
   AO22CHD U3320 (.O(n1895), 
	.B2(n215), 
	.B1(\ram[82][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n88));
   AO22CHD U3321 (.O(n1896), 
	.B2(n215), 
	.B1(\ram[82][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n88));
   AO22CHD U3322 (.O(n1897), 
	.B2(n215), 
	.B1(\ram[82][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n88));
   AO22CHD U3323 (.O(n1898), 
	.B2(n215), 
	.B1(\ram[82][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n88));
   AO22CHD U3324 (.O(n1899), 
	.B2(n215), 
	.B1(\ram[82][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n88));
   AO22CHD U3325 (.O(n1900), 
	.B2(n215), 
	.B1(\ram[82][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n88));
   AO22CHD U3326 (.O(n1901), 
	.B2(n215), 
	.B1(\ram[82][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n88));
   AO22CHD U3327 (.O(n1902), 
	.B2(n215), 
	.B1(\ram[82][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n88));
   AO22CHD U3328 (.O(n1903), 
	.B2(n215), 
	.B1(\ram[82][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n88));
   AO22CHD U3329 (.O(n1904), 
	.B2(n215), 
	.B1(\ram[82][10] ), 
	.A2(FE_OFN73_n18), 
	.A1(n88));
   AO22CHD U3330 (.O(n1905), 
	.B2(n215), 
	.B1(\ram[82][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n88));
   AO22CHD U3331 (.O(n1906), 
	.B2(n215), 
	.B1(\ram[82][12] ), 
	.A2(n20), 
	.A1(n88));
   AO22CHD U3332 (.O(n1907), 
	.B2(n215), 
	.B1(\ram[82][13] ), 
	.A2(n21), 
	.A1(n88));
   AO22CHD U3333 (.O(n1908), 
	.B2(n215), 
	.B1(\ram[82][14] ), 
	.A2(n22), 
	.A1(n88));
   AO22CHD U3334 (.O(n1909), 
	.B2(n215), 
	.B1(\ram[82][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n88));
   AO22CHD U3335 (.O(n1910), 
	.B2(n217), 
	.B1(\ram[83][0] ), 
	.A2(n6), 
	.A1(n90));
   AO22CHD U3336 (.O(n1911), 
	.B2(n217), 
	.B1(\ram[83][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n90));
   AO22CHD U3337 (.O(n1912), 
	.B2(n217), 
	.B1(\ram[83][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n90));
   AO22CHD U3338 (.O(n1913), 
	.B2(n217), 
	.B1(\ram[83][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n90));
   AO22CHD U3339 (.O(n1914), 
	.B2(n217), 
	.B1(\ram[83][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n90));
   AO22CHD U3340 (.O(n1915), 
	.B2(n217), 
	.B1(\ram[83][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n90));
   AO22CHD U3341 (.O(n1916), 
	.B2(n217), 
	.B1(\ram[83][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n90));
   AO22CHD U3342 (.O(n1917), 
	.B2(n217), 
	.B1(\ram[83][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n90));
   AO22CHD U3343 (.O(n1918), 
	.B2(n217), 
	.B1(\ram[83][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n90));
   AO22CHD U3344 (.O(n1919), 
	.B2(n217), 
	.B1(\ram[83][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n90));
   AO22CHD U3345 (.O(n1920), 
	.B2(n217), 
	.B1(\ram[83][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n90));
   AO22CHD U3346 (.O(n1921), 
	.B2(n217), 
	.B1(\ram[83][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n90));
   AO22CHD U3347 (.O(n1922), 
	.B2(n217), 
	.B1(\ram[83][12] ), 
	.A2(n20), 
	.A1(n90));
   AO22CHD U3348 (.O(n1923), 
	.B2(n217), 
	.B1(\ram[83][13] ), 
	.A2(n21), 
	.A1(n90));
   AO22CHD U3349 (.O(n1924), 
	.B2(n217), 
	.B1(\ram[83][14] ), 
	.A2(n22), 
	.A1(n90));
   AO22CHD U3350 (.O(n1925), 
	.B2(n217), 
	.B1(\ram[83][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n90));
   AO22CHD U3351 (.O(n1926), 
	.B2(n219), 
	.B1(\ram[84][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n92));
   AO22CHD U3352 (.O(n1927), 
	.B2(n219), 
	.B1(\ram[84][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n92));
   AO22CHD U3353 (.O(n1928), 
	.B2(n219), 
	.B1(\ram[84][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n92));
   AO22CHD U3354 (.O(n1929), 
	.B2(n219), 
	.B1(\ram[84][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n92));
   AO22CHD U3355 (.O(n1930), 
	.B2(n219), 
	.B1(\ram[84][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n92));
   AO22CHD U3356 (.O(n1931), 
	.B2(n219), 
	.B1(\ram[84][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n92));
   AO22CHD U3357 (.O(n1932), 
	.B2(n219), 
	.B1(\ram[84][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n92));
   AO22CHD U3358 (.O(n1933), 
	.B2(n219), 
	.B1(\ram[84][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n92));
   AO22CHD U3359 (.O(n1934), 
	.B2(n219), 
	.B1(\ram[84][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n92));
   AO22CHD U3360 (.O(n1935), 
	.B2(n219), 
	.B1(\ram[84][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n92));
   AO22CHD U3361 (.O(n1936), 
	.B2(n219), 
	.B1(\ram[84][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n92));
   AO22CHD U3362 (.O(n1937), 
	.B2(n219), 
	.B1(\ram[84][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n92));
   AO22CHD U3363 (.O(n1938), 
	.B2(n219), 
	.B1(\ram[84][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n92));
   AO22CHD U3364 (.O(n1939), 
	.B2(n219), 
	.B1(\ram[84][13] ), 
	.A2(n21), 
	.A1(n92));
   AO22CHD U3365 (.O(n1940), 
	.B2(n219), 
	.B1(\ram[84][14] ), 
	.A2(n22), 
	.A1(n92));
   AO22CHD U3366 (.O(n1941), 
	.B2(n219), 
	.B1(\ram[84][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n92));
   AO22CHD U3367 (.O(n1942), 
	.B2(n221), 
	.B1(\ram[85][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n94));
   AO22CHD U3368 (.O(n1943), 
	.B2(n221), 
	.B1(\ram[85][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n94));
   AO22CHD U3369 (.O(n1944), 
	.B2(n221), 
	.B1(\ram[85][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n94));
   AO22CHD U3370 (.O(n1945), 
	.B2(n221), 
	.B1(\ram[85][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n94));
   AO22CHD U3371 (.O(n1946), 
	.B2(n221), 
	.B1(\ram[85][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n94));
   AO22CHD U3372 (.O(n1947), 
	.B2(n221), 
	.B1(\ram[85][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n94));
   AO22CHD U3373 (.O(n1948), 
	.B2(n221), 
	.B1(\ram[85][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n94));
   AO22CHD U3374 (.O(n1949), 
	.B2(n221), 
	.B1(\ram[85][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n94));
   AO22CHD U3375 (.O(n1950), 
	.B2(n221), 
	.B1(\ram[85][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n94));
   AO22CHD U3376 (.O(n1951), 
	.B2(n221), 
	.B1(\ram[85][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n94));
   AO22CHD U3377 (.O(n1952), 
	.B2(n221), 
	.B1(FE_PHN1962_ram_85__10_), 
	.A2(FE_OFN74_n18), 
	.A1(n94));
   AO22CHD U3378 (.O(n1953), 
	.B2(n221), 
	.B1(\ram[85][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n94));
   AO22CHD U3379 (.O(n1954), 
	.B2(n221), 
	.B1(\ram[85][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n94));
   AO22CHD U3380 (.O(n1955), 
	.B2(n221), 
	.B1(\ram[85][13] ), 
	.A2(n21), 
	.A1(n94));
   AO22CHD U3381 (.O(n1956), 
	.B2(n221), 
	.B1(\ram[85][14] ), 
	.A2(n22), 
	.A1(n94));
   AO22CHD U3382 (.O(n1957), 
	.B2(n221), 
	.B1(\ram[85][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n94));
   AO22CHD U3383 (.O(n1958), 
	.B2(n223), 
	.B1(\ram[86][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n96));
   AO22CHD U3384 (.O(n1959), 
	.B2(n223), 
	.B1(\ram[86][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n96));
   AO22CHD U3385 (.O(n1960), 
	.B2(n223), 
	.B1(\ram[86][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n96));
   AO22CHD U3386 (.O(n1961), 
	.B2(n223), 
	.B1(\ram[86][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n96));
   AO22CHD U3387 (.O(n1962), 
	.B2(n223), 
	.B1(\ram[86][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n96));
   AO22CHD U3388 (.O(n1963), 
	.B2(n223), 
	.B1(\ram[86][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n96));
   AO22CHD U3389 (.O(n1964), 
	.B2(n223), 
	.B1(\ram[86][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n96));
   AO22CHD U3390 (.O(n1965), 
	.B2(n223), 
	.B1(\ram[86][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n96));
   AO22CHD U3391 (.O(n1966), 
	.B2(n223), 
	.B1(\ram[86][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n96));
   AO22CHD U3392 (.O(n1967), 
	.B2(n223), 
	.B1(\ram[86][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n96));
   AO22CHD U3393 (.O(n1968), 
	.B2(n223), 
	.B1(\ram[86][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n96));
   AO22CHD U3394 (.O(n1969), 
	.B2(n223), 
	.B1(\ram[86][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n96));
   AO22CHD U3395 (.O(n1970), 
	.B2(n223), 
	.B1(\ram[86][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n96));
   AO22CHD U3396 (.O(n1971), 
	.B2(n223), 
	.B1(\ram[86][13] ), 
	.A2(n21), 
	.A1(n96));
   AO22CHD U3397 (.O(n1972), 
	.B2(n223), 
	.B1(\ram[86][14] ), 
	.A2(n22), 
	.A1(n96));
   AO22CHD U3398 (.O(n1973), 
	.B2(n223), 
	.B1(\ram[86][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n96));
   AO22CHD U3399 (.O(n1974), 
	.B2(n225), 
	.B1(\ram[87][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n98));
   AO22CHD U3400 (.O(n1975), 
	.B2(n225), 
	.B1(\ram[87][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n98));
   AO22CHD U3401 (.O(n1976), 
	.B2(n225), 
	.B1(\ram[87][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n98));
   AO22CHD U3402 (.O(n1977), 
	.B2(n225), 
	.B1(\ram[87][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n98));
   AO22CHD U3403 (.O(n1978), 
	.B2(n225), 
	.B1(\ram[87][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n98));
   AO22CHD U3404 (.O(n1979), 
	.B2(n225), 
	.B1(\ram[87][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n98));
   AO22CHD U3405 (.O(n1980), 
	.B2(n225), 
	.B1(\ram[87][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n98));
   AO22CHD U3406 (.O(n1981), 
	.B2(n225), 
	.B1(\ram[87][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n98));
   AO22CHD U3407 (.O(n1982), 
	.B2(n225), 
	.B1(\ram[87][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n98));
   AO22CHD U3408 (.O(n1983), 
	.B2(n225), 
	.B1(\ram[87][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n98));
   AO22CHD U3409 (.O(n1984), 
	.B2(n225), 
	.B1(\ram[87][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n98));
   AO22CHD U3410 (.O(n1985), 
	.B2(n225), 
	.B1(\ram[87][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n98));
   AO22CHD U3411 (.O(n1986), 
	.B2(n225), 
	.B1(\ram[87][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n98));
   AO22CHD U3412 (.O(n1987), 
	.B2(n225), 
	.B1(\ram[87][13] ), 
	.A2(n21), 
	.A1(n98));
   AO22CHD U3413 (.O(n1988), 
	.B2(n225), 
	.B1(\ram[87][14] ), 
	.A2(n22), 
	.A1(n98));
   AO22CHD U3414 (.O(n1989), 
	.B2(n225), 
	.B1(\ram[87][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n98));
   AO22CHD U3415 (.O(n1990), 
	.B2(n227), 
	.B1(\ram[88][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n100));
   AO22CHD U3416 (.O(n1991), 
	.B2(n227), 
	.B1(\ram[88][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n100));
   AO22CHD U3417 (.O(n1992), 
	.B2(n227), 
	.B1(\ram[88][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n100));
   AO22CHD U3418 (.O(n1993), 
	.B2(n227), 
	.B1(\ram[88][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n100));
   AO22CHD U3419 (.O(n1994), 
	.B2(n227), 
	.B1(\ram[88][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n100));
   AO22CHD U3420 (.O(n1995), 
	.B2(n227), 
	.B1(\ram[88][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n100));
   AO22CHD U3421 (.O(n1996), 
	.B2(n227), 
	.B1(\ram[88][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n100));
   AO22CHD U3422 (.O(n1997), 
	.B2(n227), 
	.B1(\ram[88][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n100));
   AO22CHD U3423 (.O(n1998), 
	.B2(n227), 
	.B1(\ram[88][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n100));
   AO22CHD U3424 (.O(n1999), 
	.B2(n227), 
	.B1(\ram[88][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n100));
   AO22CHD U3425 (.O(n2000), 
	.B2(n227), 
	.B1(\ram[88][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n100));
   AO22CHD U3426 (.O(n2001), 
	.B2(n227), 
	.B1(\ram[88][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n100));
   AO22CHD U3427 (.O(n2002), 
	.B2(n227), 
	.B1(\ram[88][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n100));
   AO22CHD U3428 (.O(n2003), 
	.B2(n227), 
	.B1(\ram[88][13] ), 
	.A2(n21), 
	.A1(n100));
   AO22CHD U3429 (.O(n2004), 
	.B2(n227), 
	.B1(\ram[88][14] ), 
	.A2(n22), 
	.A1(n100));
   AO22CHD U3430 (.O(n2005), 
	.B2(n227), 
	.B1(\ram[88][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n100));
   AO22CHD U3431 (.O(n2006), 
	.B2(n229), 
	.B1(\ram[89][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n102));
   AO22CHD U3432 (.O(n2007), 
	.B2(n229), 
	.B1(\ram[89][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n102));
   AO22CHD U3433 (.O(n2008), 
	.B2(n229), 
	.B1(\ram[89][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n102));
   AO22CHD U3434 (.O(n2009), 
	.B2(n229), 
	.B1(\ram[89][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n102));
   AO22CHD U3435 (.O(n2010), 
	.B2(n229), 
	.B1(\ram[89][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n102));
   AO22CHD U3436 (.O(n2011), 
	.B2(n229), 
	.B1(\ram[89][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n102));
   AO22CHD U3437 (.O(n2012), 
	.B2(n229), 
	.B1(\ram[89][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n102));
   AO22CHD U3438 (.O(n2013), 
	.B2(n229), 
	.B1(\ram[89][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n102));
   AO22CHD U3439 (.O(n2014), 
	.B2(n229), 
	.B1(\ram[89][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n102));
   AO22CHD U3440 (.O(n2015), 
	.B2(n229), 
	.B1(\ram[89][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n102));
   AO22CHD U3441 (.O(n2016), 
	.B2(n229), 
	.B1(\ram[89][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n102));
   AO22CHD U3442 (.O(n2017), 
	.B2(n229), 
	.B1(\ram[89][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n102));
   AO22CHD U3443 (.O(n2018), 
	.B2(n229), 
	.B1(\ram[89][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n102));
   AO22CHD U3444 (.O(n2019), 
	.B2(n229), 
	.B1(\ram[89][13] ), 
	.A2(n21), 
	.A1(n102));
   AO22CHD U3445 (.O(n2020), 
	.B2(n229), 
	.B1(\ram[89][14] ), 
	.A2(n22), 
	.A1(n102));
   AO22CHD U3446 (.O(n2021), 
	.B2(n229), 
	.B1(\ram[89][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n102));
   AO22CHD U3447 (.O(n2022), 
	.B2(n231), 
	.B1(\ram[90][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n104));
   AO22CHD U3448 (.O(n2023), 
	.B2(n231), 
	.B1(\ram[90][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n104));
   AO22CHD U3449 (.O(n2024), 
	.B2(n231), 
	.B1(\ram[90][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n104));
   AO22CHD U3450 (.O(n2025), 
	.B2(n231), 
	.B1(\ram[90][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n104));
   AO22CHD U3451 (.O(n2026), 
	.B2(n231), 
	.B1(\ram[90][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n104));
   AO22CHD U3452 (.O(n2027), 
	.B2(n231), 
	.B1(\ram[90][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n104));
   AO22CHD U3453 (.O(n2028), 
	.B2(n231), 
	.B1(\ram[90][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n104));
   AO22CHD U3454 (.O(n2029), 
	.B2(n231), 
	.B1(\ram[90][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n104));
   AO22CHD U3455 (.O(n2030), 
	.B2(n231), 
	.B1(\ram[90][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n104));
   AO22CHD U3456 (.O(n2031), 
	.B2(n231), 
	.B1(\ram[90][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n104));
   AO22CHD U3457 (.O(n2032), 
	.B2(n231), 
	.B1(\ram[90][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n104));
   AO22CHD U3458 (.O(n2033), 
	.B2(n231), 
	.B1(\ram[90][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n104));
   AO22CHD U3459 (.O(n2034), 
	.B2(n231), 
	.B1(\ram[90][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n104));
   AO22CHD U3460 (.O(n2035), 
	.B2(n231), 
	.B1(\ram[90][13] ), 
	.A2(n21), 
	.A1(n104));
   AO22CHD U3461 (.O(n2036), 
	.B2(n231), 
	.B1(\ram[90][14] ), 
	.A2(n22), 
	.A1(n104));
   AO22CHD U3462 (.O(n2037), 
	.B2(n231), 
	.B1(\ram[90][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n104));
   AO22CHD U3463 (.O(n2038), 
	.B2(n233), 
	.B1(\ram[91][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n107));
   AO22CHD U3464 (.O(n2039), 
	.B2(n233), 
	.B1(\ram[91][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n107));
   AO22CHD U3465 (.O(n2040), 
	.B2(n233), 
	.B1(\ram[91][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n107));
   AO22CHD U3466 (.O(n2041), 
	.B2(n233), 
	.B1(\ram[91][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n107));
   AO22CHD U3467 (.O(n2042), 
	.B2(n233), 
	.B1(\ram[91][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n107));
   AO22CHD U3468 (.O(n2043), 
	.B2(n233), 
	.B1(\ram[91][5] ), 
	.A2(FE_OFN58_n13), 
	.A1(n107));
   AO22CHD U3469 (.O(n2044), 
	.B2(n233), 
	.B1(\ram[91][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n107));
   AO22CHD U3470 (.O(n2045), 
	.B2(n233), 
	.B1(\ram[91][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n107));
   AO22CHD U3471 (.O(n2046), 
	.B2(n233), 
	.B1(\ram[91][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n107));
   AO22CHD U3472 (.O(n2047), 
	.B2(n233), 
	.B1(\ram[91][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n107));
   AO22CHD U3473 (.O(n2048), 
	.B2(n233), 
	.B1(\ram[91][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n107));
   AO22CHD U3474 (.O(n2049), 
	.B2(n233), 
	.B1(\ram[91][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n107));
   AO22CHD U3475 (.O(n2050), 
	.B2(n233), 
	.B1(\ram[91][12] ), 
	.A2(FE_OFN80_n20), 
	.A1(n107));
   AO22CHD U3476 (.O(n2051), 
	.B2(n233), 
	.B1(\ram[91][13] ), 
	.A2(n21), 
	.A1(n107));
   AO22CHD U3477 (.O(n2052), 
	.B2(n233), 
	.B1(\ram[91][14] ), 
	.A2(n22), 
	.A1(n107));
   AO22CHD U3478 (.O(n2053), 
	.B2(n233), 
	.B1(\ram[91][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n107));
   AO22CHD U3479 (.O(n2054), 
	.B2(n235), 
	.B1(\ram[92][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n109));
   AO22CHD U3480 (.O(n2055), 
	.B2(n235), 
	.B1(\ram[92][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n109));
   AO22CHD U3481 (.O(n2056), 
	.B2(n235), 
	.B1(\ram[92][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n109));
   AO22CHD U3482 (.O(n2057), 
	.B2(n235), 
	.B1(\ram[92][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n109));
   AO22CHD U3483 (.O(n2058), 
	.B2(n235), 
	.B1(\ram[92][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n109));
   AO22CHD U3484 (.O(n2059), 
	.B2(n235), 
	.B1(\ram[92][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n109));
   AO22CHD U3485 (.O(n2060), 
	.B2(n235), 
	.B1(\ram[92][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n109));
   AO22CHD U3486 (.O(n2061), 
	.B2(n235), 
	.B1(\ram[92][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n109));
   AO22CHD U3487 (.O(n2062), 
	.B2(n235), 
	.B1(\ram[92][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n109));
   AO22CHD U3488 (.O(n2063), 
	.B2(n235), 
	.B1(\ram[92][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n109));
   AO22CHD U3489 (.O(n2064), 
	.B2(n235), 
	.B1(\ram[92][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n109));
   AO22CHD U3490 (.O(n2065), 
	.B2(n235), 
	.B1(\ram[92][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n109));
   AO22CHD U3491 (.O(n2066), 
	.B2(n235), 
	.B1(\ram[92][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n109));
   AO22CHD U3492 (.O(n2067), 
	.B2(n235), 
	.B1(\ram[92][13] ), 
	.A2(n21), 
	.A1(n109));
   AO22CHD U3493 (.O(n2068), 
	.B2(n235), 
	.B1(\ram[92][14] ), 
	.A2(n22), 
	.A1(n109));
   AO22CHD U3494 (.O(n2069), 
	.B2(n235), 
	.B1(\ram[92][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n109));
   AO22CHD U3495 (.O(n2070), 
	.B2(n237), 
	.B1(\ram[93][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n110));
   AO22CHD U3496 (.O(n2071), 
	.B2(n237), 
	.B1(\ram[93][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n110));
   AO22CHD U3497 (.O(n2072), 
	.B2(n237), 
	.B1(\ram[93][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n110));
   AO22CHD U3498 (.O(n2073), 
	.B2(n237), 
	.B1(FE_PHN2597_ram_93__3_), 
	.A2(FE_OFN52_n11), 
	.A1(n110));
   AO22CHD U3499 (.O(n2074), 
	.B2(n237), 
	.B1(\ram[93][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n110));
   AO22CHD U3500 (.O(n2075), 
	.B2(n237), 
	.B1(\ram[93][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n110));
   AO22CHD U3501 (.O(n2076), 
	.B2(n237), 
	.B1(\ram[93][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n110));
   AO22CHD U3502 (.O(n2077), 
	.B2(n237), 
	.B1(\ram[93][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n110));
   AO22CHD U3503 (.O(n2078), 
	.B2(n237), 
	.B1(\ram[93][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n110));
   AO22CHD U3504 (.O(n2079), 
	.B2(n237), 
	.B1(\ram[93][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n110));
   AO22CHD U3505 (.O(n2080), 
	.B2(n237), 
	.B1(\ram[93][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n110));
   AO22CHD U3506 (.O(n2081), 
	.B2(n237), 
	.B1(\ram[93][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n110));
   AO22CHD U3507 (.O(n2082), 
	.B2(n237), 
	.B1(\ram[93][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n110));
   AO22CHD U3508 (.O(n2083), 
	.B2(n237), 
	.B1(\ram[93][13] ), 
	.A2(n21), 
	.A1(n110));
   AO22CHD U3509 (.O(n2084), 
	.B2(n237), 
	.B1(\ram[93][14] ), 
	.A2(n22), 
	.A1(n110));
   AO22CHD U3510 (.O(n2085), 
	.B2(n237), 
	.B1(\ram[93][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n110));
   AO22CHD U3511 (.O(n2086), 
	.B2(n239), 
	.B1(\ram[94][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n112));
   AO22CHD U3512 (.O(n2087), 
	.B2(n239), 
	.B1(\ram[94][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n112));
   AO22CHD U3513 (.O(n2088), 
	.B2(n239), 
	.B1(\ram[94][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n112));
   AO22CHD U3514 (.O(n2089), 
	.B2(n239), 
	.B1(\ram[94][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n112));
   AO22CHD U3515 (.O(n2090), 
	.B2(n239), 
	.B1(\ram[94][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n112));
   AO22CHD U3516 (.O(n2091), 
	.B2(n239), 
	.B1(\ram[94][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n112));
   AO22CHD U3517 (.O(n2092), 
	.B2(n239), 
	.B1(\ram[94][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n112));
   AO22CHD U3518 (.O(n2093), 
	.B2(n239), 
	.B1(\ram[94][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n112));
   AO22CHD U3519 (.O(n2094), 
	.B2(n239), 
	.B1(\ram[94][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n112));
   AO22CHD U3520 (.O(n2095), 
	.B2(n239), 
	.B1(\ram[94][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n112));
   AO22CHD U3521 (.O(n2096), 
	.B2(n239), 
	.B1(\ram[94][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n112));
   AO22CHD U3522 (.O(n2097), 
	.B2(n239), 
	.B1(\ram[94][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n112));
   AO22CHD U3523 (.O(n2098), 
	.B2(n239), 
	.B1(\ram[94][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n112));
   AO22CHD U3524 (.O(n2099), 
	.B2(n239), 
	.B1(\ram[94][13] ), 
	.A2(n21), 
	.A1(n112));
   AO22CHD U3525 (.O(n2100), 
	.B2(n239), 
	.B1(\ram[94][14] ), 
	.A2(n22), 
	.A1(n112));
   AO22CHD U3526 (.O(n2101), 
	.B2(n239), 
	.B1(\ram[94][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n112));
   AO22CHD U3527 (.O(n2102), 
	.B2(n241), 
	.B1(\ram[95][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n114));
   AO22CHD U3528 (.O(n2103), 
	.B2(n241), 
	.B1(\ram[95][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n114));
   AO22CHD U3529 (.O(n2104), 
	.B2(n241), 
	.B1(\ram[95][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n114));
   AO22CHD U3530 (.O(n2105), 
	.B2(n241), 
	.B1(\ram[95][3] ), 
	.A2(FE_OFN52_n11), 
	.A1(n114));
   AO22CHD U3531 (.O(n2106), 
	.B2(n241), 
	.B1(\ram[95][4] ), 
	.A2(FE_OFN55_n12), 
	.A1(n114));
   AO22CHD U3532 (.O(n2107), 
	.B2(n241), 
	.B1(\ram[95][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n114));
   AO22CHD U3533 (.O(n2108), 
	.B2(n241), 
	.B1(\ram[95][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n114));
   AO22CHD U3534 (.O(n2109), 
	.B2(n241), 
	.B1(\ram[95][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n114));
   AO22CHD U3535 (.O(n2110), 
	.B2(n241), 
	.B1(\ram[95][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n114));
   AO22CHD U3536 (.O(n2111), 
	.B2(n241), 
	.B1(\ram[95][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n114));
   AO22CHD U3537 (.O(n2112), 
	.B2(n241), 
	.B1(\ram[95][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n114));
   AO22CHD U3538 (.O(n2113), 
	.B2(n241), 
	.B1(\ram[95][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n114));
   AO22CHD U3539 (.O(n2114), 
	.B2(n241), 
	.B1(\ram[95][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n114));
   AO22CHD U3540 (.O(n2115), 
	.B2(n241), 
	.B1(\ram[95][13] ), 
	.A2(n21), 
	.A1(n114));
   AO22CHD U3541 (.O(n2116), 
	.B2(n241), 
	.B1(\ram[95][14] ), 
	.A2(n22), 
	.A1(n114));
   AO22CHD U3542 (.O(n2117), 
	.B2(n241), 
	.B1(\ram[95][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n114));
   AO22CHD U3543 (.O(n2118), 
	.B2(n243), 
	.B1(\ram[96][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n116));
   AO22CHD U3544 (.O(n2119), 
	.B2(n243), 
	.B1(\ram[96][1] ), 
	.A2(n9), 
	.A1(n116));
   AO22CHD U3545 (.O(n2120), 
	.B2(n243), 
	.B1(\ram[96][2] ), 
	.A2(n10), 
	.A1(n116));
   AO22CHD U3546 (.O(n2121), 
	.B2(n243), 
	.B1(\ram[96][3] ), 
	.A2(n11), 
	.A1(n116));
   AO22CHD U3547 (.O(n2122), 
	.B2(n243), 
	.B1(\ram[96][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n116));
   AO22CHD U3548 (.O(n2123), 
	.B2(n243), 
	.B1(\ram[96][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n116));
   AO22CHD U3549 (.O(n2124), 
	.B2(n243), 
	.B1(\ram[96][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n116));
   AO22CHD U3550 (.O(n2125), 
	.B2(n243), 
	.B1(\ram[96][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n116));
   AO22CHD U3551 (.O(n2126), 
	.B2(n243), 
	.B1(\ram[96][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n116));
   AO22CHD U3552 (.O(n2127), 
	.B2(n243), 
	.B1(\ram[96][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n116));
   AO22CHD U3553 (.O(n2128), 
	.B2(n243), 
	.B1(\ram[96][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n116));
   AO22CHD U3554 (.O(n2129), 
	.B2(n243), 
	.B1(\ram[96][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n116));
   AO22CHD U3555 (.O(n2130), 
	.B2(n243), 
	.B1(\ram[96][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n116));
   AO22CHD U3556 (.O(n2131), 
	.B2(n243), 
	.B1(\ram[96][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n116));
   AO22CHD U3557 (.O(n2132), 
	.B2(n243), 
	.B1(\ram[96][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n116));
   AO22CHD U3558 (.O(n2133), 
	.B2(n243), 
	.B1(\ram[96][15] ), 
	.A2(n23), 
	.A1(n116));
   AO22CHD U3559 (.O(n2134), 
	.B2(n246), 
	.B1(\ram[97][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n118));
   AO22CHD U3560 (.O(n2135), 
	.B2(n246), 
	.B1(\ram[97][1] ), 
	.A2(n9), 
	.A1(n118));
   AO22CHD U3561 (.O(n2136), 
	.B2(n246), 
	.B1(\ram[97][2] ), 
	.A2(n10), 
	.A1(n118));
   AO22CHD U3562 (.O(n2137), 
	.B2(n246), 
	.B1(\ram[97][3] ), 
	.A2(n11), 
	.A1(n118));
   AO22CHD U3563 (.O(n2138), 
	.B2(n246), 
	.B1(\ram[97][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n118));
   AO22CHD U3564 (.O(n2139), 
	.B2(n246), 
	.B1(\ram[97][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n118));
   AO22CHD U3565 (.O(n2140), 
	.B2(n246), 
	.B1(\ram[97][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n118));
   AO22CHD U3566 (.O(n2141), 
	.B2(n246), 
	.B1(\ram[97][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n118));
   AO22CHD U3567 (.O(n2142), 
	.B2(n246), 
	.B1(\ram[97][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n118));
   AO22CHD U3568 (.O(n2143), 
	.B2(n246), 
	.B1(\ram[97][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n118));
   AO22CHD U3569 (.O(n2144), 
	.B2(n246), 
	.B1(\ram[97][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n118));
   AO22CHD U3570 (.O(n2145), 
	.B2(n246), 
	.B1(\ram[97][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n118));
   AO22CHD U3571 (.O(n2146), 
	.B2(n246), 
	.B1(\ram[97][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n118));
   AO22CHD U3572 (.O(n2147), 
	.B2(n246), 
	.B1(\ram[97][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n118));
   AO22CHD U3573 (.O(n2148), 
	.B2(n246), 
	.B1(\ram[97][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n118));
   AO22CHD U3574 (.O(n2149), 
	.B2(n246), 
	.B1(\ram[97][15] ), 
	.A2(n23), 
	.A1(n118));
   AO22CHD U3575 (.O(n2150), 
	.B2(n248), 
	.B1(\ram[98][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n120));
   AO22CHD U3576 (.O(n2151), 
	.B2(n248), 
	.B1(\ram[98][1] ), 
	.A2(n9), 
	.A1(n120));
   AO22CHD U3577 (.O(n2152), 
	.B2(n248), 
	.B1(\ram[98][2] ), 
	.A2(n10), 
	.A1(n120));
   AO22CHD U3578 (.O(n2153), 
	.B2(n248), 
	.B1(FE_PHN4971_ram_98__3_), 
	.A2(n11), 
	.A1(n120));
   AO22CHD U3579 (.O(n2154), 
	.B2(n248), 
	.B1(\ram[98][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n120));
   AO22CHD U3580 (.O(n2155), 
	.B2(n248), 
	.B1(\ram[98][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n120));
   AO22CHD U3581 (.O(n2156), 
	.B2(n248), 
	.B1(\ram[98][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n120));
   AO22CHD U3582 (.O(n2157), 
	.B2(n248), 
	.B1(\ram[98][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n120));
   AO22CHD U3583 (.O(n2158), 
	.B2(n248), 
	.B1(\ram[98][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n120));
   AO22CHD U3584 (.O(n2159), 
	.B2(n248), 
	.B1(\ram[98][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n120));
   AO22CHD U3585 (.O(n2160), 
	.B2(n248), 
	.B1(\ram[98][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n120));
   AO22CHD U3586 (.O(n2161), 
	.B2(n248), 
	.B1(\ram[98][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n120));
   AO22CHD U3587 (.O(n2162), 
	.B2(n248), 
	.B1(\ram[98][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n120));
   AO22CHD U3588 (.O(n2163), 
	.B2(n248), 
	.B1(\ram[98][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n120));
   AO22CHD U3589 (.O(n2164), 
	.B2(n248), 
	.B1(\ram[98][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n120));
   AO22CHD U3590 (.O(n2165), 
	.B2(n248), 
	.B1(\ram[98][15] ), 
	.A2(n23), 
	.A1(n120));
   AO22CHD U3591 (.O(n2166), 
	.B2(n250), 
	.B1(\ram[99][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n122));
   AO22CHD U3592 (.O(n2167), 
	.B2(n250), 
	.B1(\ram[99][1] ), 
	.A2(n9), 
	.A1(n122));
   AO22CHD U3593 (.O(n2168), 
	.B2(n250), 
	.B1(\ram[99][2] ), 
	.A2(n10), 
	.A1(n122));
   AO22CHD U3594 (.O(n2169), 
	.B2(n250), 
	.B1(\ram[99][3] ), 
	.A2(n11), 
	.A1(n122));
   AO22CHD U3595 (.O(n2170), 
	.B2(n250), 
	.B1(\ram[99][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n122));
   AO22CHD U3596 (.O(n2171), 
	.B2(n250), 
	.B1(\ram[99][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n122));
   AO22CHD U3597 (.O(n2172), 
	.B2(n250), 
	.B1(\ram[99][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n122));
   AO22CHD U3598 (.O(n2173), 
	.B2(n250), 
	.B1(\ram[99][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n122));
   AO22CHD U3599 (.O(n2174), 
	.B2(n250), 
	.B1(\ram[99][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n122));
   AO22CHD U3600 (.O(n2175), 
	.B2(n250), 
	.B1(\ram[99][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n122));
   AO22CHD U3601 (.O(n2176), 
	.B2(n250), 
	.B1(\ram[99][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n122));
   AO22CHD U3602 (.O(n2177), 
	.B2(n250), 
	.B1(\ram[99][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n122));
   AO22CHD U3603 (.O(n2178), 
	.B2(n250), 
	.B1(\ram[99][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n122));
   AO22CHD U3604 (.O(n2179), 
	.B2(n250), 
	.B1(\ram[99][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n122));
   AO22CHD U3605 (.O(n2180), 
	.B2(n250), 
	.B1(\ram[99][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n122));
   AO22CHD U3606 (.O(n2181), 
	.B2(n250), 
	.B1(\ram[99][15] ), 
	.A2(n23), 
	.A1(n122));
   AO22CHD U3607 (.O(n2182), 
	.B2(n252), 
	.B1(\ram[100][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n124));
   AO22CHD U3608 (.O(n2183), 
	.B2(n252), 
	.B1(\ram[100][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n124));
   AO22CHD U3609 (.O(n2184), 
	.B2(n252), 
	.B1(\ram[100][2] ), 
	.A2(n10), 
	.A1(n124));
   AO22CHD U3610 (.O(n2185), 
	.B2(n252), 
	.B1(\ram[100][3] ), 
	.A2(n11), 
	.A1(n124));
   AO22CHD U3611 (.O(n2186), 
	.B2(n252), 
	.B1(\ram[100][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n124));
   AO22CHD U3612 (.O(n2187), 
	.B2(n252), 
	.B1(\ram[100][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n124));
   AO22CHD U3613 (.O(n2188), 
	.B2(n252), 
	.B1(\ram[100][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n124));
   AO22CHD U3614 (.O(n2189), 
	.B2(n252), 
	.B1(\ram[100][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n124));
   AO22CHD U3615 (.O(n2190), 
	.B2(n252), 
	.B1(\ram[100][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n124));
   AO22CHD U3616 (.O(n2191), 
	.B2(n252), 
	.B1(\ram[100][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n124));
   AO22CHD U3617 (.O(n2192), 
	.B2(n252), 
	.B1(\ram[100][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n124));
   AO22CHD U3618 (.O(n2193), 
	.B2(n252), 
	.B1(\ram[100][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n124));
   AO22CHD U3619 (.O(n2194), 
	.B2(n252), 
	.B1(\ram[100][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n124));
   AO22CHD U3620 (.O(n2195), 
	.B2(n252), 
	.B1(\ram[100][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n124));
   AO22CHD U3621 (.O(n2196), 
	.B2(n252), 
	.B1(\ram[100][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n124));
   AO22CHD U3622 (.O(n2197), 
	.B2(n252), 
	.B1(\ram[100][15] ), 
	.A2(n23), 
	.A1(n124));
   AO22CHD U3623 (.O(n2198), 
	.B2(n254), 
	.B1(\ram[101][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n126));
   AO22CHD U3624 (.O(n2199), 
	.B2(n254), 
	.B1(\ram[101][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n126));
   AO22CHD U3625 (.O(n2200), 
	.B2(n254), 
	.B1(\ram[101][2] ), 
	.A2(n10), 
	.A1(n126));
   AO22CHD U3626 (.O(n2201), 
	.B2(n254), 
	.B1(\ram[101][3] ), 
	.A2(n11), 
	.A1(n126));
   AO22CHD U3627 (.O(n2202), 
	.B2(n254), 
	.B1(\ram[101][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n126));
   AO22CHD U3628 (.O(n2203), 
	.B2(n254), 
	.B1(\ram[101][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n126));
   AO22CHD U3629 (.O(n2204), 
	.B2(n254), 
	.B1(\ram[101][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n126));
   AO22CHD U3630 (.O(n2205), 
	.B2(n254), 
	.B1(\ram[101][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n126));
   AO22CHD U3631 (.O(n2206), 
	.B2(n254), 
	.B1(\ram[101][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n126));
   AO22CHD U3632 (.O(n2207), 
	.B2(n254), 
	.B1(\ram[101][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n126));
   AO22CHD U3633 (.O(n2208), 
	.B2(n254), 
	.B1(\ram[101][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n126));
   AO22CHD U3634 (.O(n2209), 
	.B2(n254), 
	.B1(\ram[101][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n126));
   AO22CHD U3635 (.O(n2210), 
	.B2(n254), 
	.B1(\ram[101][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n126));
   AO22CHD U3636 (.O(n2211), 
	.B2(n254), 
	.B1(\ram[101][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n126));
   AO22CHD U3637 (.O(n2212), 
	.B2(n254), 
	.B1(\ram[101][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n126));
   AO22CHD U3638 (.O(n2213), 
	.B2(n254), 
	.B1(\ram[101][15] ), 
	.A2(n23), 
	.A1(n126));
   AO22CHD U3639 (.O(n2214), 
	.B2(n256), 
	.B1(\ram[102][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n128));
   AO22CHD U3640 (.O(n2215), 
	.B2(n256), 
	.B1(\ram[102][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n128));
   AO22CHD U3641 (.O(n2216), 
	.B2(n256), 
	.B1(\ram[102][2] ), 
	.A2(n10), 
	.A1(n128));
   AO22CHD U3642 (.O(n2217), 
	.B2(n256), 
	.B1(\ram[102][3] ), 
	.A2(n11), 
	.A1(n128));
   AO22CHD U3643 (.O(n2218), 
	.B2(n256), 
	.B1(\ram[102][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n128));
   AO22CHD U3644 (.O(n2219), 
	.B2(n256), 
	.B1(\ram[102][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n128));
   AO22CHD U3645 (.O(n2220), 
	.B2(n256), 
	.B1(\ram[102][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n128));
   AO22CHD U3646 (.O(n2221), 
	.B2(n256), 
	.B1(\ram[102][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n128));
   AO22CHD U3647 (.O(n2222), 
	.B2(n256), 
	.B1(\ram[102][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n128));
   AO22CHD U3648 (.O(n2223), 
	.B2(n256), 
	.B1(\ram[102][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n128));
   AO22CHD U3649 (.O(n2224), 
	.B2(n256), 
	.B1(\ram[102][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n128));
   AO22CHD U3650 (.O(n2225), 
	.B2(n256), 
	.B1(\ram[102][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n128));
   AO22CHD U3651 (.O(n2226), 
	.B2(n256), 
	.B1(\ram[102][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n128));
   AO22CHD U3652 (.O(n2227), 
	.B2(n256), 
	.B1(\ram[102][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n128));
   AO22CHD U3653 (.O(n2228), 
	.B2(n256), 
	.B1(\ram[102][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n128));
   AO22CHD U3654 (.O(n2229), 
	.B2(n256), 
	.B1(\ram[102][15] ), 
	.A2(n23), 
	.A1(n128));
   AO22CHD U3655 (.O(n2230), 
	.B2(n258), 
	.B1(\ram[103][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n130));
   AO22CHD U3656 (.O(n2231), 
	.B2(n258), 
	.B1(\ram[103][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n130));
   AO22CHD U3657 (.O(n2232), 
	.B2(n258), 
	.B1(\ram[103][2] ), 
	.A2(n10), 
	.A1(n130));
   AO22CHD U3658 (.O(n2233), 
	.B2(n258), 
	.B1(\ram[103][3] ), 
	.A2(n11), 
	.A1(n130));
   AO22CHD U3659 (.O(n2234), 
	.B2(n258), 
	.B1(\ram[103][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n130));
   AO22CHD U3660 (.O(n2235), 
	.B2(n258), 
	.B1(\ram[103][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n130));
   AO22CHD U3661 (.O(n2236), 
	.B2(n258), 
	.B1(\ram[103][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n130));
   AO22CHD U3662 (.O(n2237), 
	.B2(n258), 
	.B1(\ram[103][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n130));
   AO22CHD U3663 (.O(n2238), 
	.B2(n258), 
	.B1(\ram[103][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n130));
   AO22CHD U3664 (.O(n2239), 
	.B2(n258), 
	.B1(\ram[103][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n130));
   AO22CHD U3665 (.O(n2240), 
	.B2(n258), 
	.B1(\ram[103][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n130));
   AO22CHD U3666 (.O(n2241), 
	.B2(n258), 
	.B1(\ram[103][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n130));
   AO22CHD U3667 (.O(n2242), 
	.B2(n258), 
	.B1(\ram[103][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n130));
   AO22CHD U3668 (.O(n2243), 
	.B2(n258), 
	.B1(\ram[103][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n130));
   AO22CHD U3669 (.O(n2244), 
	.B2(n258), 
	.B1(\ram[103][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n130));
   AO22CHD U3670 (.O(n2245), 
	.B2(n258), 
	.B1(\ram[103][15] ), 
	.A2(n23), 
	.A1(n130));
   AO22CHD U3671 (.O(n2246), 
	.B2(n260), 
	.B1(\ram[104][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n132));
   AO22CHD U3672 (.O(n2247), 
	.B2(n260), 
	.B1(\ram[104][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n132));
   AO22CHD U3673 (.O(n2248), 
	.B2(n260), 
	.B1(\ram[104][2] ), 
	.A2(n10), 
	.A1(n132));
   AO22CHD U3674 (.O(n2249), 
	.B2(n260), 
	.B1(\ram[104][3] ), 
	.A2(n11), 
	.A1(n132));
   AO22CHD U3675 (.O(n2250), 
	.B2(n260), 
	.B1(\ram[104][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n132));
   AO22CHD U3676 (.O(n2251), 
	.B2(n260), 
	.B1(\ram[104][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n132));
   AO22CHD U3677 (.O(n2252), 
	.B2(n260), 
	.B1(\ram[104][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n132));
   AO22CHD U3678 (.O(n2253), 
	.B2(n260), 
	.B1(\ram[104][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n132));
   AO22CHD U3679 (.O(n2254), 
	.B2(n260), 
	.B1(\ram[104][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n132));
   AO22CHD U3680 (.O(n2255), 
	.B2(n260), 
	.B1(\ram[104][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n132));
   AO22CHD U3681 (.O(n2256), 
	.B2(n260), 
	.B1(\ram[104][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n132));
   AO22CHD U3682 (.O(n2257), 
	.B2(n260), 
	.B1(\ram[104][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n132));
   AO22CHD U3683 (.O(n2258), 
	.B2(n260), 
	.B1(\ram[104][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n132));
   AO22CHD U3684 (.O(n2259), 
	.B2(n260), 
	.B1(FE_PHN2849_ram_104__13_), 
	.A2(FE_OFN83_n21), 
	.A1(n132));
   AO22CHD U3685 (.O(n2260), 
	.B2(n260), 
	.B1(\ram[104][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n132));
   AO22CHD U3686 (.O(n2261), 
	.B2(n260), 
	.B1(\ram[104][15] ), 
	.A2(n23), 
	.A1(n132));
   AO22CHD U3687 (.O(n2262), 
	.B2(n262), 
	.B1(\ram[105][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n134));
   AO22CHD U3688 (.O(n2263), 
	.B2(n262), 
	.B1(\ram[105][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n134));
   AO22CHD U3689 (.O(n2264), 
	.B2(n262), 
	.B1(\ram[105][2] ), 
	.A2(n10), 
	.A1(n134));
   AO22CHD U3690 (.O(n2265), 
	.B2(n262), 
	.B1(\ram[105][3] ), 
	.A2(n11), 
	.A1(n134));
   AO22CHD U3691 (.O(n2266), 
	.B2(n262), 
	.B1(\ram[105][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n134));
   AO22CHD U3692 (.O(n2267), 
	.B2(n262), 
	.B1(\ram[105][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n134));
   AO22CHD U3693 (.O(n2268), 
	.B2(n262), 
	.B1(\ram[105][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n134));
   AO22CHD U3694 (.O(n2269), 
	.B2(n262), 
	.B1(\ram[105][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n134));
   AO22CHD U3695 (.O(n2270), 
	.B2(n262), 
	.B1(\ram[105][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n134));
   AO22CHD U3696 (.O(n2271), 
	.B2(n262), 
	.B1(\ram[105][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n134));
   AO22CHD U3697 (.O(n2272), 
	.B2(n262), 
	.B1(\ram[105][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n134));
   AO22CHD U3698 (.O(n2273), 
	.B2(n262), 
	.B1(\ram[105][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n134));
   AO22CHD U3699 (.O(n2274), 
	.B2(n262), 
	.B1(\ram[105][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n134));
   AO22CHD U3700 (.O(n2275), 
	.B2(n262), 
	.B1(\ram[105][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n134));
   AO22CHD U3701 (.O(n2276), 
	.B2(n262), 
	.B1(\ram[105][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n134));
   AO22CHD U3702 (.O(n2277), 
	.B2(n262), 
	.B1(\ram[105][15] ), 
	.A2(n23), 
	.A1(n134));
   AO22CHD U3703 (.O(n2278), 
	.B2(n264), 
	.B1(\ram[106][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n136));
   AO22CHD U3704 (.O(n2279), 
	.B2(n264), 
	.B1(\ram[106][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n136));
   AO22CHD U3705 (.O(n2280), 
	.B2(n264), 
	.B1(\ram[106][2] ), 
	.A2(n10), 
	.A1(n136));
   AO22CHD U3706 (.O(n2281), 
	.B2(n264), 
	.B1(\ram[106][3] ), 
	.A2(n11), 
	.A1(n136));
   AO22CHD U3707 (.O(n2282), 
	.B2(n264), 
	.B1(\ram[106][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n136));
   AO22CHD U3708 (.O(n2283), 
	.B2(n264), 
	.B1(\ram[106][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n136));
   AO22CHD U3709 (.O(n2284), 
	.B2(n264), 
	.B1(\ram[106][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n136));
   AO22CHD U3710 (.O(n2285), 
	.B2(n264), 
	.B1(\ram[106][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n136));
   AO22CHD U3711 (.O(n2286), 
	.B2(n264), 
	.B1(\ram[106][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n136));
   AO22CHD U3712 (.O(n2287), 
	.B2(n264), 
	.B1(\ram[106][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n136));
   AO22CHD U3713 (.O(n2288), 
	.B2(n264), 
	.B1(\ram[106][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n136));
   AO22CHD U3714 (.O(n2289), 
	.B2(n264), 
	.B1(\ram[106][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n136));
   AO22CHD U3715 (.O(n2290), 
	.B2(n264), 
	.B1(\ram[106][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n136));
   AO22CHD U3716 (.O(n2291), 
	.B2(n264), 
	.B1(\ram[106][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n136));
   AO22CHD U3717 (.O(n2292), 
	.B2(n264), 
	.B1(\ram[106][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n136));
   AO22CHD U3718 (.O(n2293), 
	.B2(n264), 
	.B1(\ram[106][15] ), 
	.A2(n23), 
	.A1(n136));
   AO22CHD U3719 (.O(n2294), 
	.B2(n266), 
	.B1(\ram[107][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n138));
   AO22CHD U3720 (.O(n2295), 
	.B2(n266), 
	.B1(\ram[107][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n138));
   AO22CHD U3721 (.O(n2296), 
	.B2(n266), 
	.B1(\ram[107][2] ), 
	.A2(n10), 
	.A1(n138));
   AO22CHD U3722 (.O(n2297), 
	.B2(n266), 
	.B1(\ram[107][3] ), 
	.A2(n11), 
	.A1(n138));
   AO22CHD U3723 (.O(n2298), 
	.B2(n266), 
	.B1(\ram[107][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n138));
   AO22CHD U3724 (.O(n2299), 
	.B2(n266), 
	.B1(\ram[107][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n138));
   AO22CHD U3725 (.O(n2300), 
	.B2(n266), 
	.B1(\ram[107][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n138));
   AO22CHD U3726 (.O(n2301), 
	.B2(n266), 
	.B1(\ram[107][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n138));
   AO22CHD U3727 (.O(n2302), 
	.B2(n266), 
	.B1(\ram[107][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n138));
   AO22CHD U3728 (.O(n2303), 
	.B2(n266), 
	.B1(\ram[107][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n138));
   AO22CHD U3729 (.O(n2304), 
	.B2(n266), 
	.B1(\ram[107][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n138));
   AO22CHD U3730 (.O(n2305), 
	.B2(n266), 
	.B1(\ram[107][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n138));
   AO22CHD U3731 (.O(n2306), 
	.B2(n266), 
	.B1(\ram[107][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n138));
   AO22CHD U3732 (.O(n2307), 
	.B2(n266), 
	.B1(\ram[107][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n138));
   AO22CHD U3733 (.O(n2308), 
	.B2(n266), 
	.B1(\ram[107][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n138));
   AO22CHD U3734 (.O(n2309), 
	.B2(n266), 
	.B1(\ram[107][15] ), 
	.A2(n23), 
	.A1(n138));
   AO22CHD U3735 (.O(n2310), 
	.B2(n268), 
	.B1(\ram[108][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n141));
   AO22CHD U3736 (.O(n2311), 
	.B2(n268), 
	.B1(\ram[108][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n141));
   AO22CHD U3737 (.O(n2312), 
	.B2(n268), 
	.B1(\ram[108][2] ), 
	.A2(n10), 
	.A1(n141));
   AO22CHD U3738 (.O(n2313), 
	.B2(n268), 
	.B1(\ram[108][3] ), 
	.A2(n11), 
	.A1(n141));
   AO22CHD U3739 (.O(n2314), 
	.B2(n268), 
	.B1(\ram[108][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n141));
   AO22CHD U3740 (.O(n2315), 
	.B2(n268), 
	.B1(\ram[108][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n141));
   AO22CHD U3741 (.O(n2316), 
	.B2(n268), 
	.B1(\ram[108][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n141));
   AO22CHD U3742 (.O(n2317), 
	.B2(n268), 
	.B1(\ram[108][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n141));
   AO22CHD U3743 (.O(n2318), 
	.B2(n268), 
	.B1(\ram[108][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n141));
   AO22CHD U3744 (.O(n2319), 
	.B2(n268), 
	.B1(\ram[108][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n141));
   AO22CHD U3745 (.O(n2320), 
	.B2(n268), 
	.B1(\ram[108][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n141));
   AO22CHD U3746 (.O(n2321), 
	.B2(n268), 
	.B1(\ram[108][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n141));
   AO22CHD U3747 (.O(n2322), 
	.B2(n268), 
	.B1(\ram[108][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n141));
   AO22CHD U3748 (.O(n2323), 
	.B2(n268), 
	.B1(\ram[108][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n141));
   AO22CHD U3749 (.O(n2324), 
	.B2(n268), 
	.B1(\ram[108][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n141));
   AO22CHD U3750 (.O(n2325), 
	.B2(n268), 
	.B1(\ram[108][15] ), 
	.A2(n23), 
	.A1(n141));
   AO22CHD U3751 (.O(n2326), 
	.B2(n270), 
	.B1(\ram[109][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n143));
   AO22CHD U3752 (.O(n2327), 
	.B2(n270), 
	.B1(\ram[109][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n143));
   AO22CHD U3753 (.O(n2328), 
	.B2(n270), 
	.B1(\ram[109][2] ), 
	.A2(n10), 
	.A1(n143));
   AO22CHD U3754 (.O(n2329), 
	.B2(n270), 
	.B1(\ram[109][3] ), 
	.A2(n11), 
	.A1(n143));
   AO22CHD U3755 (.O(n2330), 
	.B2(n270), 
	.B1(\ram[109][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n143));
   AO22CHD U3756 (.O(n2331), 
	.B2(n270), 
	.B1(FE_PHN663_ram_109__5_), 
	.A2(FE_OFN57_n13), 
	.A1(n143));
   AO22CHD U3757 (.O(n2332), 
	.B2(n270), 
	.B1(\ram[109][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n143));
   AO22CHD U3758 (.O(n2333), 
	.B2(n270), 
	.B1(\ram[109][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n143));
   AO22CHD U3759 (.O(n2334), 
	.B2(n270), 
	.B1(\ram[109][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n143));
   AO22CHD U3760 (.O(n2335), 
	.B2(n270), 
	.B1(\ram[109][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n143));
   AO22CHD U3761 (.O(n2336), 
	.B2(n270), 
	.B1(\ram[109][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n143));
   AO22CHD U3762 (.O(n2337), 
	.B2(n270), 
	.B1(\ram[109][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n143));
   AO22CHD U3763 (.O(n2338), 
	.B2(n270), 
	.B1(\ram[109][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n143));
   AO22CHD U3764 (.O(n2339), 
	.B2(n270), 
	.B1(\ram[109][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n143));
   AO22CHD U3765 (.O(n2340), 
	.B2(n270), 
	.B1(\ram[109][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n143));
   AO22CHD U3766 (.O(n2341), 
	.B2(n270), 
	.B1(\ram[109][15] ), 
	.A2(n23), 
	.A1(n143));
   AO22CHD U3767 (.O(n2342), 
	.B2(n272), 
	.B1(\ram[110][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n144));
   AO22CHD U3768 (.O(n2343), 
	.B2(n272), 
	.B1(\ram[110][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n144));
   AO22CHD U3769 (.O(n2344), 
	.B2(n272), 
	.B1(\ram[110][2] ), 
	.A2(n10), 
	.A1(n144));
   AO22CHD U3770 (.O(n2345), 
	.B2(n272), 
	.B1(\ram[110][3] ), 
	.A2(n11), 
	.A1(n144));
   AO22CHD U3771 (.O(n2346), 
	.B2(n272), 
	.B1(\ram[110][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n144));
   AO22CHD U3772 (.O(n2347), 
	.B2(n272), 
	.B1(\ram[110][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n144));
   AO22CHD U3773 (.O(n2348), 
	.B2(n272), 
	.B1(\ram[110][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n144));
   AO22CHD U3774 (.O(n2349), 
	.B2(n272), 
	.B1(\ram[110][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n144));
   AO22CHD U3775 (.O(n2350), 
	.B2(n272), 
	.B1(\ram[110][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n144));
   AO22CHD U3776 (.O(n2351), 
	.B2(n272), 
	.B1(\ram[110][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n144));
   AO22CHD U3777 (.O(n2352), 
	.B2(n272), 
	.B1(\ram[110][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n144));
   AO22CHD U3778 (.O(n2353), 
	.B2(n272), 
	.B1(\ram[110][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n144));
   AO22CHD U3779 (.O(n2354), 
	.B2(n272), 
	.B1(\ram[110][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n144));
   AO22CHD U3780 (.O(n2355), 
	.B2(n272), 
	.B1(\ram[110][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n144));
   AO22CHD U3781 (.O(n2356), 
	.B2(n272), 
	.B1(\ram[110][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n144));
   AO22CHD U3782 (.O(n2357), 
	.B2(n272), 
	.B1(\ram[110][15] ), 
	.A2(n23), 
	.A1(n144));
   AO22CHD U3783 (.O(n2358), 
	.B2(n274), 
	.B1(\ram[111][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n146));
   AO22CHD U3784 (.O(n2359), 
	.B2(n274), 
	.B1(\ram[111][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n146));
   AO22CHD U3785 (.O(n2360), 
	.B2(n274), 
	.B1(\ram[111][2] ), 
	.A2(n10), 
	.A1(n146));
   AO22CHD U3786 (.O(n2361), 
	.B2(n274), 
	.B1(\ram[111][3] ), 
	.A2(n11), 
	.A1(n146));
   AO22CHD U3787 (.O(n2362), 
	.B2(n274), 
	.B1(\ram[111][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n146));
   AO22CHD U3788 (.O(n2363), 
	.B2(n274), 
	.B1(\ram[111][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n146));
   AO22CHD U3789 (.O(n2364), 
	.B2(n274), 
	.B1(\ram[111][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n146));
   AO22CHD U3790 (.O(n2365), 
	.B2(n274), 
	.B1(\ram[111][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n146));
   AO22CHD U3791 (.O(n2366), 
	.B2(n274), 
	.B1(\ram[111][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n146));
   AO22CHD U3792 (.O(n2367), 
	.B2(n274), 
	.B1(\ram[111][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n146));
   AO22CHD U3793 (.O(n2368), 
	.B2(n274), 
	.B1(\ram[111][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n146));
   AO22CHD U3794 (.O(n2369), 
	.B2(n274), 
	.B1(\ram[111][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n146));
   AO22CHD U3795 (.O(n2370), 
	.B2(n274), 
	.B1(\ram[111][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n146));
   AO22CHD U3796 (.O(n2371), 
	.B2(n274), 
	.B1(\ram[111][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n146));
   AO22CHD U3797 (.O(n2372), 
	.B2(n274), 
	.B1(\ram[111][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n146));
   AO22CHD U3798 (.O(n2373), 
	.B2(n274), 
	.B1(\ram[111][15] ), 
	.A2(n23), 
	.A1(n146));
   AO22CHD U3799 (.O(n2374), 
	.B2(n276), 
	.B1(\ram[112][0] ), 
	.A2(n6), 
	.A1(n148));
   AO22CHD U3800 (.O(n2375), 
	.B2(n276), 
	.B1(\ram[112][1] ), 
	.A2(n9), 
	.A1(n148));
   AO22CHD U3801 (.O(n2376), 
	.B2(n276), 
	.B1(\ram[112][2] ), 
	.A2(n10), 
	.A1(n148));
   AO22CHD U3802 (.O(n2377), 
	.B2(n276), 
	.B1(\ram[112][3] ), 
	.A2(n11), 
	.A1(n148));
   AO22CHD U3803 (.O(n2378), 
	.B2(n276), 
	.B1(\ram[112][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n148));
   AO22CHD U3804 (.O(n2379), 
	.B2(n276), 
	.B1(\ram[112][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n148));
   AO22CHD U3805 (.O(n2380), 
	.B2(n276), 
	.B1(\ram[112][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n148));
   AO22CHD U3806 (.O(n2381), 
	.B2(n276), 
	.B1(\ram[112][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n148));
   AO22CHD U3807 (.O(n2382), 
	.B2(n276), 
	.B1(\ram[112][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n148));
   AO22CHD U3808 (.O(n2383), 
	.B2(n276), 
	.B1(\ram[112][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n148));
   AO22CHD U3809 (.O(n2384), 
	.B2(n276), 
	.B1(\ram[112][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n148));
   AO22CHD U3810 (.O(n2385), 
	.B2(n276), 
	.B1(\ram[112][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n148));
   AO22CHD U3811 (.O(n2386), 
	.B2(n276), 
	.B1(\ram[112][12] ), 
	.A2(n20), 
	.A1(n148));
   AO22CHD U3812 (.O(n2387), 
	.B2(n276), 
	.B1(\ram[112][13] ), 
	.A2(n21), 
	.A1(n148));
   AO22CHD U3813 (.O(n2388), 
	.B2(n276), 
	.B1(\ram[112][14] ), 
	.A2(n22), 
	.A1(n148));
   AO22CHD U3814 (.O(n2389), 
	.B2(n276), 
	.B1(\ram[112][15] ), 
	.A2(n23), 
	.A1(n148));
   AO22CHD U3815 (.O(n2390), 
	.B2(n279), 
	.B1(\ram[113][0] ), 
	.A2(n6), 
	.A1(n150));
   AO22CHD U3816 (.O(n2391), 
	.B2(n279), 
	.B1(\ram[113][1] ), 
	.A2(n9), 
	.A1(n150));
   AO22CHD U3817 (.O(n2392), 
	.B2(n279), 
	.B1(\ram[113][2] ), 
	.A2(n10), 
	.A1(n150));
   AO22CHD U3818 (.O(n2393), 
	.B2(n279), 
	.B1(\ram[113][3] ), 
	.A2(n11), 
	.A1(n150));
   AO22CHD U3819 (.O(n2394), 
	.B2(n279), 
	.B1(\ram[113][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n150));
   AO22CHD U3820 (.O(n2395), 
	.B2(n279), 
	.B1(\ram[113][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n150));
   AO22CHD U3821 (.O(n2396), 
	.B2(n279), 
	.B1(\ram[113][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n150));
   AO22CHD U3822 (.O(n2397), 
	.B2(n279), 
	.B1(\ram[113][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n150));
   AO22CHD U3823 (.O(n2398), 
	.B2(n279), 
	.B1(\ram[113][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n150));
   AO22CHD U3824 (.O(n2399), 
	.B2(n279), 
	.B1(\ram[113][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n150));
   AO22CHD U3825 (.O(n2400), 
	.B2(n279), 
	.B1(\ram[113][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n150));
   AO22CHD U3826 (.O(n2401), 
	.B2(n279), 
	.B1(\ram[113][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n150));
   AO22CHD U3827 (.O(n2402), 
	.B2(n279), 
	.B1(\ram[113][12] ), 
	.A2(n20), 
	.A1(n150));
   AO22CHD U3828 (.O(n2403), 
	.B2(n279), 
	.B1(\ram[113][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n150));
   AO22CHD U3829 (.O(n2404), 
	.B2(n279), 
	.B1(\ram[113][14] ), 
	.A2(n22), 
	.A1(n150));
   AO22CHD U3830 (.O(n2405), 
	.B2(n279), 
	.B1(\ram[113][15] ), 
	.A2(n23), 
	.A1(n150));
   AO22CHD U3831 (.O(n2406), 
	.B2(n281), 
	.B1(\ram[114][0] ), 
	.A2(n6), 
	.A1(n152));
   AO22CHD U3832 (.O(n2407), 
	.B2(n281), 
	.B1(\ram[114][1] ), 
	.A2(n9), 
	.A1(n152));
   AO22CHD U3833 (.O(n2408), 
	.B2(n281), 
	.B1(\ram[114][2] ), 
	.A2(n10), 
	.A1(n152));
   AO22CHD U3834 (.O(n2409), 
	.B2(n281), 
	.B1(\ram[114][3] ), 
	.A2(n11), 
	.A1(n152));
   AO22CHD U3835 (.O(n2410), 
	.B2(n281), 
	.B1(\ram[114][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n152));
   AO22CHD U3836 (.O(n2411), 
	.B2(n281), 
	.B1(\ram[114][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n152));
   AO22CHD U3837 (.O(n2412), 
	.B2(n281), 
	.B1(\ram[114][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n152));
   AO22CHD U3838 (.O(n2413), 
	.B2(n281), 
	.B1(\ram[114][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n152));
   AO22CHD U3839 (.O(n2414), 
	.B2(n281), 
	.B1(\ram[114][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n152));
   AO22CHD U3840 (.O(n2415), 
	.B2(n281), 
	.B1(\ram[114][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n152));
   AO22CHD U3841 (.O(n2416), 
	.B2(n281), 
	.B1(\ram[114][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n152));
   AO22CHD U3842 (.O(FE_PHN7462_n2417), 
	.B2(n281), 
	.B1(\ram[114][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n152));
   AO22CHD U3843 (.O(n2418), 
	.B2(n281), 
	.B1(\ram[114][12] ), 
	.A2(n20), 
	.A1(n152));
   AO22CHD U3844 (.O(n2419), 
	.B2(n281), 
	.B1(\ram[114][13] ), 
	.A2(n21), 
	.A1(n152));
   AO22CHD U3845 (.O(n2420), 
	.B2(n281), 
	.B1(\ram[114][14] ), 
	.A2(n22), 
	.A1(n152));
   AO22CHD U3846 (.O(n2421), 
	.B2(n281), 
	.B1(\ram[114][15] ), 
	.A2(n23), 
	.A1(n152));
   AO22CHD U3847 (.O(n2422), 
	.B2(n283), 
	.B1(\ram[115][0] ), 
	.A2(n6), 
	.A1(n154));
   AO22CHD U3848 (.O(n2423), 
	.B2(n283), 
	.B1(\ram[115][1] ), 
	.A2(n9), 
	.A1(n154));
   AO22CHD U3849 (.O(n2424), 
	.B2(n283), 
	.B1(\ram[115][2] ), 
	.A2(n10), 
	.A1(n154));
   AO22CHD U3850 (.O(n2425), 
	.B2(n283), 
	.B1(\ram[115][3] ), 
	.A2(n11), 
	.A1(n154));
   AO22CHD U3851 (.O(n2426), 
	.B2(n283), 
	.B1(\ram[115][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n154));
   AO22CHD U3852 (.O(n2427), 
	.B2(n283), 
	.B1(\ram[115][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n154));
   AO22CHD U3853 (.O(n2428), 
	.B2(n283), 
	.B1(\ram[115][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n154));
   AO22CHD U3854 (.O(n2429), 
	.B2(n283), 
	.B1(\ram[115][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n154));
   AO22CHD U3855 (.O(n2430), 
	.B2(n283), 
	.B1(\ram[115][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n154));
   AO22CHD U3856 (.O(n2431), 
	.B2(n283), 
	.B1(\ram[115][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n154));
   AO22CHD U3857 (.O(n2432), 
	.B2(n283), 
	.B1(\ram[115][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n154));
   AO22CHD U3858 (.O(n2433), 
	.B2(n283), 
	.B1(\ram[115][11] ), 
	.A2(FE_OFN76_n19), 
	.A1(n154));
   AO22CHD U3859 (.O(n2434), 
	.B2(n283), 
	.B1(\ram[115][12] ), 
	.A2(n20), 
	.A1(n154));
   AO22CHD U3860 (.O(n2435), 
	.B2(n283), 
	.B1(\ram[115][13] ), 
	.A2(n21), 
	.A1(n154));
   AO22CHD U3861 (.O(n2436), 
	.B2(n283), 
	.B1(\ram[115][14] ), 
	.A2(n22), 
	.A1(n154));
   AO22CHD U3862 (.O(n2437), 
	.B2(n283), 
	.B1(\ram[115][15] ), 
	.A2(n23), 
	.A1(n154));
   AO22CHD U3863 (.O(n2438), 
	.B2(n285), 
	.B1(\ram[116][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n156));
   AO22CHD U3864 (.O(n2439), 
	.B2(n285), 
	.B1(\ram[116][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n156));
   AO22CHD U3865 (.O(n2440), 
	.B2(n285), 
	.B1(\ram[116][2] ), 
	.A2(n10), 
	.A1(n156));
   AO22CHD U3866 (.O(n2441), 
	.B2(n285), 
	.B1(\ram[116][3] ), 
	.A2(n11), 
	.A1(n156));
   AO22CHD U3867 (.O(n2442), 
	.B2(n285), 
	.B1(\ram[116][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n156));
   AO22CHD U3868 (.O(n2443), 
	.B2(n285), 
	.B1(\ram[116][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n156));
   AO22CHD U3869 (.O(n2444), 
	.B2(n285), 
	.B1(\ram[116][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n156));
   AO22CHD U3870 (.O(n2445), 
	.B2(n285), 
	.B1(\ram[116][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n156));
   AO22CHD U3871 (.O(n2446), 
	.B2(n285), 
	.B1(\ram[116][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n156));
   AO22CHD U3872 (.O(n2447), 
	.B2(n285), 
	.B1(\ram[116][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n156));
   AO22CHD U3873 (.O(n2448), 
	.B2(n285), 
	.B1(\ram[116][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n156));
   AO22CHD U3874 (.O(n2449), 
	.B2(n285), 
	.B1(\ram[116][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n156));
   AO22CHD U3875 (.O(n2450), 
	.B2(n285), 
	.B1(\ram[116][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n156));
   AO22CHD U3876 (.O(n2451), 
	.B2(n285), 
	.B1(\ram[116][13] ), 
	.A2(n21), 
	.A1(n156));
   AO22CHD U3877 (.O(n2452), 
	.B2(n285), 
	.B1(\ram[116][14] ), 
	.A2(n22), 
	.A1(n156));
   AO22CHD U3878 (.O(n2453), 
	.B2(n285), 
	.B1(\ram[116][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n156));
   AO22CHD U3879 (.O(n2454), 
	.B2(n287), 
	.B1(\ram[117][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n158));
   AO22CHD U3880 (.O(n2455), 
	.B2(n287), 
	.B1(\ram[117][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n158));
   AO22CHD U3881 (.O(n2456), 
	.B2(n287), 
	.B1(\ram[117][2] ), 
	.A2(n10), 
	.A1(n158));
   AO22CHD U3882 (.O(n2457), 
	.B2(n287), 
	.B1(\ram[117][3] ), 
	.A2(n11), 
	.A1(n158));
   AO22CHD U3883 (.O(n2458), 
	.B2(n287), 
	.B1(\ram[117][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n158));
   AO22CHD U3884 (.O(n2459), 
	.B2(n287), 
	.B1(\ram[117][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n158));
   AO22CHD U3885 (.O(n2460), 
	.B2(n287), 
	.B1(FE_PHN1720_ram_117__6_), 
	.A2(FE_OFN59_n14), 
	.A1(n158));
   AO22CHD U3886 (.O(n2461), 
	.B2(n287), 
	.B1(\ram[117][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n158));
   AO22CHD U3887 (.O(n2462), 
	.B2(n287), 
	.B1(\ram[117][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n158));
   AO22CHD U3888 (.O(n2463), 
	.B2(n287), 
	.B1(\ram[117][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n158));
   AO22CHD U3889 (.O(n2464), 
	.B2(n287), 
	.B1(\ram[117][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n158));
   AO22CHD U3890 (.O(n2465), 
	.B2(n287), 
	.B1(\ram[117][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n158));
   AO22CHD U3891 (.O(n2466), 
	.B2(n287), 
	.B1(\ram[117][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n158));
   AO22CHD U3892 (.O(n2467), 
	.B2(n287), 
	.B1(\ram[117][13] ), 
	.A2(n21), 
	.A1(n158));
   AO22CHD U3893 (.O(n2468), 
	.B2(n287), 
	.B1(\ram[117][14] ), 
	.A2(n22), 
	.A1(n158));
   AO22CHD U3894 (.O(n2469), 
	.B2(n287), 
	.B1(\ram[117][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n158));
   AO22CHD U3895 (.O(n2470), 
	.B2(n289), 
	.B1(\ram[118][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n160));
   AO22CHD U3896 (.O(n2471), 
	.B2(n289), 
	.B1(\ram[118][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n160));
   AO22CHD U3897 (.O(n2472), 
	.B2(n289), 
	.B1(\ram[118][2] ), 
	.A2(n10), 
	.A1(n160));
   AO22CHD U3898 (.O(n2473), 
	.B2(n289), 
	.B1(\ram[118][3] ), 
	.A2(n11), 
	.A1(n160));
   AO22CHD U3899 (.O(n2474), 
	.B2(n289), 
	.B1(\ram[118][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n160));
   AO22CHD U3900 (.O(n2475), 
	.B2(n289), 
	.B1(\ram[118][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n160));
   AO22CHD U3901 (.O(n2476), 
	.B2(n289), 
	.B1(\ram[118][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n160));
   AO22CHD U3902 (.O(n2477), 
	.B2(n289), 
	.B1(\ram[118][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n160));
   AO22CHD U3903 (.O(n2478), 
	.B2(n289), 
	.B1(\ram[118][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n160));
   AO22CHD U3904 (.O(n2479), 
	.B2(n289), 
	.B1(\ram[118][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n160));
   AO22CHD U3905 (.O(n2480), 
	.B2(n289), 
	.B1(\ram[118][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n160));
   AO22CHD U3906 (.O(n2481), 
	.B2(n289), 
	.B1(\ram[118][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n160));
   AO22CHD U3907 (.O(n2482), 
	.B2(n289), 
	.B1(\ram[118][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n160));
   AO22CHD U3908 (.O(n2483), 
	.B2(n289), 
	.B1(\ram[118][13] ), 
	.A2(n21), 
	.A1(n160));
   AO22CHD U3909 (.O(n2484), 
	.B2(n289), 
	.B1(\ram[118][14] ), 
	.A2(n22), 
	.A1(n160));
   AO22CHD U3910 (.O(n2485), 
	.B2(n289), 
	.B1(\ram[118][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n160));
   AO22CHD U3911 (.O(n2486), 
	.B2(n291), 
	.B1(\ram[119][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n162));
   AO22CHD U3912 (.O(n2487), 
	.B2(n291), 
	.B1(\ram[119][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n162));
   AO22CHD U3913 (.O(n2488), 
	.B2(n291), 
	.B1(\ram[119][2] ), 
	.A2(n10), 
	.A1(n162));
   AO22CHD U3914 (.O(n2489), 
	.B2(n291), 
	.B1(\ram[119][3] ), 
	.A2(n11), 
	.A1(n162));
   AO22CHD U3915 (.O(n2490), 
	.B2(n291), 
	.B1(\ram[119][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n162));
   AO22CHD U3916 (.O(n2491), 
	.B2(n291), 
	.B1(\ram[119][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n162));
   AO22CHD U3917 (.O(n2492), 
	.B2(n291), 
	.B1(\ram[119][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n162));
   AO22CHD U3918 (.O(n2493), 
	.B2(n291), 
	.B1(\ram[119][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n162));
   AO22CHD U3919 (.O(n2494), 
	.B2(n291), 
	.B1(\ram[119][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n162));
   AO22CHD U3920 (.O(n2495), 
	.B2(n291), 
	.B1(\ram[119][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n162));
   AO22CHD U3921 (.O(n2496), 
	.B2(n291), 
	.B1(\ram[119][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n162));
   AO22CHD U3922 (.O(n2497), 
	.B2(n291), 
	.B1(\ram[119][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n162));
   AO22CHD U3923 (.O(n2498), 
	.B2(n291), 
	.B1(\ram[119][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n162));
   AO22CHD U3924 (.O(n2499), 
	.B2(n291), 
	.B1(\ram[119][13] ), 
	.A2(n21), 
	.A1(n162));
   AO22CHD U3925 (.O(n2500), 
	.B2(n291), 
	.B1(\ram[119][14] ), 
	.A2(n22), 
	.A1(n162));
   AO22CHD U3926 (.O(n2501), 
	.B2(n291), 
	.B1(\ram[119][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n162));
   AO22CHD U3927 (.O(n2502), 
	.B2(n293), 
	.B1(\ram[120][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n164));
   AO22CHD U3928 (.O(n2503), 
	.B2(n293), 
	.B1(\ram[120][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n164));
   AO22CHD U3929 (.O(n2504), 
	.B2(n293), 
	.B1(\ram[120][2] ), 
	.A2(n10), 
	.A1(n164));
   AO22CHD U3930 (.O(n2505), 
	.B2(n293), 
	.B1(\ram[120][3] ), 
	.A2(n11), 
	.A1(n164));
   AO22CHD U3931 (.O(n2506), 
	.B2(n293), 
	.B1(\ram[120][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n164));
   AO22CHD U3932 (.O(n2507), 
	.B2(n293), 
	.B1(\ram[120][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n164));
   AO22CHD U3933 (.O(n2508), 
	.B2(n293), 
	.B1(\ram[120][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n164));
   AO22CHD U3934 (.O(n2509), 
	.B2(n293), 
	.B1(\ram[120][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n164));
   AO22CHD U3935 (.O(n2510), 
	.B2(n293), 
	.B1(\ram[120][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n164));
   AO22CHD U3936 (.O(n2511), 
	.B2(n293), 
	.B1(\ram[120][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n164));
   AO22CHD U3937 (.O(n2512), 
	.B2(n293), 
	.B1(\ram[120][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n164));
   AO22CHD U3938 (.O(n2513), 
	.B2(n293), 
	.B1(\ram[120][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n164));
   AO22CHD U3939 (.O(n2514), 
	.B2(n293), 
	.B1(\ram[120][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n164));
   AO22CHD U3940 (.O(n2515), 
	.B2(n293), 
	.B1(\ram[120][13] ), 
	.A2(n21), 
	.A1(n164));
   AO22CHD U3941 (.O(n2516), 
	.B2(n293), 
	.B1(FE_PHN2828_ram_120__14_), 
	.A2(n22), 
	.A1(n164));
   AO22CHD U3942 (.O(n2517), 
	.B2(n293), 
	.B1(\ram[120][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n164));
   AO22CHD U3943 (.O(n2518), 
	.B2(n295), 
	.B1(\ram[121][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n166));
   AO22CHD U3944 (.O(n2519), 
	.B2(n295), 
	.B1(\ram[121][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n166));
   AO22CHD U3945 (.O(n2520), 
	.B2(n295), 
	.B1(\ram[121][2] ), 
	.A2(n10), 
	.A1(n166));
   AO22CHD U3946 (.O(n2521), 
	.B2(n295), 
	.B1(\ram[121][3] ), 
	.A2(n11), 
	.A1(n166));
   AO22CHD U3947 (.O(n2522), 
	.B2(n295), 
	.B1(\ram[121][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n166));
   AO22CHD U3948 (.O(n2523), 
	.B2(n295), 
	.B1(\ram[121][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n166));
   AO22CHD U3949 (.O(n2524), 
	.B2(n295), 
	.B1(\ram[121][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n166));
   AO22CHD U3950 (.O(n2525), 
	.B2(n295), 
	.B1(\ram[121][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n166));
   AO22CHD U3951 (.O(n2526), 
	.B2(n295), 
	.B1(\ram[121][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n166));
   AO22CHD U3952 (.O(n2527), 
	.B2(n295), 
	.B1(\ram[121][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n166));
   AO22CHD U3953 (.O(n2528), 
	.B2(n295), 
	.B1(\ram[121][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n166));
   AO22CHD U3954 (.O(n2529), 
	.B2(n295), 
	.B1(\ram[121][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n166));
   AO22CHD U3955 (.O(n2530), 
	.B2(n295), 
	.B1(\ram[121][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n166));
   AO22CHD U3956 (.O(n2531), 
	.B2(n295), 
	.B1(\ram[121][13] ), 
	.A2(n21), 
	.A1(n166));
   AO22CHD U3957 (.O(n2532), 
	.B2(n295), 
	.B1(\ram[121][14] ), 
	.A2(n22), 
	.A1(n166));
   AO22CHD U3958 (.O(n2533), 
	.B2(n295), 
	.B1(\ram[121][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n166));
   AO22CHD U3959 (.O(n2534), 
	.B2(n297), 
	.B1(\ram[122][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n168));
   AO22CHD U3960 (.O(n2535), 
	.B2(n297), 
	.B1(\ram[122][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n168));
   AO22CHD U3961 (.O(n2536), 
	.B2(n297), 
	.B1(FE_PHN1470_ram_122__2_), 
	.A2(n10), 
	.A1(n168));
   AO22CHD U3962 (.O(n2537), 
	.B2(n297), 
	.B1(\ram[122][3] ), 
	.A2(n11), 
	.A1(n168));
   AO22CHD U3963 (.O(n2538), 
	.B2(n297), 
	.B1(\ram[122][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n168));
   AO22CHD U3964 (.O(n2539), 
	.B2(n297), 
	.B1(\ram[122][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n168));
   AO22CHD U3965 (.O(n2540), 
	.B2(n297), 
	.B1(\ram[122][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n168));
   AO22CHD U3966 (.O(n2541), 
	.B2(n297), 
	.B1(\ram[122][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n168));
   AO22CHD U3967 (.O(n2542), 
	.B2(n297), 
	.B1(\ram[122][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n168));
   AO22CHD U3968 (.O(n2543), 
	.B2(n297), 
	.B1(\ram[122][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n168));
   AO22CHD U3969 (.O(n2544), 
	.B2(n297), 
	.B1(\ram[122][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n168));
   AO22CHD U3970 (.O(n2545), 
	.B2(n297), 
	.B1(\ram[122][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n168));
   AO22CHD U3971 (.O(n2546), 
	.B2(n297), 
	.B1(\ram[122][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n168));
   AO22CHD U3972 (.O(n2547), 
	.B2(n297), 
	.B1(\ram[122][13] ), 
	.A2(n21), 
	.A1(n168));
   AO22CHD U3973 (.O(n2548), 
	.B2(n297), 
	.B1(\ram[122][14] ), 
	.A2(n22), 
	.A1(n168));
   AO22CHD U3974 (.O(n2549), 
	.B2(n297), 
	.B1(\ram[122][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n168));
   AO22CHD U3975 (.O(n2550), 
	.B2(n299), 
	.B1(\ram[123][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n170));
   AO22CHD U3976 (.O(n2551), 
	.B2(n299), 
	.B1(\ram[123][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n170));
   AO22CHD U3977 (.O(n2552), 
	.B2(n299), 
	.B1(\ram[123][2] ), 
	.A2(n10), 
	.A1(n170));
   AO22CHD U3978 (.O(n2553), 
	.B2(n299), 
	.B1(\ram[123][3] ), 
	.A2(n11), 
	.A1(n170));
   AO22CHD U3979 (.O(n2554), 
	.B2(n299), 
	.B1(\ram[123][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n170));
   AO22CHD U3980 (.O(n2555), 
	.B2(n299), 
	.B1(\ram[123][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n170));
   AO22CHD U3981 (.O(n2556), 
	.B2(n299), 
	.B1(\ram[123][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n170));
   AO22CHD U3982 (.O(n2557), 
	.B2(n299), 
	.B1(\ram[123][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n170));
   AO22CHD U3983 (.O(n2558), 
	.B2(n299), 
	.B1(\ram[123][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n170));
   AO22CHD U3984 (.O(n2559), 
	.B2(n299), 
	.B1(\ram[123][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n170));
   AO22CHD U3985 (.O(n2560), 
	.B2(n299), 
	.B1(\ram[123][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n170));
   AO22CHD U3986 (.O(n2561), 
	.B2(n299), 
	.B1(\ram[123][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n170));
   AO22CHD U3987 (.O(n2562), 
	.B2(n299), 
	.B1(\ram[123][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n170));
   AO22CHD U3988 (.O(n2563), 
	.B2(n299), 
	.B1(\ram[123][13] ), 
	.A2(n21), 
	.A1(n170));
   AO22CHD U3989 (.O(n2564), 
	.B2(n299), 
	.B1(\ram[123][14] ), 
	.A2(n22), 
	.A1(n170));
   AO22CHD U3990 (.O(n2565), 
	.B2(n299), 
	.B1(\ram[123][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n170));
   AO22CHD U3991 (.O(n2566), 
	.B2(n301), 
	.B1(\ram[124][0] ), 
	.A2(n6), 
	.A1(n172));
   AO22CHD U3992 (.O(n2567), 
	.B2(n301), 
	.B1(\ram[124][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n172));
   AO22CHD U3993 (.O(n2568), 
	.B2(n301), 
	.B1(\ram[124][2] ), 
	.A2(n10), 
	.A1(n172));
   AO22CHD U3994 (.O(n2569), 
	.B2(n301), 
	.B1(\ram[124][3] ), 
	.A2(n11), 
	.A1(n172));
   AO22CHD U3995 (.O(n2570), 
	.B2(n301), 
	.B1(\ram[124][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n172));
   AO22CHD U3996 (.O(n2571), 
	.B2(n301), 
	.B1(\ram[124][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n172));
   AO22CHD U3997 (.O(n2572), 
	.B2(n301), 
	.B1(\ram[124][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n172));
   AO22CHD U3998 (.O(n2573), 
	.B2(n301), 
	.B1(\ram[124][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n172));
   AO22CHD U3999 (.O(n2574), 
	.B2(n301), 
	.B1(\ram[124][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n172));
   AO22CHD U4000 (.O(n2575), 
	.B2(n301), 
	.B1(\ram[124][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n172));
   AO22CHD U4001 (.O(n2576), 
	.B2(n301), 
	.B1(\ram[124][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n172));
   AO22CHD U4002 (.O(n2577), 
	.B2(n301), 
	.B1(\ram[124][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n172));
   AO22CHD U4003 (.O(n2578), 
	.B2(n301), 
	.B1(\ram[124][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n172));
   AO22CHD U4004 (.O(n2579), 
	.B2(n301), 
	.B1(\ram[124][13] ), 
	.A2(n21), 
	.A1(n172));
   AO22CHD U4005 (.O(n2580), 
	.B2(n301), 
	.B1(\ram[124][14] ), 
	.A2(n22), 
	.A1(n172));
   AO22CHD U4006 (.O(n2581), 
	.B2(n301), 
	.B1(\ram[124][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n172));
   AO22CHD U4007 (.O(FE_PHN7461_n2582), 
	.B2(n303), 
	.B1(\ram[125][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n175));
   AO22CHD U4008 (.O(n2583), 
	.B2(n303), 
	.B1(\ram[125][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n175));
   AO22CHD U4009 (.O(n2584), 
	.B2(n303), 
	.B1(\ram[125][2] ), 
	.A2(n10), 
	.A1(n175));
   AO22CHD U4010 (.O(n2585), 
	.B2(n303), 
	.B1(\ram[125][3] ), 
	.A2(n11), 
	.A1(n175));
   AO22CHD U4011 (.O(n2586), 
	.B2(n303), 
	.B1(\ram[125][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n175));
   AO22CHD U4012 (.O(n2587), 
	.B2(n303), 
	.B1(\ram[125][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n175));
   AO22CHD U4013 (.O(n2588), 
	.B2(n303), 
	.B1(\ram[125][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n175));
   AO22CHD U4014 (.O(n2589), 
	.B2(n303), 
	.B1(\ram[125][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n175));
   AO22CHD U4015 (.O(n2590), 
	.B2(n303), 
	.B1(\ram[125][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n175));
   AO22CHD U4016 (.O(n2591), 
	.B2(n303), 
	.B1(\ram[125][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n175));
   AO22CHD U4017 (.O(n2592), 
	.B2(n303), 
	.B1(\ram[125][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n175));
   AO22CHD U4018 (.O(n2593), 
	.B2(n303), 
	.B1(\ram[125][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n175));
   AO22CHD U4019 (.O(n2594), 
	.B2(n303), 
	.B1(\ram[125][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n175));
   AO22CHD U4020 (.O(n2595), 
	.B2(n303), 
	.B1(\ram[125][13] ), 
	.A2(n21), 
	.A1(n175));
   AO22CHD U4021 (.O(n2596), 
	.B2(n303), 
	.B1(\ram[125][14] ), 
	.A2(n22), 
	.A1(n175));
   AO22CHD U4022 (.O(n2597), 
	.B2(n303), 
	.B1(\ram[125][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n175));
   AO22CHD U4023 (.O(n2598), 
	.B2(n305), 
	.B1(\ram[126][0] ), 
	.A2(FE_OFN41_n6), 
	.A1(n177));
   AO22CHD U4024 (.O(n2599), 
	.B2(n305), 
	.B1(\ram[126][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n177));
   AO22CHD U4025 (.O(n2600), 
	.B2(n305), 
	.B1(\ram[126][2] ), 
	.A2(n10), 
	.A1(n177));
   AO22CHD U4026 (.O(n2601), 
	.B2(n305), 
	.B1(\ram[126][3] ), 
	.A2(n11), 
	.A1(n177));
   AO22CHD U4027 (.O(n2602), 
	.B2(n305), 
	.B1(\ram[126][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n177));
   AO22CHD U4028 (.O(n2603), 
	.B2(n305), 
	.B1(\ram[126][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n177));
   AO22CHD U4029 (.O(n2604), 
	.B2(n305), 
	.B1(\ram[126][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n177));
   AO22CHD U4030 (.O(n2605), 
	.B2(n305), 
	.B1(\ram[126][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n177));
   AO22CHD U4031 (.O(n2606), 
	.B2(n305), 
	.B1(\ram[126][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n177));
   AO22CHD U4032 (.O(n2607), 
	.B2(n305), 
	.B1(\ram[126][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n177));
   AO22CHD U4033 (.O(n2608), 
	.B2(n305), 
	.B1(\ram[126][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n177));
   AO22CHD U4034 (.O(n2609), 
	.B2(n305), 
	.B1(\ram[126][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n177));
   AO22CHD U4035 (.O(n2610), 
	.B2(n305), 
	.B1(\ram[126][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n177));
   AO22CHD U4036 (.O(n2611), 
	.B2(n305), 
	.B1(\ram[126][13] ), 
	.A2(n21), 
	.A1(n177));
   AO22CHD U4037 (.O(n2612), 
	.B2(n305), 
	.B1(\ram[126][14] ), 
	.A2(n22), 
	.A1(n177));
   AO22CHD U4038 (.O(n2613), 
	.B2(n305), 
	.B1(\ram[126][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n177));
   AO22CHD U4039 (.O(n2614), 
	.B2(n307), 
	.B1(\ram[127][0] ), 
	.A2(n6), 
	.A1(n178));
   AO22CHD U4040 (.O(n2615), 
	.B2(n307), 
	.B1(\ram[127][1] ), 
	.A2(FE_OFN44_n9), 
	.A1(n178));
   AO22CHD U4041 (.O(n2616), 
	.B2(n307), 
	.B1(\ram[127][2] ), 
	.A2(n10), 
	.A1(n178));
   AO22CHD U4042 (.O(n2617), 
	.B2(n307), 
	.B1(\ram[127][3] ), 
	.A2(n11), 
	.A1(n178));
   AO22CHD U4043 (.O(n2618), 
	.B2(n307), 
	.B1(\ram[127][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n178));
   AO22CHD U4044 (.O(n2619), 
	.B2(n307), 
	.B1(\ram[127][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n178));
   AO22CHD U4045 (.O(n2620), 
	.B2(n307), 
	.B1(\ram[127][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n178));
   AO22CHD U4046 (.O(n2621), 
	.B2(n307), 
	.B1(\ram[127][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n178));
   AO22CHD U4047 (.O(n2622), 
	.B2(n307), 
	.B1(\ram[127][8] ), 
	.A2(FE_OFN69_n16), 
	.A1(n178));
   AO22CHD U4048 (.O(n2623), 
	.B2(n307), 
	.B1(\ram[127][9] ), 
	.A2(FE_OFN70_n17), 
	.A1(n178));
   AO22CHD U4049 (.O(n2624), 
	.B2(n307), 
	.B1(\ram[127][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n178));
   AO22CHD U4050 (.O(n2625), 
	.B2(n307), 
	.B1(\ram[127][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n178));
   AO22CHD U4051 (.O(n2626), 
	.B2(n307), 
	.B1(\ram[127][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n178));
   AO22CHD U4052 (.O(n2627), 
	.B2(n307), 
	.B1(\ram[127][13] ), 
	.A2(n21), 
	.A1(n178));
   AO22CHD U4053 (.O(n2628), 
	.B2(n307), 
	.B1(\ram[127][14] ), 
	.A2(n22), 
	.A1(n178));
   AO22CHD U4054 (.O(n2629), 
	.B2(n307), 
	.B1(\ram[127][15] ), 
	.A2(FE_OFN89_n23), 
	.A1(n178));
   AO22CHD U4055 (.O(n2630), 
	.B2(n309), 
	.B1(\ram[128][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n180));
   AO22CHD U4056 (.O(n2631), 
	.B2(n309), 
	.B1(\ram[128][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n180));
   AO22CHD U4057 (.O(n2632), 
	.B2(n309), 
	.B1(\ram[128][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n180));
   AO22CHD U4058 (.O(n2633), 
	.B2(n309), 
	.B1(\ram[128][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n180));
   AO22CHD U4059 (.O(n2634), 
	.B2(n309), 
	.B1(\ram[128][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n180));
   AO22CHD U4060 (.O(n2635), 
	.B2(n309), 
	.B1(\ram[128][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n180));
   AO22CHD U4061 (.O(n2636), 
	.B2(n309), 
	.B1(\ram[128][6] ), 
	.A2(n14), 
	.A1(n180));
   AO22CHD U4062 (.O(n2637), 
	.B2(n309), 
	.B1(\ram[128][7] ), 
	.A2(n15), 
	.A1(n180));
   AO22CHD U4063 (.O(n2638), 
	.B2(n309), 
	.B1(\ram[128][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n180));
   AO22CHD U4064 (.O(n2639), 
	.B2(n309), 
	.B1(\ram[128][9] ), 
	.A2(n17), 
	.A1(n180));
   AO22CHD U4065 (.O(n2640), 
	.B2(n309), 
	.B1(\ram[128][10] ), 
	.A2(n18), 
	.A1(n180));
   AO22CHD U4066 (.O(n2641), 
	.B2(n309), 
	.B1(\ram[128][11] ), 
	.A2(n19), 
	.A1(n180));
   AO22CHD U4067 (.O(n2642), 
	.B2(n309), 
	.B1(\ram[128][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n180));
   AO22CHD U4068 (.O(n2643), 
	.B2(n309), 
	.B1(\ram[128][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n180));
   AO22CHD U4069 (.O(n2644), 
	.B2(n309), 
	.B1(\ram[128][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n180));
   AO22CHD U4070 (.O(n2645), 
	.B2(n309), 
	.B1(\ram[128][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n180));
   AO22CHD U4071 (.O(n2646), 
	.B2(n312), 
	.B1(\ram[129][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n182));
   AO22CHD U4072 (.O(n2647), 
	.B2(n312), 
	.B1(\ram[129][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n182));
   AO22CHD U4073 (.O(n2648), 
	.B2(n312), 
	.B1(\ram[129][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n182));
   AO22CHD U4074 (.O(n2649), 
	.B2(n312), 
	.B1(\ram[129][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n182));
   AO22CHD U4075 (.O(n2650), 
	.B2(n312), 
	.B1(\ram[129][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n182));
   AO22CHD U4076 (.O(n2651), 
	.B2(n312), 
	.B1(\ram[129][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n182));
   AO22CHD U4077 (.O(n2652), 
	.B2(n312), 
	.B1(\ram[129][6] ), 
	.A2(n14), 
	.A1(n182));
   AO22CHD U4078 (.O(n2653), 
	.B2(n312), 
	.B1(FE_PHN1322_ram_129__7_), 
	.A2(n15), 
	.A1(n182));
   AO22CHD U4079 (.O(n2654), 
	.B2(n312), 
	.B1(\ram[129][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n182));
   AO22CHD U4080 (.O(n2655), 
	.B2(n312), 
	.B1(\ram[129][9] ), 
	.A2(n17), 
	.A1(n182));
   AO22CHD U4081 (.O(n2656), 
	.B2(n312), 
	.B1(\ram[129][10] ), 
	.A2(n18), 
	.A1(n182));
   AO22CHD U4082 (.O(n2657), 
	.B2(n312), 
	.B1(\ram[129][11] ), 
	.A2(n19), 
	.A1(n182));
   AO22CHD U4083 (.O(n2658), 
	.B2(n312), 
	.B1(\ram[129][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n182));
   AO22CHD U4084 (.O(n2659), 
	.B2(n312), 
	.B1(\ram[129][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n182));
   AO22CHD U4085 (.O(n2660), 
	.B2(n312), 
	.B1(\ram[129][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n182));
   AO22CHD U4086 (.O(n2661), 
	.B2(n312), 
	.B1(\ram[129][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n182));
   AO22CHD U4087 (.O(n2662), 
	.B2(n314), 
	.B1(\ram[130][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n184));
   AO22CHD U4088 (.O(n2663), 
	.B2(n314), 
	.B1(\ram[130][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n184));
   AO22CHD U4089 (.O(n2664), 
	.B2(n314), 
	.B1(\ram[130][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n184));
   AO22CHD U4090 (.O(n2665), 
	.B2(n314), 
	.B1(\ram[130][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n184));
   AO22CHD U4091 (.O(n2666), 
	.B2(n314), 
	.B1(\ram[130][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n184));
   AO22CHD U4092 (.O(n2667), 
	.B2(n314), 
	.B1(\ram[130][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n184));
   AO22CHD U4093 (.O(n2668), 
	.B2(n314), 
	.B1(\ram[130][6] ), 
	.A2(n14), 
	.A1(n184));
   AO22CHD U4094 (.O(n2669), 
	.B2(n314), 
	.B1(\ram[130][7] ), 
	.A2(n15), 
	.A1(n184));
   AO22CHD U4095 (.O(n2670), 
	.B2(n314), 
	.B1(\ram[130][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n184));
   AO22CHD U4096 (.O(n2671), 
	.B2(n314), 
	.B1(\ram[130][9] ), 
	.A2(n17), 
	.A1(n184));
   AO22CHD U4097 (.O(n2672), 
	.B2(n314), 
	.B1(\ram[130][10] ), 
	.A2(n18), 
	.A1(n184));
   AO22CHD U4098 (.O(n2673), 
	.B2(n314), 
	.B1(\ram[130][11] ), 
	.A2(n19), 
	.A1(n184));
   AO22CHD U4099 (.O(n2674), 
	.B2(n314), 
	.B1(\ram[130][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n184));
   AO22CHD U4100 (.O(n2675), 
	.B2(n314), 
	.B1(\ram[130][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n184));
   AO22CHD U4101 (.O(n2676), 
	.B2(n314), 
	.B1(\ram[130][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n184));
   AO22CHD U4102 (.O(n2677), 
	.B2(n314), 
	.B1(\ram[130][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n184));
   AO22CHD U4103 (.O(n2678), 
	.B2(n316), 
	.B1(\ram[131][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n186));
   AO22CHD U4104 (.O(n2679), 
	.B2(n316), 
	.B1(\ram[131][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n186));
   AO22CHD U4105 (.O(n2680), 
	.B2(n316), 
	.B1(\ram[131][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n186));
   AO22CHD U4106 (.O(n2681), 
	.B2(n316), 
	.B1(\ram[131][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n186));
   AO22CHD U4107 (.O(n2682), 
	.B2(n316), 
	.B1(\ram[131][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n186));
   AO22CHD U4108 (.O(n2683), 
	.B2(n316), 
	.B1(\ram[131][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n186));
   AO22CHD U4109 (.O(n2684), 
	.B2(n316), 
	.B1(\ram[131][6] ), 
	.A2(n14), 
	.A1(n186));
   AO22CHD U4110 (.O(n2685), 
	.B2(n316), 
	.B1(\ram[131][7] ), 
	.A2(n15), 
	.A1(n186));
   AO22CHD U4111 (.O(n2686), 
	.B2(n316), 
	.B1(\ram[131][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n186));
   AO22CHD U4112 (.O(n2687), 
	.B2(n316), 
	.B1(\ram[131][9] ), 
	.A2(n17), 
	.A1(n186));
   AO22CHD U4113 (.O(n2688), 
	.B2(n316), 
	.B1(\ram[131][10] ), 
	.A2(n18), 
	.A1(n186));
   AO22CHD U4114 (.O(n2689), 
	.B2(n316), 
	.B1(\ram[131][11] ), 
	.A2(n19), 
	.A1(n186));
   AO22CHD U4115 (.O(n2690), 
	.B2(n316), 
	.B1(\ram[131][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n186));
   AO22CHD U4116 (.O(n2691), 
	.B2(n316), 
	.B1(\ram[131][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n186));
   AO22CHD U4117 (.O(n2692), 
	.B2(n316), 
	.B1(\ram[131][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n186));
   AO22CHD U4118 (.O(n2693), 
	.B2(n316), 
	.B1(\ram[131][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n186));
   AO22CHD U4119 (.O(n2694), 
	.B2(n318), 
	.B1(\ram[132][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n188));
   AO22CHD U4120 (.O(n2695), 
	.B2(n318), 
	.B1(\ram[132][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n188));
   AO22CHD U4121 (.O(n2696), 
	.B2(n318), 
	.B1(\ram[132][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n188));
   AO22CHD U4122 (.O(n2697), 
	.B2(n318), 
	.B1(\ram[132][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n188));
   AO22CHD U4123 (.O(n2698), 
	.B2(n318), 
	.B1(\ram[132][4] ), 
	.A2(n12), 
	.A1(n188));
   AO22CHD U4124 (.O(n2699), 
	.B2(n318), 
	.B1(\ram[132][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n188));
   AO22CHD U4125 (.O(n2700), 
	.B2(n318), 
	.B1(\ram[132][6] ), 
	.A2(n14), 
	.A1(n188));
   AO22CHD U4126 (.O(n2701), 
	.B2(n318), 
	.B1(\ram[132][7] ), 
	.A2(n15), 
	.A1(n188));
   AO22CHD U4127 (.O(n2702), 
	.B2(n318), 
	.B1(FE_PHN2193_ram_132__8_), 
	.A2(FE_OFN68_n16), 
	.A1(n188));
   AO22CHD U4128 (.O(n2703), 
	.B2(n318), 
	.B1(\ram[132][9] ), 
	.A2(n17), 
	.A1(n188));
   AO22CHD U4129 (.O(n2704), 
	.B2(n318), 
	.B1(\ram[132][10] ), 
	.A2(n18), 
	.A1(n188));
   AO22CHD U4130 (.O(n2705), 
	.B2(n318), 
	.B1(\ram[132][11] ), 
	.A2(n19), 
	.A1(n188));
   AO22CHD U4131 (.O(n2706), 
	.B2(n318), 
	.B1(\ram[132][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n188));
   AO22CHD U4132 (.O(n2707), 
	.B2(n318), 
	.B1(\ram[132][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n188));
   AO22CHD U4133 (.O(n2708), 
	.B2(n318), 
	.B1(\ram[132][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n188));
   AO22CHD U4134 (.O(n2709), 
	.B2(n318), 
	.B1(\ram[132][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n188));
   AO22CHD U4135 (.O(n2710), 
	.B2(n320), 
	.B1(\ram[133][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n190));
   AO22CHD U4136 (.O(n2711), 
	.B2(n320), 
	.B1(\ram[133][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n190));
   AO22CHD U4137 (.O(n2712), 
	.B2(n320), 
	.B1(\ram[133][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n190));
   AO22CHD U4138 (.O(n2713), 
	.B2(n320), 
	.B1(\ram[133][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n190));
   AO22CHD U4139 (.O(n2714), 
	.B2(n320), 
	.B1(\ram[133][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n190));
   AO22CHD U4140 (.O(n2715), 
	.B2(n320), 
	.B1(\ram[133][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n190));
   AO22CHD U4141 (.O(n2716), 
	.B2(n320), 
	.B1(\ram[133][6] ), 
	.A2(n14), 
	.A1(n190));
   AO22CHD U4142 (.O(n2717), 
	.B2(n320), 
	.B1(\ram[133][7] ), 
	.A2(n15), 
	.A1(n190));
   AO22CHD U4143 (.O(n2718), 
	.B2(n320), 
	.B1(\ram[133][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n190));
   AO22CHD U4144 (.O(n2719), 
	.B2(n320), 
	.B1(FE_PHN5386_ram_133__9_), 
	.A2(n17), 
	.A1(n190));
   AO22CHD U4145 (.O(n2720), 
	.B2(n320), 
	.B1(\ram[133][10] ), 
	.A2(n18), 
	.A1(n190));
   AO22CHD U4146 (.O(n2721), 
	.B2(n320), 
	.B1(\ram[133][11] ), 
	.A2(n19), 
	.A1(n190));
   AO22CHD U4147 (.O(n2722), 
	.B2(n320), 
	.B1(\ram[133][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n190));
   AO22CHD U4148 (.O(n2723), 
	.B2(n320), 
	.B1(\ram[133][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n190));
   AO22CHD U4149 (.O(n2724), 
	.B2(n320), 
	.B1(\ram[133][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n190));
   AO22CHD U4150 (.O(n2725), 
	.B2(n320), 
	.B1(\ram[133][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n190));
   AO22CHD U4151 (.O(n2726), 
	.B2(n322), 
	.B1(\ram[134][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n192));
   AO22CHD U4152 (.O(n2727), 
	.B2(n322), 
	.B1(\ram[134][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n192));
   AO22CHD U4153 (.O(n2728), 
	.B2(n322), 
	.B1(\ram[134][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n192));
   AO22CHD U4154 (.O(n2729), 
	.B2(n322), 
	.B1(\ram[134][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n192));
   AO22CHD U4155 (.O(n2730), 
	.B2(n322), 
	.B1(\ram[134][4] ), 
	.A2(n12), 
	.A1(n192));
   AO22CHD U4156 (.O(n2731), 
	.B2(n322), 
	.B1(\ram[134][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n192));
   AO22CHD U4157 (.O(n2732), 
	.B2(n322), 
	.B1(\ram[134][6] ), 
	.A2(n14), 
	.A1(n192));
   AO22CHD U4158 (.O(n2733), 
	.B2(n322), 
	.B1(\ram[134][7] ), 
	.A2(n15), 
	.A1(n192));
   AO22CHD U4159 (.O(n2734), 
	.B2(n322), 
	.B1(\ram[134][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n192));
   AO22CHD U4160 (.O(n2735), 
	.B2(n322), 
	.B1(\ram[134][9] ), 
	.A2(n17), 
	.A1(n192));
   AO22CHD U4161 (.O(n2736), 
	.B2(n322), 
	.B1(\ram[134][10] ), 
	.A2(n18), 
	.A1(n192));
   AO22CHD U4162 (.O(n2737), 
	.B2(n322), 
	.B1(\ram[134][11] ), 
	.A2(n19), 
	.A1(n192));
   AO22CHD U4163 (.O(n2738), 
	.B2(n322), 
	.B1(\ram[134][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n192));
   AO22CHD U4164 (.O(n2739), 
	.B2(n322), 
	.B1(\ram[134][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n192));
   AO22CHD U4165 (.O(n2740), 
	.B2(n322), 
	.B1(\ram[134][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n192));
   AO22CHD U4166 (.O(n2741), 
	.B2(n322), 
	.B1(\ram[134][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n192));
   AO22CHD U4167 (.O(n2742), 
	.B2(n324), 
	.B1(\ram[135][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n194));
   AO22CHD U4168 (.O(n2743), 
	.B2(n324), 
	.B1(\ram[135][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n194));
   AO22CHD U4169 (.O(n2744), 
	.B2(n324), 
	.B1(\ram[135][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n194));
   AO22CHD U4170 (.O(n2745), 
	.B2(n324), 
	.B1(\ram[135][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n194));
   AO22CHD U4171 (.O(n2746), 
	.B2(n324), 
	.B1(\ram[135][4] ), 
	.A2(n12), 
	.A1(n194));
   AO22CHD U4172 (.O(n2747), 
	.B2(n324), 
	.B1(\ram[135][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n194));
   AO22CHD U4173 (.O(n2748), 
	.B2(n324), 
	.B1(\ram[135][6] ), 
	.A2(n14), 
	.A1(n194));
   AO22CHD U4174 (.O(n2749), 
	.B2(n324), 
	.B1(\ram[135][7] ), 
	.A2(n15), 
	.A1(n194));
   AO22CHD U4175 (.O(n2750), 
	.B2(n324), 
	.B1(\ram[135][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n194));
   AO22CHD U4176 (.O(n2751), 
	.B2(n324), 
	.B1(\ram[135][9] ), 
	.A2(n17), 
	.A1(n194));
   AO22CHD U4177 (.O(n2752), 
	.B2(n324), 
	.B1(\ram[135][10] ), 
	.A2(n18), 
	.A1(n194));
   AO22CHD U4178 (.O(n2753), 
	.B2(n324), 
	.B1(\ram[135][11] ), 
	.A2(n19), 
	.A1(n194));
   AO22CHD U4179 (.O(n2754), 
	.B2(n324), 
	.B1(\ram[135][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n194));
   AO22CHD U4180 (.O(n2755), 
	.B2(n324), 
	.B1(\ram[135][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n194));
   AO22CHD U4181 (.O(n2756), 
	.B2(n324), 
	.B1(\ram[135][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n194));
   AO22CHD U4182 (.O(n2757), 
	.B2(n324), 
	.B1(\ram[135][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n194));
   AO22CHD U4183 (.O(n2758), 
	.B2(n326), 
	.B1(\ram[136][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n196));
   AO22CHD U4184 (.O(n2759), 
	.B2(n326), 
	.B1(\ram[136][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n196));
   AO22CHD U4185 (.O(n2760), 
	.B2(n326), 
	.B1(\ram[136][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n196));
   AO22CHD U4186 (.O(n2761), 
	.B2(n326), 
	.B1(\ram[136][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n196));
   AO22CHD U4187 (.O(n2762), 
	.B2(n326), 
	.B1(\ram[136][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n196));
   AO22CHD U4188 (.O(n2763), 
	.B2(n326), 
	.B1(\ram[136][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n196));
   AO22CHD U4189 (.O(n2764), 
	.B2(n326), 
	.B1(\ram[136][6] ), 
	.A2(n14), 
	.A1(n196));
   AO22CHD U4190 (.O(n2765), 
	.B2(n326), 
	.B1(\ram[136][7] ), 
	.A2(n15), 
	.A1(n196));
   AO22CHD U4191 (.O(n2766), 
	.B2(n326), 
	.B1(\ram[136][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n196));
   AO22CHD U4192 (.O(n2767), 
	.B2(n326), 
	.B1(\ram[136][9] ), 
	.A2(n17), 
	.A1(n196));
   AO22CHD U4193 (.O(n2768), 
	.B2(n326), 
	.B1(\ram[136][10] ), 
	.A2(n18), 
	.A1(n196));
   AO22CHD U4194 (.O(n2769), 
	.B2(n326), 
	.B1(\ram[136][11] ), 
	.A2(n19), 
	.A1(n196));
   AO22CHD U4195 (.O(n2770), 
	.B2(n326), 
	.B1(\ram[136][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n196));
   AO22CHD U4196 (.O(n2771), 
	.B2(n326), 
	.B1(\ram[136][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n196));
   AO22CHD U4197 (.O(n2772), 
	.B2(n326), 
	.B1(\ram[136][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n196));
   AO22CHD U4198 (.O(n2773), 
	.B2(n326), 
	.B1(\ram[136][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n196));
   AO22CHD U4199 (.O(n2774), 
	.B2(n328), 
	.B1(\ram[137][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n198));
   AO22CHD U4200 (.O(n2775), 
	.B2(n328), 
	.B1(\ram[137][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n198));
   AO22CHD U4201 (.O(n2776), 
	.B2(n328), 
	.B1(\ram[137][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n198));
   AO22CHD U4202 (.O(n2777), 
	.B2(n328), 
	.B1(\ram[137][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n198));
   AO22CHD U4203 (.O(n2778), 
	.B2(n328), 
	.B1(\ram[137][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n198));
   AO22CHD U4204 (.O(n2779), 
	.B2(n328), 
	.B1(\ram[137][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n198));
   AO22CHD U4205 (.O(n2780), 
	.B2(n328), 
	.B1(\ram[137][6] ), 
	.A2(n14), 
	.A1(n198));
   AO22CHD U4206 (.O(n2781), 
	.B2(n328), 
	.B1(\ram[137][7] ), 
	.A2(n15), 
	.A1(n198));
   AO22CHD U4207 (.O(n2782), 
	.B2(n328), 
	.B1(\ram[137][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n198));
   AO22CHD U4208 (.O(n2783), 
	.B2(n328), 
	.B1(\ram[137][9] ), 
	.A2(n17), 
	.A1(n198));
   AO22CHD U4209 (.O(n2784), 
	.B2(n328), 
	.B1(\ram[137][10] ), 
	.A2(n18), 
	.A1(n198));
   AO22CHD U4210 (.O(n2785), 
	.B2(n328), 
	.B1(\ram[137][11] ), 
	.A2(n19), 
	.A1(n198));
   AO22CHD U4211 (.O(n2786), 
	.B2(n328), 
	.B1(\ram[137][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n198));
   AO22CHD U4212 (.O(n2787), 
	.B2(n328), 
	.B1(\ram[137][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n198));
   AO22CHD U4213 (.O(n2788), 
	.B2(n328), 
	.B1(\ram[137][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n198));
   AO22CHD U4214 (.O(n2789), 
	.B2(n328), 
	.B1(\ram[137][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n198));
   AO22CHD U4215 (.O(n2790), 
	.B2(n330), 
	.B1(\ram[138][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n200));
   AO22CHD U4216 (.O(n2791), 
	.B2(n330), 
	.B1(\ram[138][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n200));
   AO22CHD U4217 (.O(n2792), 
	.B2(n330), 
	.B1(\ram[138][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n200));
   AO22CHD U4218 (.O(n2793), 
	.B2(n330), 
	.B1(\ram[138][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n200));
   AO22CHD U4219 (.O(n2794), 
	.B2(n330), 
	.B1(\ram[138][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n200));
   AO22CHD U4220 (.O(n2795), 
	.B2(n330), 
	.B1(\ram[138][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n200));
   AO22CHD U4221 (.O(n2796), 
	.B2(n330), 
	.B1(\ram[138][6] ), 
	.A2(n14), 
	.A1(n200));
   AO22CHD U4222 (.O(n2797), 
	.B2(n330), 
	.B1(\ram[138][7] ), 
	.A2(n15), 
	.A1(n200));
   AO22CHD U4223 (.O(n2798), 
	.B2(n330), 
	.B1(\ram[138][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n200));
   AO22CHD U4224 (.O(n2799), 
	.B2(n330), 
	.B1(\ram[138][9] ), 
	.A2(n17), 
	.A1(n200));
   AO22CHD U4225 (.O(n2800), 
	.B2(n330), 
	.B1(\ram[138][10] ), 
	.A2(n18), 
	.A1(n200));
   AO22CHD U4226 (.O(n2801), 
	.B2(n330), 
	.B1(\ram[138][11] ), 
	.A2(n19), 
	.A1(n200));
   AO22CHD U4227 (.O(n2802), 
	.B2(n330), 
	.B1(\ram[138][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n200));
   AO22CHD U4228 (.O(n2803), 
	.B2(n330), 
	.B1(\ram[138][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n200));
   AO22CHD U4229 (.O(n2804), 
	.B2(n330), 
	.B1(\ram[138][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n200));
   AO22CHD U4230 (.O(n2805), 
	.B2(n330), 
	.B1(\ram[138][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n200));
   AO22CHD U4231 (.O(n2806), 
	.B2(n332), 
	.B1(\ram[139][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n202));
   AO22CHD U4232 (.O(n2807), 
	.B2(n332), 
	.B1(\ram[139][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n202));
   AO22CHD U4233 (.O(n2808), 
	.B2(n332), 
	.B1(\ram[139][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n202));
   AO22CHD U4234 (.O(n2809), 
	.B2(n332), 
	.B1(\ram[139][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n202));
   AO22CHD U4235 (.O(n2810), 
	.B2(n332), 
	.B1(\ram[139][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n202));
   AO22CHD U4236 (.O(n2811), 
	.B2(n332), 
	.B1(\ram[139][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n202));
   AO22CHD U4237 (.O(n2812), 
	.B2(n332), 
	.B1(\ram[139][6] ), 
	.A2(n14), 
	.A1(n202));
   AO22CHD U4238 (.O(n2813), 
	.B2(n332), 
	.B1(\ram[139][7] ), 
	.A2(n15), 
	.A1(n202));
   AO22CHD U4239 (.O(n2814), 
	.B2(n332), 
	.B1(\ram[139][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n202));
   AO22CHD U4240 (.O(n2815), 
	.B2(n332), 
	.B1(\ram[139][9] ), 
	.A2(n17), 
	.A1(n202));
   AO22CHD U4241 (.O(n2816), 
	.B2(n332), 
	.B1(\ram[139][10] ), 
	.A2(n18), 
	.A1(n202));
   AO22CHD U4242 (.O(n2817), 
	.B2(n332), 
	.B1(\ram[139][11] ), 
	.A2(n19), 
	.A1(n202));
   AO22CHD U4243 (.O(n2818), 
	.B2(n332), 
	.B1(\ram[139][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n202));
   AO22CHD U4244 (.O(n2819), 
	.B2(n332), 
	.B1(\ram[139][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n202));
   AO22CHD U4245 (.O(n2820), 
	.B2(n332), 
	.B1(\ram[139][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n202));
   AO22CHD U4246 (.O(n2821), 
	.B2(n332), 
	.B1(\ram[139][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n202));
   AO22CHD U4247 (.O(n2822), 
	.B2(n334), 
	.B1(\ram[140][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n204));
   AO22CHD U4248 (.O(n2823), 
	.B2(n334), 
	.B1(\ram[140][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n204));
   AO22CHD U4249 (.O(n2824), 
	.B2(n334), 
	.B1(\ram[140][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n204));
   AO22CHD U4250 (.O(n2825), 
	.B2(n334), 
	.B1(\ram[140][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n204));
   AO22CHD U4251 (.O(n2826), 
	.B2(n334), 
	.B1(\ram[140][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n204));
   AO22CHD U4252 (.O(n2827), 
	.B2(n334), 
	.B1(\ram[140][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n204));
   AO22CHD U4253 (.O(n2828), 
	.B2(n334), 
	.B1(\ram[140][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n204));
   AO22CHD U4254 (.O(n2829), 
	.B2(n334), 
	.B1(\ram[140][7] ), 
	.A2(n15), 
	.A1(n204));
   AO22CHD U4255 (.O(n2830), 
	.B2(n334), 
	.B1(\ram[140][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n204));
   AO22CHD U4256 (.O(n2831), 
	.B2(n334), 
	.B1(\ram[140][9] ), 
	.A2(n17), 
	.A1(n204));
   AO22CHD U4257 (.O(n2832), 
	.B2(n334), 
	.B1(\ram[140][10] ), 
	.A2(n18), 
	.A1(n204));
   AO22CHD U4258 (.O(n2833), 
	.B2(n334), 
	.B1(\ram[140][11] ), 
	.A2(n19), 
	.A1(n204));
   AO22CHD U4259 (.O(n2834), 
	.B2(n334), 
	.B1(\ram[140][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n204));
   AO22CHD U4260 (.O(n2835), 
	.B2(n334), 
	.B1(\ram[140][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n204));
   AO22CHD U4261 (.O(n2836), 
	.B2(n334), 
	.B1(\ram[140][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n204));
   AO22CHD U4262 (.O(n2837), 
	.B2(n334), 
	.B1(\ram[140][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n204));
   AO22CHD U4263 (.O(n2838), 
	.B2(n336), 
	.B1(\ram[141][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n206));
   AO22CHD U4264 (.O(n2839), 
	.B2(n336), 
	.B1(\ram[141][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n206));
   AO22CHD U4265 (.O(n2840), 
	.B2(n336), 
	.B1(\ram[141][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n206));
   AO22CHD U4266 (.O(n2841), 
	.B2(n336), 
	.B1(\ram[141][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n206));
   AO22CHD U4267 (.O(n2842), 
	.B2(n336), 
	.B1(\ram[141][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n206));
   AO22CHD U4268 (.O(n2843), 
	.B2(n336), 
	.B1(\ram[141][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n206));
   AO22CHD U4269 (.O(n2844), 
	.B2(n336), 
	.B1(\ram[141][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n206));
   AO22CHD U4270 (.O(n2845), 
	.B2(n336), 
	.B1(\ram[141][7] ), 
	.A2(n15), 
	.A1(n206));
   AO22CHD U4271 (.O(n2846), 
	.B2(n336), 
	.B1(\ram[141][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n206));
   AO22CHD U4272 (.O(n2847), 
	.B2(n336), 
	.B1(\ram[141][9] ), 
	.A2(n17), 
	.A1(n206));
   AO22CHD U4273 (.O(n2848), 
	.B2(n336), 
	.B1(\ram[141][10] ), 
	.A2(n18), 
	.A1(n206));
   AO22CHD U4274 (.O(n2849), 
	.B2(n336), 
	.B1(\ram[141][11] ), 
	.A2(n19), 
	.A1(n206));
   AO22CHD U4275 (.O(n2850), 
	.B2(n336), 
	.B1(\ram[141][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n206));
   AO22CHD U4276 (.O(n2851), 
	.B2(n336), 
	.B1(\ram[141][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n206));
   AO22CHD U4277 (.O(n2852), 
	.B2(n336), 
	.B1(\ram[141][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n206));
   AO22CHD U4278 (.O(n2853), 
	.B2(n336), 
	.B1(\ram[141][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n206));
   AO22CHD U4279 (.O(n2854), 
	.B2(n338), 
	.B1(\ram[142][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n209));
   AO22CHD U4280 (.O(n2855), 
	.B2(n338), 
	.B1(\ram[142][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n209));
   AO22CHD U4281 (.O(n2856), 
	.B2(n338), 
	.B1(\ram[142][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n209));
   AO22CHD U4282 (.O(n2857), 
	.B2(n338), 
	.B1(\ram[142][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n209));
   AO22CHD U4283 (.O(n2858), 
	.B2(n338), 
	.B1(\ram[142][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n209));
   AO22CHD U4284 (.O(n2859), 
	.B2(n338), 
	.B1(\ram[142][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n209));
   AO22CHD U4285 (.O(n2860), 
	.B2(n338), 
	.B1(\ram[142][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n209));
   AO22CHD U4286 (.O(n2861), 
	.B2(n338), 
	.B1(\ram[142][7] ), 
	.A2(n15), 
	.A1(n209));
   AO22CHD U4287 (.O(n2862), 
	.B2(n338), 
	.B1(\ram[142][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n209));
   AO22CHD U4288 (.O(n2863), 
	.B2(n338), 
	.B1(\ram[142][9] ), 
	.A2(n17), 
	.A1(n209));
   AO22CHD U4289 (.O(n2864), 
	.B2(n338), 
	.B1(\ram[142][10] ), 
	.A2(n18), 
	.A1(n209));
   AO22CHD U4290 (.O(n2865), 
	.B2(n338), 
	.B1(\ram[142][11] ), 
	.A2(n19), 
	.A1(n209));
   AO22CHD U4291 (.O(n2866), 
	.B2(n338), 
	.B1(\ram[142][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n209));
   AO22CHD U4292 (.O(n2867), 
	.B2(n338), 
	.B1(\ram[142][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n209));
   AO22CHD U4293 (.O(n2868), 
	.B2(n338), 
	.B1(\ram[142][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n209));
   AO22CHD U4294 (.O(n2869), 
	.B2(n338), 
	.B1(\ram[142][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n209));
   AO22CHD U4295 (.O(n2870), 
	.B2(n340), 
	.B1(\ram[143][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n211));
   AO22CHD U4296 (.O(n2871), 
	.B2(n340), 
	.B1(\ram[143][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n211));
   AO22CHD U4297 (.O(n2872), 
	.B2(n340), 
	.B1(\ram[143][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n211));
   AO22CHD U4298 (.O(n2873), 
	.B2(n340), 
	.B1(\ram[143][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n211));
   AO22CHD U4299 (.O(n2874), 
	.B2(n340), 
	.B1(\ram[143][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n211));
   AO22CHD U4300 (.O(n2875), 
	.B2(n340), 
	.B1(\ram[143][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n211));
   AO22CHD U4301 (.O(n2876), 
	.B2(n340), 
	.B1(\ram[143][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n211));
   AO22CHD U4302 (.O(n2877), 
	.B2(n340), 
	.B1(\ram[143][7] ), 
	.A2(n15), 
	.A1(n211));
   AO22CHD U4303 (.O(n2878), 
	.B2(n340), 
	.B1(\ram[143][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n211));
   AO22CHD U4304 (.O(n2879), 
	.B2(n340), 
	.B1(\ram[143][9] ), 
	.A2(n17), 
	.A1(n211));
   AO22CHD U4305 (.O(n2880), 
	.B2(n340), 
	.B1(FE_PHN3074_ram_143__10_), 
	.A2(n18), 
	.A1(n211));
   AO22CHD U4306 (.O(n2881), 
	.B2(n340), 
	.B1(\ram[143][11] ), 
	.A2(n19), 
	.A1(n211));
   AO22CHD U4307 (.O(n2882), 
	.B2(n340), 
	.B1(\ram[143][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n211));
   AO22CHD U4308 (.O(n2883), 
	.B2(n340), 
	.B1(\ram[143][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n211));
   AO22CHD U4309 (.O(n2884), 
	.B2(n340), 
	.B1(\ram[143][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n211));
   AO22CHD U4310 (.O(n2885), 
	.B2(n340), 
	.B1(\ram[143][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n211));
   AO22CHD U4311 (.O(n2886), 
	.B2(n343), 
	.B1(\ram[144][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n212));
   AO22CHD U4312 (.O(n2887), 
	.B2(n343), 
	.B1(\ram[144][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n212));
   AO22CHD U4313 (.O(n2888), 
	.B2(n343), 
	.B1(\ram[144][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n212));
   AO22CHD U4314 (.O(n2889), 
	.B2(n343), 
	.B1(\ram[144][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n212));
   AO22CHD U4315 (.O(FE_PHN7249_n2890), 
	.B2(n343), 
	.B1(\ram[144][4] ), 
	.A2(n12), 
	.A1(n212));
   AO22CHD U4316 (.O(n2891), 
	.B2(n343), 
	.B1(\ram[144][5] ), 
	.A2(n13), 
	.A1(n212));
   AO22CHD U4317 (.O(n2892), 
	.B2(n343), 
	.B1(\ram[144][6] ), 
	.A2(n14), 
	.A1(n212));
   AO22CHD U4318 (.O(n2893), 
	.B2(n343), 
	.B1(\ram[144][7] ), 
	.A2(n15), 
	.A1(n212));
   AO22CHD U4319 (.O(n2894), 
	.B2(n343), 
	.B1(FE_PHN4185_ram_144__8_), 
	.A2(n16), 
	.A1(n212));
   AO22CHD U4320 (.O(n2895), 
	.B2(n343), 
	.B1(\ram[144][9] ), 
	.A2(n17), 
	.A1(n212));
   AO22CHD U4321 (.O(n2896), 
	.B2(n343), 
	.B1(\ram[144][10] ), 
	.A2(n18), 
	.A1(n212));
   AO22CHD U4322 (.O(n2897), 
	.B2(n343), 
	.B1(\ram[144][11] ), 
	.A2(n19), 
	.A1(n212));
   AO22CHD U4323 (.O(n2898), 
	.B2(n343), 
	.B1(\ram[144][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n212));
   AO22CHD U4324 (.O(n2899), 
	.B2(n343), 
	.B1(\ram[144][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n212));
   AO22CHD U4325 (.O(n2900), 
	.B2(n343), 
	.B1(\ram[144][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n212));
   AO22CHD U4326 (.O(n2901), 
	.B2(n343), 
	.B1(\ram[144][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n212));
   AO22CHD U4327 (.O(n2902), 
	.B2(n346), 
	.B1(FE_PHN4161_ram_145__0_), 
	.A2(FE_OFN43_n6), 
	.A1(n214));
   AO22CHD U4328 (.O(n2903), 
	.B2(n346), 
	.B1(FE_PHN5534_ram_145__1_), 
	.A2(FE_OFN45_n9), 
	.A1(n214));
   AO22CHD U4329 (.O(n2904), 
	.B2(n346), 
	.B1(\ram[145][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n214));
   AO22CHD U4330 (.O(n2905), 
	.B2(n346), 
	.B1(\ram[145][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n214));
   AO22CHD U4331 (.O(n2906), 
	.B2(n346), 
	.B1(\ram[145][4] ), 
	.A2(n12), 
	.A1(n214));
   AO22CHD U4332 (.O(n2907), 
	.B2(n346), 
	.B1(\ram[145][5] ), 
	.A2(n13), 
	.A1(n214));
   AO22CHD U4333 (.O(n2908), 
	.B2(n346), 
	.B1(\ram[145][6] ), 
	.A2(n14), 
	.A1(n214));
   AO22CHD U4334 (.O(n2909), 
	.B2(n346), 
	.B1(FE_PHN5447_ram_145__7_), 
	.A2(n15), 
	.A1(n214));
   AO22CHD U4335 (.O(n2910), 
	.B2(n346), 
	.B1(\ram[145][8] ), 
	.A2(n16), 
	.A1(n214));
   AO22CHD U4336 (.O(n2911), 
	.B2(n346), 
	.B1(\ram[145][9] ), 
	.A2(n17), 
	.A1(n214));
   AO22CHD U4337 (.O(n2912), 
	.B2(n346), 
	.B1(FE_PHN4026_ram_145__10_), 
	.A2(n18), 
	.A1(n214));
   AO22CHD U4338 (.O(n2913), 
	.B2(n346), 
	.B1(\ram[145][11] ), 
	.A2(n19), 
	.A1(n214));
   AO22CHD U4339 (.O(n2914), 
	.B2(n346), 
	.B1(\ram[145][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n214));
   AO22CHD U4340 (.O(n2915), 
	.B2(n346), 
	.B1(\ram[145][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n214));
   AO22CHD U4341 (.O(n2916), 
	.B2(n346), 
	.B1(\ram[145][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n214));
   AO22CHD U4342 (.O(n2917), 
	.B2(n346), 
	.B1(\ram[145][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n214));
   AO22CHD U4343 (.O(n2918), 
	.B2(n348), 
	.B1(\ram[146][0] ), 
	.A2(n6), 
	.A1(n216));
   AO22CHD U4344 (.O(n2919), 
	.B2(n348), 
	.B1(\ram[146][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n216));
   AO22CHD U4345 (.O(n2920), 
	.B2(n348), 
	.B1(\ram[146][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n216));
   AO22CHD U4346 (.O(n2921), 
	.B2(n348), 
	.B1(\ram[146][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n216));
   AO22CHD U4347 (.O(n2922), 
	.B2(n348), 
	.B1(\ram[146][4] ), 
	.A2(n12), 
	.A1(n216));
   AO22CHD U4348 (.O(n2923), 
	.B2(n348), 
	.B1(\ram[146][5] ), 
	.A2(n13), 
	.A1(n216));
   AO22CHD U4349 (.O(n2924), 
	.B2(n348), 
	.B1(\ram[146][6] ), 
	.A2(n14), 
	.A1(n216));
   AO22CHD U4350 (.O(n2925), 
	.B2(n348), 
	.B1(\ram[146][7] ), 
	.A2(n15), 
	.A1(n216));
   AO22CHD U4351 (.O(n2926), 
	.B2(n348), 
	.B1(\ram[146][8] ), 
	.A2(n16), 
	.A1(n216));
   AO22CHD U4352 (.O(n2927), 
	.B2(n348), 
	.B1(\ram[146][9] ), 
	.A2(n17), 
	.A1(n216));
   AO22CHD U4353 (.O(n2928), 
	.B2(n348), 
	.B1(\ram[146][10] ), 
	.A2(n18), 
	.A1(n216));
   AO22CHD U4354 (.O(n2929), 
	.B2(n348), 
	.B1(\ram[146][11] ), 
	.A2(n19), 
	.A1(n216));
   AO22CHD U4355 (.O(n2930), 
	.B2(n348), 
	.B1(\ram[146][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n216));
   AO22CHD U4356 (.O(n2931), 
	.B2(n348), 
	.B1(\ram[146][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n216));
   AO22CHD U4357 (.O(n2932), 
	.B2(n348), 
	.B1(\ram[146][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n216));
   AO22CHD U4358 (.O(n2933), 
	.B2(n348), 
	.B1(\ram[146][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n216));
   AO22CHD U4359 (.O(n2934), 
	.B2(n350), 
	.B1(\ram[147][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n218));
   AO22CHD U4360 (.O(n2935), 
	.B2(n350), 
	.B1(\ram[147][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n218));
   AO22CHD U4361 (.O(n2936), 
	.B2(n350), 
	.B1(\ram[147][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n218));
   AO22CHD U4362 (.O(n2937), 
	.B2(n350), 
	.B1(\ram[147][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n218));
   AO22CHD U4363 (.O(n2938), 
	.B2(n350), 
	.B1(\ram[147][4] ), 
	.A2(n12), 
	.A1(n218));
   AO22CHD U4364 (.O(n2939), 
	.B2(n350), 
	.B1(\ram[147][5] ), 
	.A2(n13), 
	.A1(n218));
   AO22CHD U4365 (.O(n2940), 
	.B2(n350), 
	.B1(\ram[147][6] ), 
	.A2(n14), 
	.A1(n218));
   AO22CHD U4366 (.O(n2941), 
	.B2(n350), 
	.B1(\ram[147][7] ), 
	.A2(n15), 
	.A1(n218));
   AO22CHD U4367 (.O(n2942), 
	.B2(n350), 
	.B1(\ram[147][8] ), 
	.A2(n16), 
	.A1(n218));
   AO22CHD U4368 (.O(n2943), 
	.B2(n350), 
	.B1(\ram[147][9] ), 
	.A2(n17), 
	.A1(n218));
   AO22CHD U4369 (.O(n2944), 
	.B2(n350), 
	.B1(\ram[147][10] ), 
	.A2(n18), 
	.A1(n218));
   AO22CHD U4370 (.O(n2945), 
	.B2(n350), 
	.B1(\ram[147][11] ), 
	.A2(n19), 
	.A1(n218));
   AO22CHD U4371 (.O(n2946), 
	.B2(n350), 
	.B1(\ram[147][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n218));
   AO22CHD U4372 (.O(n2947), 
	.B2(n350), 
	.B1(\ram[147][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n218));
   AO22CHD U4373 (.O(n2948), 
	.B2(n350), 
	.B1(\ram[147][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n218));
   AO22CHD U4374 (.O(n2949), 
	.B2(n350), 
	.B1(\ram[147][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n218));
   AO22CHD U4375 (.O(n2950), 
	.B2(n352), 
	.B1(\ram[148][0] ), 
	.A2(n6), 
	.A1(n220));
   AO22CHD U4376 (.O(n2951), 
	.B2(n352), 
	.B1(\ram[148][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n220));
   AO22CHD U4377 (.O(n2952), 
	.B2(n352), 
	.B1(\ram[148][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n220));
   AO22CHD U4378 (.O(n2953), 
	.B2(n352), 
	.B1(\ram[148][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n220));
   AO22CHD U4379 (.O(n2954), 
	.B2(n352), 
	.B1(\ram[148][4] ), 
	.A2(n12), 
	.A1(n220));
   AO22CHD U4380 (.O(n2955), 
	.B2(n352), 
	.B1(\ram[148][5] ), 
	.A2(n13), 
	.A1(n220));
   AO22CHD U4381 (.O(n2956), 
	.B2(n352), 
	.B1(\ram[148][6] ), 
	.A2(n14), 
	.A1(n220));
   AO22CHD U4382 (.O(n2957), 
	.B2(n352), 
	.B1(\ram[148][7] ), 
	.A2(n15), 
	.A1(n220));
   AO22CHD U4383 (.O(n2958), 
	.B2(n352), 
	.B1(\ram[148][8] ), 
	.A2(n16), 
	.A1(n220));
   AO22CHD U4384 (.O(n2959), 
	.B2(n352), 
	.B1(\ram[148][9] ), 
	.A2(n17), 
	.A1(n220));
   AO22CHD U4385 (.O(n2960), 
	.B2(n352), 
	.B1(\ram[148][10] ), 
	.A2(n18), 
	.A1(n220));
   AO22CHD U4386 (.O(n2961), 
	.B2(n352), 
	.B1(\ram[148][11] ), 
	.A2(n19), 
	.A1(n220));
   AO22CHD U4387 (.O(n2962), 
	.B2(n352), 
	.B1(\ram[148][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n220));
   AO22CHD U4388 (.O(n2963), 
	.B2(n352), 
	.B1(\ram[148][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n220));
   AO22CHD U4389 (.O(n2964), 
	.B2(n352), 
	.B1(\ram[148][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n220));
   AO22CHD U4390 (.O(n2965), 
	.B2(n352), 
	.B1(\ram[148][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n220));
   AO22CHD U4391 (.O(n2966), 
	.B2(n354), 
	.B1(\ram[149][0] ), 
	.A2(n6), 
	.A1(n222));
   AO22CHD U4392 (.O(n2967), 
	.B2(n354), 
	.B1(\ram[149][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n222));
   AO22CHD U4393 (.O(n2968), 
	.B2(n354), 
	.B1(\ram[149][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n222));
   AO22CHD U4394 (.O(n2969), 
	.B2(n354), 
	.B1(\ram[149][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n222));
   AO22CHD U4395 (.O(n2970), 
	.B2(n354), 
	.B1(\ram[149][4] ), 
	.A2(n12), 
	.A1(n222));
   AO22CHD U4396 (.O(n2971), 
	.B2(n354), 
	.B1(\ram[149][5] ), 
	.A2(n13), 
	.A1(n222));
   AO22CHD U4397 (.O(n2972), 
	.B2(n354), 
	.B1(\ram[149][6] ), 
	.A2(n14), 
	.A1(n222));
   AO22CHD U4398 (.O(n2973), 
	.B2(n354), 
	.B1(\ram[149][7] ), 
	.A2(n15), 
	.A1(n222));
   AO22CHD U4399 (.O(n2974), 
	.B2(n354), 
	.B1(\ram[149][8] ), 
	.A2(n16), 
	.A1(n222));
   AO22CHD U4400 (.O(n2975), 
	.B2(n354), 
	.B1(\ram[149][9] ), 
	.A2(n17), 
	.A1(n222));
   AO22CHD U4401 (.O(n2976), 
	.B2(n354), 
	.B1(\ram[149][10] ), 
	.A2(n18), 
	.A1(n222));
   AO22CHD U4402 (.O(n2977), 
	.B2(n354), 
	.B1(\ram[149][11] ), 
	.A2(n19), 
	.A1(n222));
   AO22CHD U4403 (.O(n2978), 
	.B2(n354), 
	.B1(\ram[149][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n222));
   AO22CHD U4404 (.O(n2979), 
	.B2(n354), 
	.B1(\ram[149][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n222));
   AO22CHD U4405 (.O(n2980), 
	.B2(n354), 
	.B1(\ram[149][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n222));
   AO22CHD U4406 (.O(n2981), 
	.B2(n354), 
	.B1(\ram[149][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n222));
   AO22CHD U4407 (.O(n2982), 
	.B2(n356), 
	.B1(\ram[150][0] ), 
	.A2(n6), 
	.A1(n224));
   AO22CHD U4408 (.O(n2983), 
	.B2(n356), 
	.B1(\ram[150][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n224));
   AO22CHD U4409 (.O(n2984), 
	.B2(n356), 
	.B1(\ram[150][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n224));
   AO22CHD U4410 (.O(n2985), 
	.B2(n356), 
	.B1(\ram[150][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n224));
   AO22CHD U4411 (.O(n2986), 
	.B2(n356), 
	.B1(\ram[150][4] ), 
	.A2(n12), 
	.A1(n224));
   AO22CHD U4412 (.O(n2987), 
	.B2(n356), 
	.B1(\ram[150][5] ), 
	.A2(n13), 
	.A1(n224));
   AO22CHD U4413 (.O(n2988), 
	.B2(n356), 
	.B1(\ram[150][6] ), 
	.A2(n14), 
	.A1(n224));
   AO22CHD U4414 (.O(n2989), 
	.B2(n356), 
	.B1(\ram[150][7] ), 
	.A2(n15), 
	.A1(n224));
   AO22CHD U4415 (.O(n2990), 
	.B2(n356), 
	.B1(\ram[150][8] ), 
	.A2(n16), 
	.A1(n224));
   AO22CHD U4416 (.O(n2991), 
	.B2(n356), 
	.B1(\ram[150][9] ), 
	.A2(n17), 
	.A1(n224));
   AO22CHD U4417 (.O(n2992), 
	.B2(n356), 
	.B1(\ram[150][10] ), 
	.A2(n18), 
	.A1(n224));
   AO22CHD U4418 (.O(n2993), 
	.B2(n356), 
	.B1(\ram[150][11] ), 
	.A2(n19), 
	.A1(n224));
   AO22CHD U4419 (.O(n2994), 
	.B2(n356), 
	.B1(\ram[150][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n224));
   AO22CHD U4420 (.O(n2995), 
	.B2(n356), 
	.B1(\ram[150][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n224));
   AO22CHD U4421 (.O(n2996), 
	.B2(n356), 
	.B1(\ram[150][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n224));
   AO22CHD U4422 (.O(n2997), 
	.B2(n356), 
	.B1(\ram[150][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n224));
   AO22CHD U4423 (.O(n2998), 
	.B2(n358), 
	.B1(\ram[151][0] ), 
	.A2(n6), 
	.A1(n226));
   AO22CHD U4424 (.O(n2999), 
	.B2(n358), 
	.B1(\ram[151][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n226));
   AO22CHD U4425 (.O(n3000), 
	.B2(n358), 
	.B1(\ram[151][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n226));
   AO22CHD U4426 (.O(n3001), 
	.B2(n358), 
	.B1(\ram[151][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n226));
   AO22CHD U4427 (.O(n3002), 
	.B2(n358), 
	.B1(\ram[151][4] ), 
	.A2(n12), 
	.A1(n226));
   AO22CHD U4428 (.O(n3003), 
	.B2(n358), 
	.B1(\ram[151][5] ), 
	.A2(n13), 
	.A1(n226));
   AO22CHD U4429 (.O(n3004), 
	.B2(n358), 
	.B1(\ram[151][6] ), 
	.A2(n14), 
	.A1(n226));
   AO22CHD U4430 (.O(n3005), 
	.B2(n358), 
	.B1(\ram[151][7] ), 
	.A2(n15), 
	.A1(n226));
   AO22CHD U4431 (.O(n3006), 
	.B2(n358), 
	.B1(\ram[151][8] ), 
	.A2(n16), 
	.A1(n226));
   AO22CHD U4432 (.O(n3007), 
	.B2(n358), 
	.B1(\ram[151][9] ), 
	.A2(n17), 
	.A1(n226));
   AO22CHD U4433 (.O(n3008), 
	.B2(n358), 
	.B1(\ram[151][10] ), 
	.A2(n18), 
	.A1(n226));
   AO22CHD U4434 (.O(n3009), 
	.B2(n358), 
	.B1(\ram[151][11] ), 
	.A2(n19), 
	.A1(n226));
   AO22CHD U4435 (.O(n3010), 
	.B2(n358), 
	.B1(\ram[151][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n226));
   AO22CHD U4436 (.O(n3011), 
	.B2(n358), 
	.B1(\ram[151][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n226));
   AO22CHD U4437 (.O(n3012), 
	.B2(n358), 
	.B1(\ram[151][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n226));
   AO22CHD U4438 (.O(n3013), 
	.B2(n358), 
	.B1(\ram[151][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n226));
   AO22CHD U4439 (.O(n3014), 
	.B2(n360), 
	.B1(\ram[152][0] ), 
	.A2(n6), 
	.A1(n228));
   AO22CHD U4440 (.O(n3015), 
	.B2(n360), 
	.B1(\ram[152][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n228));
   AO22CHD U4441 (.O(n3016), 
	.B2(n360), 
	.B1(\ram[152][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n228));
   AO22CHD U4442 (.O(n3017), 
	.B2(n360), 
	.B1(\ram[152][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n228));
   AO22CHD U4443 (.O(n3018), 
	.B2(n360), 
	.B1(\ram[152][4] ), 
	.A2(n12), 
	.A1(n228));
   AO22CHD U4444 (.O(n3019), 
	.B2(n360), 
	.B1(\ram[152][5] ), 
	.A2(n13), 
	.A1(n228));
   AO22CHD U4445 (.O(n3020), 
	.B2(n360), 
	.B1(\ram[152][6] ), 
	.A2(n14), 
	.A1(n228));
   AO22CHD U4446 (.O(n3021), 
	.B2(n360), 
	.B1(\ram[152][7] ), 
	.A2(n15), 
	.A1(n228));
   AO22CHD U4447 (.O(n3022), 
	.B2(n360), 
	.B1(\ram[152][8] ), 
	.A2(n16), 
	.A1(n228));
   AO22CHD U4448 (.O(n3023), 
	.B2(n360), 
	.B1(\ram[152][9] ), 
	.A2(n17), 
	.A1(n228));
   AO22CHD U4449 (.O(n3024), 
	.B2(n360), 
	.B1(\ram[152][10] ), 
	.A2(n18), 
	.A1(n228));
   AO22CHD U4450 (.O(n3025), 
	.B2(n360), 
	.B1(\ram[152][11] ), 
	.A2(n19), 
	.A1(n228));
   AO22CHD U4451 (.O(n3026), 
	.B2(n360), 
	.B1(\ram[152][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n228));
   AO22CHD U4452 (.O(n3027), 
	.B2(n360), 
	.B1(\ram[152][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n228));
   AO22CHD U4453 (.O(n3028), 
	.B2(n360), 
	.B1(\ram[152][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n228));
   AO22CHD U4454 (.O(n3029), 
	.B2(n360), 
	.B1(\ram[152][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n228));
   AO22CHD U4455 (.O(n3030), 
	.B2(n362), 
	.B1(\ram[153][0] ), 
	.A2(n6), 
	.A1(n230));
   AO22CHD U4456 (.O(n3031), 
	.B2(n362), 
	.B1(\ram[153][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n230));
   AO22CHD U4457 (.O(n3032), 
	.B2(n362), 
	.B1(\ram[153][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n230));
   AO22CHD U4458 (.O(n3033), 
	.B2(n362), 
	.B1(\ram[153][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n230));
   AO22CHD U4459 (.O(n3034), 
	.B2(n362), 
	.B1(\ram[153][4] ), 
	.A2(n12), 
	.A1(n230));
   AO22CHD U4460 (.O(n3035), 
	.B2(n362), 
	.B1(\ram[153][5] ), 
	.A2(n13), 
	.A1(n230));
   AO22CHD U4461 (.O(n3036), 
	.B2(n362), 
	.B1(\ram[153][6] ), 
	.A2(n14), 
	.A1(n230));
   AO22CHD U4462 (.O(n3037), 
	.B2(n362), 
	.B1(FE_PHN4257_ram_153__7_), 
	.A2(n15), 
	.A1(n230));
   AO22CHD U4463 (.O(n3038), 
	.B2(n362), 
	.B1(\ram[153][8] ), 
	.A2(n16), 
	.A1(n230));
   AO22CHD U4464 (.O(n3039), 
	.B2(n362), 
	.B1(\ram[153][9] ), 
	.A2(n17), 
	.A1(n230));
   AO22CHD U4465 (.O(n3040), 
	.B2(n362), 
	.B1(\ram[153][10] ), 
	.A2(n18), 
	.A1(n230));
   AO22CHD U4466 (.O(n3041), 
	.B2(n362), 
	.B1(FE_PHN4406_ram_153__11_), 
	.A2(n19), 
	.A1(n230));
   AO22CHD U4467 (.O(n3042), 
	.B2(n362), 
	.B1(\ram[153][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n230));
   AO22CHD U4468 (.O(n3043), 
	.B2(n362), 
	.B1(\ram[153][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n230));
   AO22CHD U4469 (.O(n3044), 
	.B2(n362), 
	.B1(\ram[153][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n230));
   AO22CHD U4470 (.O(n3045), 
	.B2(n362), 
	.B1(\ram[153][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n230));
   AO22CHD U4471 (.O(n3046), 
	.B2(n364), 
	.B1(\ram[154][0] ), 
	.A2(n6), 
	.A1(n232));
   AO22CHD U4472 (.O(n3047), 
	.B2(n364), 
	.B1(\ram[154][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n232));
   AO22CHD U4473 (.O(n3048), 
	.B2(n364), 
	.B1(\ram[154][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n232));
   AO22CHD U4474 (.O(n3049), 
	.B2(n364), 
	.B1(\ram[154][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n232));
   AO22CHD U4475 (.O(n3050), 
	.B2(n364), 
	.B1(\ram[154][4] ), 
	.A2(n12), 
	.A1(n232));
   AO22CHD U4476 (.O(n3051), 
	.B2(n364), 
	.B1(FE_PHN4358_ram_154__5_), 
	.A2(n13), 
	.A1(n232));
   AO22CHD U4477 (.O(FE_PHN7307_n3052), 
	.B2(n364), 
	.B1(\ram[154][6] ), 
	.A2(n14), 
	.A1(n232));
   AO22CHD U4478 (.O(n3053), 
	.B2(n364), 
	.B1(\ram[154][7] ), 
	.A2(n15), 
	.A1(n232));
   AO22CHD U4479 (.O(n3054), 
	.B2(n364), 
	.B1(\ram[154][8] ), 
	.A2(n16), 
	.A1(n232));
   AO22CHD U4480 (.O(n3055), 
	.B2(n364), 
	.B1(\ram[154][9] ), 
	.A2(n17), 
	.A1(n232));
   AO22CHD U4481 (.O(n3056), 
	.B2(n364), 
	.B1(\ram[154][10] ), 
	.A2(n18), 
	.A1(n232));
   AO22CHD U4482 (.O(n3057), 
	.B2(n364), 
	.B1(\ram[154][11] ), 
	.A2(n19), 
	.A1(n232));
   AO22CHD U4483 (.O(n3058), 
	.B2(n364), 
	.B1(\ram[154][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n232));
   AO22CHD U4484 (.O(n3059), 
	.B2(n364), 
	.B1(\ram[154][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n232));
   AO22CHD U4485 (.O(n3060), 
	.B2(n364), 
	.B1(\ram[154][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n232));
   AO22CHD U4486 (.O(n3061), 
	.B2(n364), 
	.B1(\ram[154][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n232));
   AO22CHD U4487 (.O(n3062), 
	.B2(n366), 
	.B1(\ram[155][0] ), 
	.A2(n6), 
	.A1(n234));
   AO22CHD U4488 (.O(n3063), 
	.B2(n366), 
	.B1(\ram[155][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n234));
   AO22CHD U4489 (.O(n3064), 
	.B2(n366), 
	.B1(\ram[155][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n234));
   AO22CHD U4490 (.O(n3065), 
	.B2(n366), 
	.B1(\ram[155][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n234));
   AO22CHD U4491 (.O(n3066), 
	.B2(n366), 
	.B1(\ram[155][4] ), 
	.A2(n12), 
	.A1(n234));
   AO22CHD U4492 (.O(n3067), 
	.B2(n366), 
	.B1(\ram[155][5] ), 
	.A2(n13), 
	.A1(n234));
   AO22CHD U4493 (.O(n3068), 
	.B2(n366), 
	.B1(\ram[155][6] ), 
	.A2(n14), 
	.A1(n234));
   AO22CHD U4494 (.O(n3069), 
	.B2(n366), 
	.B1(\ram[155][7] ), 
	.A2(n15), 
	.A1(n234));
   AO22CHD U4495 (.O(n3070), 
	.B2(n366), 
	.B1(\ram[155][8] ), 
	.A2(n16), 
	.A1(n234));
   AO22CHD U4496 (.O(n3071), 
	.B2(n366), 
	.B1(\ram[155][9] ), 
	.A2(n17), 
	.A1(n234));
   AO22CHD U4497 (.O(n3072), 
	.B2(n366), 
	.B1(\ram[155][10] ), 
	.A2(n18), 
	.A1(n234));
   AO22CHD U4498 (.O(n3073), 
	.B2(n366), 
	.B1(\ram[155][11] ), 
	.A2(n19), 
	.A1(n234));
   AO22CHD U4499 (.O(n3074), 
	.B2(n366), 
	.B1(\ram[155][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n234));
   AO22CHD U4500 (.O(n3075), 
	.B2(n366), 
	.B1(\ram[155][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n234));
   AO22CHD U4501 (.O(n3076), 
	.B2(n366), 
	.B1(\ram[155][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n234));
   AO22CHD U4502 (.O(n3077), 
	.B2(n366), 
	.B1(\ram[155][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n234));
   AO22CHD U4503 (.O(n3078), 
	.B2(n368), 
	.B1(\ram[156][0] ), 
	.A2(n6), 
	.A1(n236));
   AO22CHD U4504 (.O(n3079), 
	.B2(n368), 
	.B1(\ram[156][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n236));
   AO22CHD U4505 (.O(n3080), 
	.B2(n368), 
	.B1(\ram[156][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n236));
   AO22CHD U4506 (.O(n3081), 
	.B2(n368), 
	.B1(\ram[156][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n236));
   AO22CHD U4507 (.O(n3082), 
	.B2(n368), 
	.B1(\ram[156][4] ), 
	.A2(n12), 
	.A1(n236));
   AO22CHD U4508 (.O(n3083), 
	.B2(n368), 
	.B1(\ram[156][5] ), 
	.A2(n13), 
	.A1(n236));
   AO22CHD U4509 (.O(n3084), 
	.B2(n368), 
	.B1(\ram[156][6] ), 
	.A2(n14), 
	.A1(n236));
   AO22CHD U4510 (.O(n3085), 
	.B2(n368), 
	.B1(\ram[156][7] ), 
	.A2(n15), 
	.A1(n236));
   AO22CHD U4511 (.O(n3086), 
	.B2(n368), 
	.B1(\ram[156][8] ), 
	.A2(n16), 
	.A1(n236));
   AO22CHD U4512 (.O(n3087), 
	.B2(n368), 
	.B1(\ram[156][9] ), 
	.A2(n17), 
	.A1(n236));
   AO22CHD U4513 (.O(n3088), 
	.B2(n368), 
	.B1(\ram[156][10] ), 
	.A2(n18), 
	.A1(n236));
   AO22CHD U4514 (.O(n3089), 
	.B2(n368), 
	.B1(\ram[156][11] ), 
	.A2(n19), 
	.A1(n236));
   AO22CHD U4515 (.O(n3090), 
	.B2(n368), 
	.B1(\ram[156][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n236));
   AO22CHD U4516 (.O(n3091), 
	.B2(n368), 
	.B1(\ram[156][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n236));
   AO22CHD U4517 (.O(n3092), 
	.B2(n368), 
	.B1(\ram[156][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n236));
   AO22CHD U4518 (.O(n3093), 
	.B2(n368), 
	.B1(\ram[156][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n236));
   AO22CHD U4519 (.O(n3094), 
	.B2(n370), 
	.B1(\ram[157][0] ), 
	.A2(n6), 
	.A1(n238));
   AO22CHD U4520 (.O(n3095), 
	.B2(n370), 
	.B1(\ram[157][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n238));
   AO22CHD U4521 (.O(n3096), 
	.B2(n370), 
	.B1(\ram[157][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n238));
   AO22CHD U4522 (.O(n3097), 
	.B2(n370), 
	.B1(\ram[157][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n238));
   AO22CHD U4523 (.O(n3098), 
	.B2(n370), 
	.B1(\ram[157][4] ), 
	.A2(n12), 
	.A1(n238));
   AO22CHD U4524 (.O(n3099), 
	.B2(n370), 
	.B1(\ram[157][5] ), 
	.A2(n13), 
	.A1(n238));
   AO22CHD U4525 (.O(n3100), 
	.B2(n370), 
	.B1(\ram[157][6] ), 
	.A2(n14), 
	.A1(n238));
   AO22CHD U4526 (.O(n3101), 
	.B2(n370), 
	.B1(\ram[157][7] ), 
	.A2(n15), 
	.A1(n238));
   AO22CHD U4527 (.O(n3102), 
	.B2(n370), 
	.B1(\ram[157][8] ), 
	.A2(n16), 
	.A1(n238));
   AO22CHD U4528 (.O(n3103), 
	.B2(n370), 
	.B1(\ram[157][9] ), 
	.A2(n17), 
	.A1(n238));
   AO22CHD U4529 (.O(n3104), 
	.B2(n370), 
	.B1(\ram[157][10] ), 
	.A2(n18), 
	.A1(n238));
   AO22CHD U4530 (.O(n3105), 
	.B2(n370), 
	.B1(\ram[157][11] ), 
	.A2(n19), 
	.A1(n238));
   AO22CHD U4531 (.O(n3106), 
	.B2(n370), 
	.B1(\ram[157][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n238));
   AO22CHD U4532 (.O(n3107), 
	.B2(n370), 
	.B1(\ram[157][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n238));
   AO22CHD U4533 (.O(n3108), 
	.B2(n370), 
	.B1(\ram[157][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n238));
   AO22CHD U4534 (.O(n3109), 
	.B2(n370), 
	.B1(\ram[157][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n238));
   AO22CHD U4535 (.O(n3110), 
	.B2(n372), 
	.B1(\ram[158][0] ), 
	.A2(n6), 
	.A1(n240));
   AO22CHD U4536 (.O(n3111), 
	.B2(n372), 
	.B1(\ram[158][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n240));
   AO22CHD U4537 (.O(n3112), 
	.B2(n372), 
	.B1(\ram[158][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n240));
   AO22CHD U4538 (.O(n3113), 
	.B2(n372), 
	.B1(\ram[158][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n240));
   AO22CHD U4539 (.O(n3114), 
	.B2(n372), 
	.B1(\ram[158][4] ), 
	.A2(n12), 
	.A1(n240));
   AO22CHD U4540 (.O(n3115), 
	.B2(n372), 
	.B1(\ram[158][5] ), 
	.A2(n13), 
	.A1(n240));
   AO22CHD U4541 (.O(n3116), 
	.B2(n372), 
	.B1(\ram[158][6] ), 
	.A2(n14), 
	.A1(n240));
   AO22CHD U4542 (.O(n3117), 
	.B2(n372), 
	.B1(\ram[158][7] ), 
	.A2(n15), 
	.A1(n240));
   AO22CHD U4543 (.O(n3118), 
	.B2(n372), 
	.B1(\ram[158][8] ), 
	.A2(n16), 
	.A1(n240));
   AO22CHD U4544 (.O(n3119), 
	.B2(n372), 
	.B1(\ram[158][9] ), 
	.A2(n17), 
	.A1(n240));
   AO22CHD U4545 (.O(n3120), 
	.B2(n372), 
	.B1(\ram[158][10] ), 
	.A2(n18), 
	.A1(n240));
   AO22CHD U4546 (.O(n3121), 
	.B2(n372), 
	.B1(FE_PHN4527_ram_158__11_), 
	.A2(n19), 
	.A1(n240));
   AO22CHD U4547 (.O(n3122), 
	.B2(n372), 
	.B1(\ram[158][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n240));
   AO22CHD U4548 (.O(n3123), 
	.B2(n372), 
	.B1(\ram[158][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n240));
   AO22CHD U4549 (.O(n3124), 
	.B2(n372), 
	.B1(\ram[158][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n240));
   AO22CHD U4550 (.O(n3125), 
	.B2(n372), 
	.B1(\ram[158][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n240));
   AO22CHD U4551 (.O(n3126), 
	.B2(n374), 
	.B1(\ram[159][0] ), 
	.A2(n6), 
	.A1(n242));
   AO22CHD U4552 (.O(n3127), 
	.B2(n374), 
	.B1(\ram[159][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n242));
   AO22CHD U4553 (.O(n3128), 
	.B2(n374), 
	.B1(\ram[159][2] ), 
	.A2(FE_OFN47_n10), 
	.A1(n242));
   AO22CHD U4554 (.O(FE_PHN7293_n3129), 
	.B2(n374), 
	.B1(\ram[159][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n242));
   AO22CHD U4555 (.O(n3130), 
	.B2(n374), 
	.B1(\ram[159][4] ), 
	.A2(n12), 
	.A1(n242));
   AO22CHD U4556 (.O(n3131), 
	.B2(n374), 
	.B1(\ram[159][5] ), 
	.A2(n13), 
	.A1(n242));
   AO22CHD U4557 (.O(n3132), 
	.B2(n374), 
	.B1(\ram[159][6] ), 
	.A2(n14), 
	.A1(n242));
   AO22CHD U4558 (.O(n3133), 
	.B2(n374), 
	.B1(\ram[159][7] ), 
	.A2(n15), 
	.A1(n242));
   AO22CHD U4559 (.O(n3134), 
	.B2(n374), 
	.B1(\ram[159][8] ), 
	.A2(n16), 
	.A1(n242));
   AO22CHD U4560 (.O(n3135), 
	.B2(n374), 
	.B1(\ram[159][9] ), 
	.A2(n17), 
	.A1(n242));
   AO22CHD U4561 (.O(n3136), 
	.B2(n374), 
	.B1(\ram[159][10] ), 
	.A2(n18), 
	.A1(n242));
   AO22CHD U4562 (.O(n3137), 
	.B2(n374), 
	.B1(\ram[159][11] ), 
	.A2(n19), 
	.A1(n242));
   AO22CHD U4563 (.O(n3138), 
	.B2(n374), 
	.B1(\ram[159][12] ), 
	.A2(FE_OFN79_n20), 
	.A1(n242));
   AO22CHD U4564 (.O(n3139), 
	.B2(n374), 
	.B1(\ram[159][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n242));
   AO22CHD U4565 (.O(n3140), 
	.B2(n374), 
	.B1(\ram[159][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n242));
   AO22CHD U4566 (.O(n3141), 
	.B2(n374), 
	.B1(\ram[159][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n242));
   AO22CHD U4567 (.O(n3142), 
	.B2(n376), 
	.B1(\ram[160][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n244));
   AO22CHD U4568 (.O(n3143), 
	.B2(n376), 
	.B1(\ram[160][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n244));
   AO22CHD U4569 (.O(n3144), 
	.B2(n376), 
	.B1(\ram[160][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n244));
   AO22CHD U4570 (.O(n3145), 
	.B2(n376), 
	.B1(\ram[160][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n244));
   AO22CHD U4571 (.O(n3146), 
	.B2(n376), 
	.B1(\ram[160][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n244));
   AO22CHD U4572 (.O(n3147), 
	.B2(n376), 
	.B1(\ram[160][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n244));
   AO22CHD U4573 (.O(n3148), 
	.B2(n376), 
	.B1(\ram[160][6] ), 
	.A2(n14), 
	.A1(n244));
   AO22CHD U4574 (.O(n3149), 
	.B2(n376), 
	.B1(\ram[160][7] ), 
	.A2(n15), 
	.A1(n244));
   AO22CHD U4575 (.O(n3150), 
	.B2(n376), 
	.B1(\ram[160][8] ), 
	.A2(n16), 
	.A1(n244));
   AO22CHD U4576 (.O(n3151), 
	.B2(n376), 
	.B1(\ram[160][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n244));
   AO22CHD U4577 (.O(n3152), 
	.B2(n376), 
	.B1(\ram[160][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n244));
   AO22CHD U4578 (.O(n3153), 
	.B2(n376), 
	.B1(\ram[160][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n244));
   AO22CHD U4579 (.O(n3154), 
	.B2(n376), 
	.B1(\ram[160][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n244));
   AO22CHD U4580 (.O(n3155), 
	.B2(n376), 
	.B1(\ram[160][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n244));
   AO22CHD U4581 (.O(n3156), 
	.B2(n376), 
	.B1(\ram[160][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n244));
   AO22CHD U4582 (.O(n3157), 
	.B2(n376), 
	.B1(\ram[160][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n244));
   AO22CHD U4583 (.O(n3158), 
	.B2(n379), 
	.B1(\ram[161][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n245));
   AO22CHD U4584 (.O(n3159), 
	.B2(n379), 
	.B1(\ram[161][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n245));
   AO22CHD U4585 (.O(n3160), 
	.B2(n379), 
	.B1(\ram[161][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n245));
   AO22CHD U4586 (.O(n3161), 
	.B2(n379), 
	.B1(\ram[161][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n245));
   AO22CHD U4587 (.O(n3162), 
	.B2(n379), 
	.B1(\ram[161][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n245));
   AO22CHD U4588 (.O(n3163), 
	.B2(n379), 
	.B1(\ram[161][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n245));
   AO22CHD U4589 (.O(n3164), 
	.B2(n379), 
	.B1(\ram[161][6] ), 
	.A2(n14), 
	.A1(n245));
   AO22CHD U4590 (.O(n3165), 
	.B2(n379), 
	.B1(\ram[161][7] ), 
	.A2(n15), 
	.A1(n245));
   AO22CHD U4591 (.O(n3166), 
	.B2(n379), 
	.B1(\ram[161][8] ), 
	.A2(n16), 
	.A1(n245));
   AO22CHD U4592 (.O(n3167), 
	.B2(n379), 
	.B1(\ram[161][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n245));
   AO22CHD U4593 (.O(n3168), 
	.B2(n379), 
	.B1(\ram[161][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n245));
   AO22CHD U4594 (.O(n3169), 
	.B2(n379), 
	.B1(\ram[161][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n245));
   AO22CHD U4595 (.O(n3170), 
	.B2(n379), 
	.B1(\ram[161][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n245));
   AO22CHD U4596 (.O(n3171), 
	.B2(n379), 
	.B1(\ram[161][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n245));
   AO22CHD U4597 (.O(n3172), 
	.B2(n379), 
	.B1(\ram[161][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n245));
   AO22CHD U4598 (.O(n3173), 
	.B2(n379), 
	.B1(\ram[161][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n245));
   AO22CHD U4599 (.O(n3174), 
	.B2(n381), 
	.B1(\ram[162][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n247));
   AO22CHD U4600 (.O(n3175), 
	.B2(n381), 
	.B1(\ram[162][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n247));
   AO22CHD U4601 (.O(n3176), 
	.B2(n381), 
	.B1(\ram[162][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n247));
   AO22CHD U4602 (.O(n3177), 
	.B2(n381), 
	.B1(\ram[162][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n247));
   AO22CHD U4603 (.O(n3178), 
	.B2(n381), 
	.B1(\ram[162][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n247));
   AO22CHD U4604 (.O(n3179), 
	.B2(n381), 
	.B1(\ram[162][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n247));
   AO22CHD U4605 (.O(n3180), 
	.B2(n381), 
	.B1(\ram[162][6] ), 
	.A2(n14), 
	.A1(n247));
   AO22CHD U4606 (.O(n3181), 
	.B2(n381), 
	.B1(\ram[162][7] ), 
	.A2(n15), 
	.A1(n247));
   AO22CHD U4607 (.O(n3182), 
	.B2(n381), 
	.B1(\ram[162][8] ), 
	.A2(n16), 
	.A1(n247));
   AO22CHD U4608 (.O(n3183), 
	.B2(n381), 
	.B1(\ram[162][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n247));
   AO22CHD U4609 (.O(n3184), 
	.B2(n381), 
	.B1(\ram[162][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n247));
   AO22CHD U4610 (.O(n3185), 
	.B2(n381), 
	.B1(\ram[162][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n247));
   AO22CHD U4611 (.O(n3186), 
	.B2(n381), 
	.B1(\ram[162][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n247));
   AO22CHD U4612 (.O(n3187), 
	.B2(n381), 
	.B1(\ram[162][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n247));
   AO22CHD U4613 (.O(n3188), 
	.B2(n381), 
	.B1(\ram[162][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n247));
   AO22CHD U4614 (.O(n3189), 
	.B2(n381), 
	.B1(\ram[162][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n247));
   AO22CHD U4615 (.O(n3190), 
	.B2(n383), 
	.B1(\ram[163][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n249));
   AO22CHD U4616 (.O(n3191), 
	.B2(n383), 
	.B1(\ram[163][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n249));
   AO22CHD U4617 (.O(n3192), 
	.B2(n383), 
	.B1(\ram[163][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n249));
   AO22CHD U4618 (.O(n3193), 
	.B2(n383), 
	.B1(\ram[163][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n249));
   AO22CHD U4619 (.O(n3194), 
	.B2(n383), 
	.B1(\ram[163][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n249));
   AO22CHD U4620 (.O(n3195), 
	.B2(n383), 
	.B1(\ram[163][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n249));
   AO22CHD U4621 (.O(n3196), 
	.B2(n383), 
	.B1(\ram[163][6] ), 
	.A2(n14), 
	.A1(n249));
   AO22CHD U4622 (.O(n3197), 
	.B2(n383), 
	.B1(\ram[163][7] ), 
	.A2(n15), 
	.A1(n249));
   AO22CHD U4623 (.O(n3198), 
	.B2(n383), 
	.B1(\ram[163][8] ), 
	.A2(n16), 
	.A1(n249));
   AO22CHD U4624 (.O(n3199), 
	.B2(n383), 
	.B1(\ram[163][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n249));
   AO22CHD U4625 (.O(n3200), 
	.B2(n383), 
	.B1(\ram[163][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n249));
   AO22CHD U4626 (.O(n3201), 
	.B2(n383), 
	.B1(\ram[163][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n249));
   AO22CHD U4627 (.O(n3202), 
	.B2(n383), 
	.B1(\ram[163][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n249));
   AO22CHD U4628 (.O(n3203), 
	.B2(n383), 
	.B1(\ram[163][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n249));
   AO22CHD U4629 (.O(n3204), 
	.B2(n383), 
	.B1(\ram[163][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n249));
   AO22CHD U4630 (.O(n3205), 
	.B2(n383), 
	.B1(\ram[163][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n249));
   AO22CHD U4631 (.O(n3206), 
	.B2(n385), 
	.B1(\ram[164][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n251));
   AO22CHD U4632 (.O(n3207), 
	.B2(n385), 
	.B1(\ram[164][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n251));
   AO22CHD U4633 (.O(n3208), 
	.B2(n385), 
	.B1(\ram[164][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n251));
   AO22CHD U4634 (.O(n3209), 
	.B2(n385), 
	.B1(\ram[164][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n251));
   AO22CHD U4635 (.O(n3210), 
	.B2(n385), 
	.B1(\ram[164][4] ), 
	.A2(n12), 
	.A1(n251));
   AO22CHD U4636 (.O(n3211), 
	.B2(n385), 
	.B1(\ram[164][5] ), 
	.A2(n13), 
	.A1(n251));
   AO22CHD U4637 (.O(n3212), 
	.B2(n385), 
	.B1(\ram[164][6] ), 
	.A2(n14), 
	.A1(n251));
   AO22CHD U4638 (.O(n3213), 
	.B2(n385), 
	.B1(\ram[164][7] ), 
	.A2(n15), 
	.A1(n251));
   AO22CHD U4639 (.O(n3214), 
	.B2(n385), 
	.B1(\ram[164][8] ), 
	.A2(n16), 
	.A1(n251));
   AO22CHD U4640 (.O(n3215), 
	.B2(n385), 
	.B1(\ram[164][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n251));
   AO22CHD U4641 (.O(n3216), 
	.B2(n385), 
	.B1(\ram[164][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n251));
   AO22CHD U4642 (.O(n3217), 
	.B2(n385), 
	.B1(\ram[164][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n251));
   AO22CHD U4643 (.O(n3218), 
	.B2(n385), 
	.B1(\ram[164][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n251));
   AO22CHD U4644 (.O(n3219), 
	.B2(n385), 
	.B1(\ram[164][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n251));
   AO22CHD U4645 (.O(n3220), 
	.B2(n385), 
	.B1(\ram[164][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n251));
   AO22CHD U4646 (.O(n3221), 
	.B2(n385), 
	.B1(\ram[164][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n251));
   AO22CHD U4647 (.O(n3222), 
	.B2(n387), 
	.B1(\ram[165][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n253));
   AO22CHD U4648 (.O(n3223), 
	.B2(n387), 
	.B1(\ram[165][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n253));
   AO22CHD U4649 (.O(n3224), 
	.B2(n387), 
	.B1(\ram[165][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n253));
   AO22CHD U4650 (.O(n3225), 
	.B2(n387), 
	.B1(\ram[165][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n253));
   AO22CHD U4651 (.O(n3226), 
	.B2(n387), 
	.B1(\ram[165][4] ), 
	.A2(n12), 
	.A1(n253));
   AO22CHD U4652 (.O(n3227), 
	.B2(n387), 
	.B1(\ram[165][5] ), 
	.A2(n13), 
	.A1(n253));
   AO22CHD U4653 (.O(n3228), 
	.B2(n387), 
	.B1(\ram[165][6] ), 
	.A2(n14), 
	.A1(n253));
   AO22CHD U4654 (.O(n3229), 
	.B2(n387), 
	.B1(\ram[165][7] ), 
	.A2(n15), 
	.A1(n253));
   AO22CHD U4655 (.O(n3230), 
	.B2(n387), 
	.B1(\ram[165][8] ), 
	.A2(n16), 
	.A1(n253));
   AO22CHD U4656 (.O(n3231), 
	.B2(n387), 
	.B1(\ram[165][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n253));
   AO22CHD U4657 (.O(n3232), 
	.B2(n387), 
	.B1(\ram[165][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n253));
   AO22CHD U4658 (.O(n3233), 
	.B2(n387), 
	.B1(\ram[165][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n253));
   AO22CHD U4659 (.O(n3234), 
	.B2(n387), 
	.B1(\ram[165][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n253));
   AO22CHD U4660 (.O(n3235), 
	.B2(n387), 
	.B1(\ram[165][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n253));
   AO22CHD U4661 (.O(n3236), 
	.B2(n387), 
	.B1(\ram[165][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n253));
   AO22CHD U4662 (.O(n3237), 
	.B2(n387), 
	.B1(\ram[165][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n253));
   AO22CHD U4663 (.O(n3238), 
	.B2(n389), 
	.B1(\ram[166][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n255));
   AO22CHD U4664 (.O(n3239), 
	.B2(n389), 
	.B1(\ram[166][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n255));
   AO22CHD U4665 (.O(n3240), 
	.B2(n389), 
	.B1(\ram[166][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n255));
   AO22CHD U4666 (.O(n3241), 
	.B2(n389), 
	.B1(\ram[166][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n255));
   AO22CHD U4667 (.O(n3242), 
	.B2(n389), 
	.B1(\ram[166][4] ), 
	.A2(n12), 
	.A1(n255));
   AO22CHD U4668 (.O(n3243), 
	.B2(n389), 
	.B1(\ram[166][5] ), 
	.A2(n13), 
	.A1(n255));
   AO22CHD U4669 (.O(n3244), 
	.B2(n389), 
	.B1(\ram[166][6] ), 
	.A2(n14), 
	.A1(n255));
   AO22CHD U4670 (.O(n3245), 
	.B2(n389), 
	.B1(\ram[166][7] ), 
	.A2(n15), 
	.A1(n255));
   AO22CHD U4671 (.O(n3246), 
	.B2(n389), 
	.B1(\ram[166][8] ), 
	.A2(n16), 
	.A1(n255));
   AO22CHD U4672 (.O(n3247), 
	.B2(n389), 
	.B1(\ram[166][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n255));
   AO22CHD U4673 (.O(n3248), 
	.B2(n389), 
	.B1(\ram[166][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n255));
   AO22CHD U4674 (.O(n3249), 
	.B2(n389), 
	.B1(\ram[166][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n255));
   AO22CHD U4675 (.O(n3250), 
	.B2(n389), 
	.B1(\ram[166][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n255));
   AO22CHD U4676 (.O(n3251), 
	.B2(n389), 
	.B1(\ram[166][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n255));
   AO22CHD U4677 (.O(n3252), 
	.B2(n389), 
	.B1(\ram[166][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n255));
   AO22CHD U4678 (.O(n3253), 
	.B2(n389), 
	.B1(\ram[166][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n255));
   AO22CHD U4679 (.O(n3254), 
	.B2(n391), 
	.B1(\ram[167][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n257));
   AO22CHD U4680 (.O(n3255), 
	.B2(n391), 
	.B1(\ram[167][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n257));
   AO22CHD U4681 (.O(n3256), 
	.B2(n391), 
	.B1(\ram[167][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n257));
   AO22CHD U4682 (.O(n3257), 
	.B2(n391), 
	.B1(\ram[167][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n257));
   AO22CHD U4683 (.O(n3258), 
	.B2(n391), 
	.B1(\ram[167][4] ), 
	.A2(n12), 
	.A1(n257));
   AO22CHD U4684 (.O(n3259), 
	.B2(n391), 
	.B1(\ram[167][5] ), 
	.A2(n13), 
	.A1(n257));
   AO22CHD U4685 (.O(n3260), 
	.B2(n391), 
	.B1(\ram[167][6] ), 
	.A2(n14), 
	.A1(n257));
   AO22CHD U4686 (.O(n3261), 
	.B2(n391), 
	.B1(\ram[167][7] ), 
	.A2(n15), 
	.A1(n257));
   AO22CHD U4687 (.O(n3262), 
	.B2(n391), 
	.B1(\ram[167][8] ), 
	.A2(n16), 
	.A1(n257));
   AO22CHD U4688 (.O(n3263), 
	.B2(n391), 
	.B1(\ram[167][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n257));
   AO22CHD U4689 (.O(n3264), 
	.B2(n391), 
	.B1(\ram[167][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n257));
   AO22CHD U4690 (.O(n3265), 
	.B2(n391), 
	.B1(\ram[167][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n257));
   AO22CHD U4691 (.O(n3266), 
	.B2(n391), 
	.B1(\ram[167][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n257));
   AO22CHD U4692 (.O(n3267), 
	.B2(n391), 
	.B1(\ram[167][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n257));
   AO22CHD U4693 (.O(n3268), 
	.B2(n391), 
	.B1(\ram[167][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n257));
   AO22CHD U4694 (.O(n3269), 
	.B2(n391), 
	.B1(\ram[167][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n257));
   AO22CHD U4695 (.O(n3270), 
	.B2(n393), 
	.B1(\ram[168][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n259));
   AO22CHD U4696 (.O(n3271), 
	.B2(n393), 
	.B1(\ram[168][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n259));
   AO22CHD U4697 (.O(n3272), 
	.B2(n393), 
	.B1(\ram[168][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n259));
   AO22CHD U4698 (.O(n3273), 
	.B2(n393), 
	.B1(\ram[168][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n259));
   AO22CHD U4699 (.O(n3274), 
	.B2(n393), 
	.B1(\ram[168][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n259));
   AO22CHD U4700 (.O(n3275), 
	.B2(n393), 
	.B1(\ram[168][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n259));
   AO22CHD U4701 (.O(n3276), 
	.B2(n393), 
	.B1(\ram[168][6] ), 
	.A2(n14), 
	.A1(n259));
   AO22CHD U4702 (.O(n3277), 
	.B2(n393), 
	.B1(\ram[168][7] ), 
	.A2(n15), 
	.A1(n259));
   AO22CHD U4703 (.O(n3278), 
	.B2(n393), 
	.B1(\ram[168][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n259));
   AO22CHD U4704 (.O(n3279), 
	.B2(n393), 
	.B1(\ram[168][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n259));
   AO22CHD U4705 (.O(n3280), 
	.B2(n393), 
	.B1(\ram[168][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n259));
   AO22CHD U4706 (.O(n3281), 
	.B2(n393), 
	.B1(\ram[168][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n259));
   AO22CHD U4707 (.O(n3282), 
	.B2(n393), 
	.B1(\ram[168][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n259));
   AO22CHD U4708 (.O(n3283), 
	.B2(n393), 
	.B1(\ram[168][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n259));
   AO22CHD U4709 (.O(n3284), 
	.B2(n393), 
	.B1(\ram[168][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n259));
   AO22CHD U4710 (.O(n3285), 
	.B2(n393), 
	.B1(\ram[168][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n259));
   AO22CHD U4711 (.O(n3286), 
	.B2(n395), 
	.B1(\ram[169][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n261));
   AO22CHD U4712 (.O(n3287), 
	.B2(n395), 
	.B1(\ram[169][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n261));
   AO22CHD U4713 (.O(n3288), 
	.B2(n395), 
	.B1(\ram[169][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n261));
   AO22CHD U4714 (.O(n3289), 
	.B2(n395), 
	.B1(\ram[169][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n261));
   AO22CHD U4715 (.O(n3290), 
	.B2(n395), 
	.B1(\ram[169][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n261));
   AO22CHD U4716 (.O(n3291), 
	.B2(n395), 
	.B1(\ram[169][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n261));
   AO22CHD U4717 (.O(n3292), 
	.B2(n395), 
	.B1(\ram[169][6] ), 
	.A2(n14), 
	.A1(n261));
   AO22CHD U4718 (.O(n3293), 
	.B2(n395), 
	.B1(\ram[169][7] ), 
	.A2(n15), 
	.A1(n261));
   AO22CHD U4719 (.O(n3294), 
	.B2(n395), 
	.B1(\ram[169][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n261));
   AO22CHD U4720 (.O(n3295), 
	.B2(n395), 
	.B1(\ram[169][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n261));
   AO22CHD U4721 (.O(n3296), 
	.B2(n395), 
	.B1(\ram[169][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n261));
   AO22CHD U4722 (.O(n3297), 
	.B2(n395), 
	.B1(\ram[169][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n261));
   AO22CHD U4723 (.O(n3298), 
	.B2(n395), 
	.B1(\ram[169][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n261));
   AO22CHD U4724 (.O(n3299), 
	.B2(n395), 
	.B1(\ram[169][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n261));
   AO22CHD U4725 (.O(n3300), 
	.B2(n395), 
	.B1(\ram[169][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n261));
   AO22CHD U4726 (.O(n3301), 
	.B2(n395), 
	.B1(\ram[169][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n261));
   AO22CHD U4727 (.O(n3302), 
	.B2(n397), 
	.B1(\ram[170][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n263));
   AO22CHD U4728 (.O(n3303), 
	.B2(n397), 
	.B1(\ram[170][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n263));
   AO22CHD U4729 (.O(n3304), 
	.B2(n397), 
	.B1(\ram[170][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n263));
   AO22CHD U4730 (.O(n3305), 
	.B2(n397), 
	.B1(\ram[170][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n263));
   AO22CHD U4731 (.O(n3306), 
	.B2(n397), 
	.B1(\ram[170][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n263));
   AO22CHD U4732 (.O(n3307), 
	.B2(n397), 
	.B1(\ram[170][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n263));
   AO22CHD U4733 (.O(n3308), 
	.B2(n397), 
	.B1(\ram[170][6] ), 
	.A2(n14), 
	.A1(n263));
   AO22CHD U4734 (.O(n3309), 
	.B2(n397), 
	.B1(\ram[170][7] ), 
	.A2(n15), 
	.A1(n263));
   AO22CHD U4735 (.O(n3310), 
	.B2(n397), 
	.B1(\ram[170][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n263));
   AO22CHD U4736 (.O(n3311), 
	.B2(n397), 
	.B1(\ram[170][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n263));
   AO22CHD U4737 (.O(n3312), 
	.B2(n397), 
	.B1(\ram[170][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n263));
   AO22CHD U4738 (.O(n3313), 
	.B2(n397), 
	.B1(\ram[170][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n263));
   AO22CHD U4739 (.O(n3314), 
	.B2(n397), 
	.B1(\ram[170][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n263));
   AO22CHD U4740 (.O(n3315), 
	.B2(n397), 
	.B1(\ram[170][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n263));
   AO22CHD U4741 (.O(n3316), 
	.B2(n397), 
	.B1(\ram[170][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n263));
   AO22CHD U4742 (.O(n3317), 
	.B2(n397), 
	.B1(\ram[170][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n263));
   AO22CHD U4743 (.O(n3318), 
	.B2(n399), 
	.B1(\ram[171][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n265));
   AO22CHD U4744 (.O(n3319), 
	.B2(n399), 
	.B1(\ram[171][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n265));
   AO22CHD U4745 (.O(n3320), 
	.B2(n399), 
	.B1(\ram[171][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n265));
   AO22CHD U4746 (.O(n3321), 
	.B2(n399), 
	.B1(\ram[171][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n265));
   AO22CHD U4747 (.O(n3322), 
	.B2(n399), 
	.B1(\ram[171][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n265));
   AO22CHD U4748 (.O(n3323), 
	.B2(n399), 
	.B1(\ram[171][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n265));
   AO22CHD U4749 (.O(n3324), 
	.B2(n399), 
	.B1(\ram[171][6] ), 
	.A2(n14), 
	.A1(n265));
   AO22CHD U4750 (.O(n3325), 
	.B2(n399), 
	.B1(\ram[171][7] ), 
	.A2(n15), 
	.A1(n265));
   AO22CHD U4751 (.O(n3326), 
	.B2(n399), 
	.B1(\ram[171][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n265));
   AO22CHD U4752 (.O(n3327), 
	.B2(n399), 
	.B1(\ram[171][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n265));
   AO22CHD U4753 (.O(n3328), 
	.B2(n399), 
	.B1(\ram[171][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n265));
   AO22CHD U4754 (.O(n3329), 
	.B2(n399), 
	.B1(\ram[171][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n265));
   AO22CHD U4755 (.O(n3330), 
	.B2(n399), 
	.B1(\ram[171][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n265));
   AO22CHD U4756 (.O(n3331), 
	.B2(n399), 
	.B1(\ram[171][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n265));
   AO22CHD U4757 (.O(n3332), 
	.B2(n399), 
	.B1(\ram[171][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n265));
   AO22CHD U4758 (.O(n3333), 
	.B2(n399), 
	.B1(\ram[171][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n265));
   AO22CHD U4759 (.O(n3334), 
	.B2(n401), 
	.B1(\ram[172][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n267));
   AO22CHD U4760 (.O(n3335), 
	.B2(n401), 
	.B1(\ram[172][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n267));
   AO22CHD U4761 (.O(n3336), 
	.B2(n401), 
	.B1(\ram[172][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n267));
   AO22CHD U4762 (.O(n3337), 
	.B2(n401), 
	.B1(\ram[172][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n267));
   AO22CHD U4763 (.O(n3338), 
	.B2(n401), 
	.B1(\ram[172][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n267));
   AO22CHD U4764 (.O(n3339), 
	.B2(n401), 
	.B1(\ram[172][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n267));
   AO22CHD U4765 (.O(n3340), 
	.B2(n401), 
	.B1(\ram[172][6] ), 
	.A2(n14), 
	.A1(n267));
   AO22CHD U4766 (.O(n3341), 
	.B2(n401), 
	.B1(\ram[172][7] ), 
	.A2(n15), 
	.A1(n267));
   AO22CHD U4767 (.O(n3342), 
	.B2(n401), 
	.B1(\ram[172][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n267));
   AO22CHD U4768 (.O(n3343), 
	.B2(n401), 
	.B1(\ram[172][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n267));
   AO22CHD U4769 (.O(n3344), 
	.B2(n401), 
	.B1(\ram[172][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n267));
   AO22CHD U4770 (.O(n3345), 
	.B2(n401), 
	.B1(\ram[172][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n267));
   AO22CHD U4771 (.O(n3346), 
	.B2(n401), 
	.B1(\ram[172][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n267));
   AO22CHD U4772 (.O(n3347), 
	.B2(n401), 
	.B1(\ram[172][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n267));
   AO22CHD U4773 (.O(n3348), 
	.B2(n401), 
	.B1(\ram[172][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n267));
   AO22CHD U4774 (.O(n3349), 
	.B2(n401), 
	.B1(\ram[172][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n267));
   AO22CHD U4775 (.O(n3350), 
	.B2(n403), 
	.B1(\ram[173][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n269));
   AO22CHD U4776 (.O(n3351), 
	.B2(n403), 
	.B1(\ram[173][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n269));
   AO22CHD U4777 (.O(n3352), 
	.B2(n403), 
	.B1(\ram[173][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n269));
   AO22CHD U4778 (.O(n3353), 
	.B2(n403), 
	.B1(\ram[173][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n269));
   AO22CHD U4779 (.O(n3354), 
	.B2(n403), 
	.B1(\ram[173][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n269));
   AO22CHD U4780 (.O(n3355), 
	.B2(n403), 
	.B1(\ram[173][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n269));
   AO22CHD U4781 (.O(n3356), 
	.B2(n403), 
	.B1(\ram[173][6] ), 
	.A2(n14), 
	.A1(n269));
   AO22CHD U4782 (.O(n3357), 
	.B2(n403), 
	.B1(\ram[173][7] ), 
	.A2(n15), 
	.A1(n269));
   AO22CHD U4783 (.O(n3358), 
	.B2(n403), 
	.B1(\ram[173][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n269));
   AO22CHD U4784 (.O(n3359), 
	.B2(n403), 
	.B1(\ram[173][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n269));
   AO22CHD U4785 (.O(n3360), 
	.B2(n403), 
	.B1(\ram[173][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n269));
   AO22CHD U4786 (.O(n3361), 
	.B2(n403), 
	.B1(\ram[173][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n269));
   AO22CHD U4787 (.O(n3362), 
	.B2(n403), 
	.B1(\ram[173][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n269));
   AO22CHD U4788 (.O(n3363), 
	.B2(n403), 
	.B1(\ram[173][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n269));
   AO22CHD U4789 (.O(n3364), 
	.B2(n403), 
	.B1(\ram[173][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n269));
   AO22CHD U4790 (.O(n3365), 
	.B2(n403), 
	.B1(\ram[173][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n269));
   AO22CHD U4791 (.O(n3366), 
	.B2(n405), 
	.B1(\ram[174][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n271));
   AO22CHD U4792 (.O(n3367), 
	.B2(n405), 
	.B1(\ram[174][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n271));
   AO22CHD U4793 (.O(n3368), 
	.B2(n405), 
	.B1(\ram[174][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n271));
   AO22CHD U4794 (.O(n3369), 
	.B2(n405), 
	.B1(\ram[174][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n271));
   AO22CHD U4795 (.O(n3370), 
	.B2(n405), 
	.B1(\ram[174][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n271));
   AO22CHD U4796 (.O(n3371), 
	.B2(n405), 
	.B1(\ram[174][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n271));
   AO22CHD U4797 (.O(n3372), 
	.B2(n405), 
	.B1(\ram[174][6] ), 
	.A2(n14), 
	.A1(n271));
   AO22CHD U4798 (.O(n3373), 
	.B2(n405), 
	.B1(\ram[174][7] ), 
	.A2(n15), 
	.A1(n271));
   AO22CHD U4799 (.O(n3374), 
	.B2(n405), 
	.B1(\ram[174][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n271));
   AO22CHD U4800 (.O(n3375), 
	.B2(n405), 
	.B1(\ram[174][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n271));
   AO22CHD U4801 (.O(n3376), 
	.B2(n405), 
	.B1(\ram[174][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n271));
   AO22CHD U4802 (.O(n3377), 
	.B2(n405), 
	.B1(\ram[174][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n271));
   AO22CHD U4803 (.O(n3378), 
	.B2(n405), 
	.B1(\ram[174][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n271));
   AO22CHD U4804 (.O(n3379), 
	.B2(n405), 
	.B1(\ram[174][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n271));
   AO22CHD U4805 (.O(n3380), 
	.B2(n405), 
	.B1(\ram[174][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n271));
   AO22CHD U4806 (.O(n3381), 
	.B2(n405), 
	.B1(\ram[174][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n271));
   AO22CHD U4807 (.O(n3382), 
	.B2(n407), 
	.B1(\ram[175][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n273));
   AO22CHD U4808 (.O(n3383), 
	.B2(n407), 
	.B1(\ram[175][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n273));
   AO22CHD U4809 (.O(n3384), 
	.B2(n407), 
	.B1(\ram[175][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n273));
   AO22CHD U4810 (.O(n3385), 
	.B2(n407), 
	.B1(\ram[175][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n273));
   AO22CHD U4811 (.O(n3386), 
	.B2(n407), 
	.B1(\ram[175][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n273));
   AO22CHD U4812 (.O(n3387), 
	.B2(n407), 
	.B1(\ram[175][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n273));
   AO22CHD U4813 (.O(n3388), 
	.B2(n407), 
	.B1(\ram[175][6] ), 
	.A2(n14), 
	.A1(n273));
   AO22CHD U4814 (.O(n3389), 
	.B2(n407), 
	.B1(\ram[175][7] ), 
	.A2(n15), 
	.A1(n273));
   AO22CHD U4815 (.O(n3390), 
	.B2(n407), 
	.B1(\ram[175][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n273));
   AO22CHD U4816 (.O(n3391), 
	.B2(n407), 
	.B1(\ram[175][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n273));
   AO22CHD U4817 (.O(n3392), 
	.B2(n407), 
	.B1(\ram[175][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n273));
   AO22CHD U4818 (.O(n3393), 
	.B2(n407), 
	.B1(\ram[175][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n273));
   AO22CHD U4819 (.O(n3394), 
	.B2(n407), 
	.B1(\ram[175][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n273));
   AO22CHD U4820 (.O(n3395), 
	.B2(n407), 
	.B1(\ram[175][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n273));
   AO22CHD U4821 (.O(n3396), 
	.B2(n407), 
	.B1(\ram[175][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n273));
   AO22CHD U4822 (.O(n3397), 
	.B2(n407), 
	.B1(\ram[175][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n273));
   AO22CHD U4823 (.O(n3398), 
	.B2(n409), 
	.B1(\ram[176][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n275));
   AO22CHD U4824 (.O(n3399), 
	.B2(n409), 
	.B1(\ram[176][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n275));
   AO22CHD U4825 (.O(n3400), 
	.B2(n409), 
	.B1(\ram[176][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n275));
   AO22CHD U4826 (.O(n3401), 
	.B2(n409), 
	.B1(\ram[176][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n275));
   AO22CHD U4827 (.O(n3402), 
	.B2(n409), 
	.B1(\ram[176][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n275));
   AO22CHD U4828 (.O(n3403), 
	.B2(n409), 
	.B1(\ram[176][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n275));
   AO22CHD U4829 (.O(n3404), 
	.B2(n409), 
	.B1(\ram[176][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n275));
   AO22CHD U4830 (.O(n3405), 
	.B2(n409), 
	.B1(\ram[176][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n275));
   AO22CHD U4831 (.O(n3406), 
	.B2(n409), 
	.B1(\ram[176][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n275));
   AO22CHD U4832 (.O(n3407), 
	.B2(n409), 
	.B1(\ram[176][9] ), 
	.A2(n17), 
	.A1(n275));
   AO22CHD U4833 (.O(n3408), 
	.B2(n409), 
	.B1(\ram[176][10] ), 
	.A2(n18), 
	.A1(n275));
   AO22CHD U4834 (.O(n3409), 
	.B2(n409), 
	.B1(\ram[176][11] ), 
	.A2(n19), 
	.A1(n275));
   AO22CHD U4835 (.O(n3410), 
	.B2(n409), 
	.B1(\ram[176][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n275));
   AO22CHD U4836 (.O(n3411), 
	.B2(n409), 
	.B1(\ram[176][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n275));
   AO22CHD U4837 (.O(n3412), 
	.B2(n409), 
	.B1(\ram[176][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n275));
   AO22CHD U4838 (.O(n3413), 
	.B2(n409), 
	.B1(\ram[176][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n275));
   AO22CHD U4839 (.O(n3414), 
	.B2(n412), 
	.B1(\ram[177][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n277));
   AO22CHD U4840 (.O(n3415), 
	.B2(n412), 
	.B1(\ram[177][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n277));
   AO22CHD U4841 (.O(n3416), 
	.B2(n412), 
	.B1(\ram[177][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n277));
   AO22CHD U4842 (.O(n3417), 
	.B2(n412), 
	.B1(\ram[177][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n277));
   AO22CHD U4843 (.O(n3418), 
	.B2(n412), 
	.B1(\ram[177][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n277));
   AO22CHD U4844 (.O(n3419), 
	.B2(n412), 
	.B1(\ram[177][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n277));
   AO22CHD U4845 (.O(n3420), 
	.B2(n412), 
	.B1(\ram[177][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n277));
   AO22CHD U4846 (.O(n3421), 
	.B2(n412), 
	.B1(\ram[177][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n277));
   AO22CHD U4847 (.O(n3422), 
	.B2(n412), 
	.B1(\ram[177][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n277));
   AO22CHD U4848 (.O(n3423), 
	.B2(n412), 
	.B1(\ram[177][9] ), 
	.A2(n17), 
	.A1(n277));
   AO22CHD U4849 (.O(n3424), 
	.B2(n412), 
	.B1(\ram[177][10] ), 
	.A2(n18), 
	.A1(n277));
   AO22CHD U4850 (.O(n3425), 
	.B2(n412), 
	.B1(\ram[177][11] ), 
	.A2(n19), 
	.A1(n277));
   AO22CHD U4851 (.O(n3426), 
	.B2(n412), 
	.B1(\ram[177][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n277));
   AO22CHD U4852 (.O(n3427), 
	.B2(n412), 
	.B1(\ram[177][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n277));
   AO22CHD U4853 (.O(n3428), 
	.B2(n412), 
	.B1(\ram[177][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n277));
   AO22CHD U4854 (.O(n3429), 
	.B2(n412), 
	.B1(\ram[177][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n277));
   AO22CHD U4855 (.O(n3430), 
	.B2(n414), 
	.B1(\ram[178][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n278));
   AO22CHD U4856 (.O(n3431), 
	.B2(n414), 
	.B1(\ram[178][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n278));
   AO22CHD U4857 (.O(n3432), 
	.B2(n414), 
	.B1(\ram[178][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n278));
   AO22CHD U4858 (.O(n3433), 
	.B2(n414), 
	.B1(\ram[178][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n278));
   AO22CHD U4859 (.O(n3434), 
	.B2(n414), 
	.B1(\ram[178][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n278));
   AO22CHD U4860 (.O(n3435), 
	.B2(n414), 
	.B1(\ram[178][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n278));
   AO22CHD U4861 (.O(n3436), 
	.B2(n414), 
	.B1(\ram[178][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n278));
   AO22CHD U4862 (.O(n3437), 
	.B2(n414), 
	.B1(\ram[178][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n278));
   AO22CHD U4863 (.O(n3438), 
	.B2(n414), 
	.B1(\ram[178][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n278));
   AO22CHD U4864 (.O(n3439), 
	.B2(n414), 
	.B1(\ram[178][9] ), 
	.A2(n17), 
	.A1(n278));
   AO22CHD U4865 (.O(n3440), 
	.B2(n414), 
	.B1(\ram[178][10] ), 
	.A2(n18), 
	.A1(n278));
   AO22CHD U4866 (.O(n3441), 
	.B2(n414), 
	.B1(\ram[178][11] ), 
	.A2(n19), 
	.A1(n278));
   AO22CHD U4867 (.O(n3442), 
	.B2(n414), 
	.B1(\ram[178][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n278));
   AO22CHD U4868 (.O(n3443), 
	.B2(n414), 
	.B1(\ram[178][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n278));
   AO22CHD U4869 (.O(n3444), 
	.B2(n414), 
	.B1(\ram[178][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n278));
   AO22CHD U4870 (.O(n3445), 
	.B2(n414), 
	.B1(\ram[178][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n278));
   AO22CHD U4871 (.O(n3446), 
	.B2(n416), 
	.B1(\ram[179][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n280));
   AO22CHD U4872 (.O(n3447), 
	.B2(n416), 
	.B1(\ram[179][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n280));
   AO22CHD U4873 (.O(n3448), 
	.B2(n416), 
	.B1(\ram[179][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n280));
   AO22CHD U4874 (.O(n3449), 
	.B2(n416), 
	.B1(\ram[179][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n280));
   AO22CHD U4875 (.O(n3450), 
	.B2(n416), 
	.B1(\ram[179][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n280));
   AO22CHD U4876 (.O(n3451), 
	.B2(n416), 
	.B1(\ram[179][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n280));
   AO22CHD U4877 (.O(n3452), 
	.B2(n416), 
	.B1(\ram[179][6] ), 
	.A2(FE_OFN62_n14), 
	.A1(n280));
   AO22CHD U4878 (.O(n3453), 
	.B2(n416), 
	.B1(\ram[179][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n280));
   AO22CHD U4879 (.O(n3454), 
	.B2(n416), 
	.B1(\ram[179][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n280));
   AO22CHD U4880 (.O(n3455), 
	.B2(n416), 
	.B1(\ram[179][9] ), 
	.A2(n17), 
	.A1(n280));
   AO22CHD U4881 (.O(n3456), 
	.B2(n416), 
	.B1(\ram[179][10] ), 
	.A2(n18), 
	.A1(n280));
   AO22CHD U4882 (.O(n3457), 
	.B2(n416), 
	.B1(\ram[179][11] ), 
	.A2(n19), 
	.A1(n280));
   AO22CHD U4883 (.O(n3458), 
	.B2(n416), 
	.B1(\ram[179][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n280));
   AO22CHD U4884 (.O(n3459), 
	.B2(n416), 
	.B1(\ram[179][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n280));
   AO22CHD U4885 (.O(n3460), 
	.B2(n416), 
	.B1(\ram[179][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n280));
   AO22CHD U4886 (.O(n3461), 
	.B2(n416), 
	.B1(\ram[179][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n280));
   AO22CHD U4887 (.O(n3462), 
	.B2(n418), 
	.B1(\ram[180][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n282));
   AO22CHD U4888 (.O(n3463), 
	.B2(n418), 
	.B1(\ram[180][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n282));
   AO22CHD U4889 (.O(n3464), 
	.B2(n418), 
	.B1(\ram[180][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n282));
   AO22CHD U4890 (.O(n3465), 
	.B2(n418), 
	.B1(\ram[180][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n282));
   AO22CHD U4891 (.O(n3466), 
	.B2(n418), 
	.B1(\ram[180][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n282));
   AO22CHD U4892 (.O(n3467), 
	.B2(n418), 
	.B1(\ram[180][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n282));
   AO22CHD U4893 (.O(n3468), 
	.B2(n418), 
	.B1(\ram[180][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n282));
   AO22CHD U4894 (.O(n3469), 
	.B2(n418), 
	.B1(\ram[180][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n282));
   AO22CHD U4895 (.O(n3470), 
	.B2(n418), 
	.B1(\ram[180][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n282));
   AO22CHD U4896 (.O(n3471), 
	.B2(n418), 
	.B1(\ram[180][9] ), 
	.A2(n17), 
	.A1(n282));
   AO22CHD U4897 (.O(n3472), 
	.B2(n418), 
	.B1(\ram[180][10] ), 
	.A2(n18), 
	.A1(n282));
   AO22CHD U4898 (.O(n3473), 
	.B2(n418), 
	.B1(\ram[180][11] ), 
	.A2(n19), 
	.A1(n282));
   AO22CHD U4899 (.O(n3474), 
	.B2(n418), 
	.B1(\ram[180][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n282));
   AO22CHD U4900 (.O(n3475), 
	.B2(n418), 
	.B1(\ram[180][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n282));
   AO22CHD U4901 (.O(n3476), 
	.B2(n418), 
	.B1(\ram[180][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n282));
   AO22CHD U4902 (.O(n3477), 
	.B2(n418), 
	.B1(\ram[180][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n282));
   AO22CHD U4903 (.O(n3478), 
	.B2(n420), 
	.B1(\ram[181][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n284));
   AO22CHD U4904 (.O(n3479), 
	.B2(n420), 
	.B1(\ram[181][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n284));
   AO22CHD U4905 (.O(n3480), 
	.B2(n420), 
	.B1(\ram[181][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n284));
   AO22CHD U4906 (.O(n3481), 
	.B2(n420), 
	.B1(\ram[181][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n284));
   AO22CHD U4907 (.O(n3482), 
	.B2(n420), 
	.B1(\ram[181][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n284));
   AO22CHD U4908 (.O(n3483), 
	.B2(n420), 
	.B1(\ram[181][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n284));
   AO22CHD U4909 (.O(n3484), 
	.B2(n420), 
	.B1(\ram[181][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n284));
   AO22CHD U4910 (.O(n3485), 
	.B2(n420), 
	.B1(\ram[181][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n284));
   AO22CHD U4911 (.O(n3486), 
	.B2(n420), 
	.B1(\ram[181][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n284));
   AO22CHD U4912 (.O(n3487), 
	.B2(n420), 
	.B1(\ram[181][9] ), 
	.A2(n17), 
	.A1(n284));
   AO22CHD U4913 (.O(n3488), 
	.B2(n420), 
	.B1(\ram[181][10] ), 
	.A2(n18), 
	.A1(n284));
   AO22CHD U4914 (.O(n3489), 
	.B2(n420), 
	.B1(\ram[181][11] ), 
	.A2(n19), 
	.A1(n284));
   AO22CHD U4915 (.O(n3490), 
	.B2(n420), 
	.B1(\ram[181][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n284));
   AO22CHD U4916 (.O(n3491), 
	.B2(n420), 
	.B1(\ram[181][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n284));
   AO22CHD U4917 (.O(n3492), 
	.B2(n420), 
	.B1(\ram[181][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n284));
   AO22CHD U4918 (.O(n3493), 
	.B2(n420), 
	.B1(\ram[181][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n284));
   AO22CHD U4919 (.O(n3494), 
	.B2(n422), 
	.B1(\ram[182][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n286));
   AO22CHD U4920 (.O(n3495), 
	.B2(n422), 
	.B1(\ram[182][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n286));
   AO22CHD U4921 (.O(n3496), 
	.B2(n422), 
	.B1(\ram[182][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n286));
   AO22CHD U4922 (.O(n3497), 
	.B2(n422), 
	.B1(\ram[182][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n286));
   AO22CHD U4923 (.O(n3498), 
	.B2(n422), 
	.B1(\ram[182][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n286));
   AO22CHD U4924 (.O(n3499), 
	.B2(n422), 
	.B1(\ram[182][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n286));
   AO22CHD U4925 (.O(n3500), 
	.B2(n422), 
	.B1(\ram[182][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n286));
   AO22CHD U4926 (.O(n3501), 
	.B2(n422), 
	.B1(\ram[182][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n286));
   AO22CHD U4927 (.O(n3502), 
	.B2(n422), 
	.B1(\ram[182][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n286));
   AO22CHD U4928 (.O(n3503), 
	.B2(n422), 
	.B1(\ram[182][9] ), 
	.A2(n17), 
	.A1(n286));
   AO22CHD U4929 (.O(n3504), 
	.B2(n422), 
	.B1(\ram[182][10] ), 
	.A2(n18), 
	.A1(n286));
   AO22CHD U4930 (.O(n3505), 
	.B2(n422), 
	.B1(\ram[182][11] ), 
	.A2(n19), 
	.A1(n286));
   AO22CHD U4931 (.O(n3506), 
	.B2(n422), 
	.B1(\ram[182][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n286));
   AO22CHD U4932 (.O(n3507), 
	.B2(n422), 
	.B1(\ram[182][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n286));
   AO22CHD U4933 (.O(n3508), 
	.B2(n422), 
	.B1(\ram[182][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n286));
   AO22CHD U4934 (.O(n3509), 
	.B2(n422), 
	.B1(\ram[182][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n286));
   AO22CHD U4935 (.O(n3510), 
	.B2(n424), 
	.B1(\ram[183][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n288));
   AO22CHD U4936 (.O(n3511), 
	.B2(n424), 
	.B1(\ram[183][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n288));
   AO22CHD U4937 (.O(n3512), 
	.B2(n424), 
	.B1(\ram[183][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n288));
   AO22CHD U4938 (.O(n3513), 
	.B2(n424), 
	.B1(\ram[183][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n288));
   AO22CHD U4939 (.O(n3514), 
	.B2(n424), 
	.B1(\ram[183][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n288));
   AO22CHD U4940 (.O(n3515), 
	.B2(n424), 
	.B1(\ram[183][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n288));
   AO22CHD U4941 (.O(n3516), 
	.B2(n424), 
	.B1(\ram[183][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n288));
   AO22CHD U4942 (.O(n3517), 
	.B2(n424), 
	.B1(\ram[183][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n288));
   AO22CHD U4943 (.O(n3518), 
	.B2(n424), 
	.B1(\ram[183][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n288));
   AO22CHD U4944 (.O(n3519), 
	.B2(n424), 
	.B1(\ram[183][9] ), 
	.A2(n17), 
	.A1(n288));
   AO22CHD U4945 (.O(n3520), 
	.B2(n424), 
	.B1(\ram[183][10] ), 
	.A2(n18), 
	.A1(n288));
   AO22CHD U4946 (.O(n3521), 
	.B2(n424), 
	.B1(\ram[183][11] ), 
	.A2(n19), 
	.A1(n288));
   AO22CHD U4947 (.O(n3522), 
	.B2(n424), 
	.B1(\ram[183][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n288));
   AO22CHD U4948 (.O(n3523), 
	.B2(n424), 
	.B1(\ram[183][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n288));
   AO22CHD U4949 (.O(n3524), 
	.B2(n424), 
	.B1(\ram[183][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n288));
   AO22CHD U4950 (.O(n3525), 
	.B2(n424), 
	.B1(\ram[183][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n288));
   AO22CHD U4951 (.O(n3526), 
	.B2(n426), 
	.B1(\ram[184][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n290));
   AO22CHD U4952 (.O(n3527), 
	.B2(n426), 
	.B1(\ram[184][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n290));
   AO22CHD U4953 (.O(n3528), 
	.B2(n426), 
	.B1(\ram[184][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n290));
   AO22CHD U4954 (.O(n3529), 
	.B2(n426), 
	.B1(\ram[184][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n290));
   AO22CHD U4955 (.O(n3530), 
	.B2(n426), 
	.B1(\ram[184][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n290));
   AO22CHD U4956 (.O(n3531), 
	.B2(n426), 
	.B1(\ram[184][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n290));
   AO22CHD U4957 (.O(n3532), 
	.B2(n426), 
	.B1(\ram[184][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n290));
   AO22CHD U4958 (.O(n3533), 
	.B2(n426), 
	.B1(\ram[184][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n290));
   AO22CHD U4959 (.O(n3534), 
	.B2(n426), 
	.B1(\ram[184][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n290));
   AO22CHD U4960 (.O(n3535), 
	.B2(n426), 
	.B1(\ram[184][9] ), 
	.A2(n17), 
	.A1(n290));
   AO22CHD U4961 (.O(n3536), 
	.B2(n426), 
	.B1(\ram[184][10] ), 
	.A2(n18), 
	.A1(n290));
   AO22CHD U4962 (.O(n3537), 
	.B2(n426), 
	.B1(\ram[184][11] ), 
	.A2(n19), 
	.A1(n290));
   AO22CHD U4963 (.O(n3538), 
	.B2(n426), 
	.B1(\ram[184][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n290));
   AO22CHD U4964 (.O(n3539), 
	.B2(n426), 
	.B1(\ram[184][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n290));
   AO22CHD U4965 (.O(n3540), 
	.B2(n426), 
	.B1(\ram[184][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n290));
   AO22CHD U4966 (.O(n3541), 
	.B2(n426), 
	.B1(\ram[184][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n290));
   AO22CHD U4967 (.O(n3542), 
	.B2(n428), 
	.B1(\ram[185][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n292));
   AO22CHD U4968 (.O(n3543), 
	.B2(n428), 
	.B1(\ram[185][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n292));
   AO22CHD U4969 (.O(n3544), 
	.B2(n428), 
	.B1(\ram[185][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n292));
   AO22CHD U4970 (.O(n3545), 
	.B2(n428), 
	.B1(\ram[185][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n292));
   AO22CHD U4971 (.O(n3546), 
	.B2(n428), 
	.B1(\ram[185][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n292));
   AO22CHD U4972 (.O(n3547), 
	.B2(n428), 
	.B1(\ram[185][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n292));
   AO22CHD U4973 (.O(n3548), 
	.B2(n428), 
	.B1(\ram[185][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n292));
   AO22CHD U4974 (.O(n3549), 
	.B2(n428), 
	.B1(\ram[185][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n292));
   AO22CHD U4975 (.O(n3550), 
	.B2(n428), 
	.B1(\ram[185][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n292));
   AO22CHD U4976 (.O(n3551), 
	.B2(n428), 
	.B1(\ram[185][9] ), 
	.A2(n17), 
	.A1(n292));
   AO22CHD U4977 (.O(n3552), 
	.B2(n428), 
	.B1(\ram[185][10] ), 
	.A2(n18), 
	.A1(n292));
   AO22CHD U4978 (.O(n3553), 
	.B2(n428), 
	.B1(\ram[185][11] ), 
	.A2(n19), 
	.A1(n292));
   AO22CHD U4979 (.O(n3554), 
	.B2(n428), 
	.B1(\ram[185][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n292));
   AO22CHD U4980 (.O(n3555), 
	.B2(n428), 
	.B1(\ram[185][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n292));
   AO22CHD U4981 (.O(n3556), 
	.B2(n428), 
	.B1(\ram[185][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n292));
   AO22CHD U4982 (.O(n3557), 
	.B2(n428), 
	.B1(\ram[185][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n292));
   AO22CHD U4983 (.O(n3558), 
	.B2(n430), 
	.B1(\ram[186][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n294));
   AO22CHD U4984 (.O(n3559), 
	.B2(n430), 
	.B1(\ram[186][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n294));
   AO22CHD U4985 (.O(n3560), 
	.B2(n430), 
	.B1(\ram[186][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n294));
   AO22CHD U4986 (.O(n3561), 
	.B2(n430), 
	.B1(\ram[186][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n294));
   AO22CHD U4987 (.O(n3562), 
	.B2(n430), 
	.B1(\ram[186][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n294));
   AO22CHD U4988 (.O(n3563), 
	.B2(n430), 
	.B1(\ram[186][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n294));
   AO22CHD U4989 (.O(n3564), 
	.B2(n430), 
	.B1(\ram[186][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n294));
   AO22CHD U4990 (.O(n3565), 
	.B2(n430), 
	.B1(\ram[186][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n294));
   AO22CHD U4991 (.O(n3566), 
	.B2(n430), 
	.B1(\ram[186][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n294));
   AO22CHD U4992 (.O(n3567), 
	.B2(n430), 
	.B1(\ram[186][9] ), 
	.A2(n17), 
	.A1(n294));
   AO22CHD U4993 (.O(n3568), 
	.B2(n430), 
	.B1(\ram[186][10] ), 
	.A2(n18), 
	.A1(n294));
   AO22CHD U4994 (.O(n3569), 
	.B2(n430), 
	.B1(\ram[186][11] ), 
	.A2(n19), 
	.A1(n294));
   AO22CHD U4995 (.O(n3570), 
	.B2(n430), 
	.B1(\ram[186][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n294));
   AO22CHD U4996 (.O(n3571), 
	.B2(n430), 
	.B1(\ram[186][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n294));
   AO22CHD U4997 (.O(n3572), 
	.B2(n430), 
	.B1(\ram[186][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n294));
   AO22CHD U4998 (.O(n3573), 
	.B2(n430), 
	.B1(\ram[186][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n294));
   AO22CHD U4999 (.O(n3574), 
	.B2(n432), 
	.B1(\ram[187][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n296));
   AO22CHD U5000 (.O(n3575), 
	.B2(n432), 
	.B1(\ram[187][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n296));
   AO22CHD U5001 (.O(n3576), 
	.B2(n432), 
	.B1(\ram[187][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n296));
   AO22CHD U5002 (.O(n3577), 
	.B2(n432), 
	.B1(\ram[187][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n296));
   AO22CHD U5003 (.O(n3578), 
	.B2(n432), 
	.B1(\ram[187][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n296));
   AO22CHD U5004 (.O(n3579), 
	.B2(n432), 
	.B1(\ram[187][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n296));
   AO22CHD U5005 (.O(n3580), 
	.B2(n432), 
	.B1(\ram[187][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n296));
   AO22CHD U5006 (.O(n3581), 
	.B2(n432), 
	.B1(\ram[187][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n296));
   AO22CHD U5007 (.O(n3582), 
	.B2(n432), 
	.B1(\ram[187][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n296));
   AO22CHD U5008 (.O(n3583), 
	.B2(n432), 
	.B1(\ram[187][9] ), 
	.A2(n17), 
	.A1(n296));
   AO22CHD U5009 (.O(n3584), 
	.B2(n432), 
	.B1(\ram[187][10] ), 
	.A2(n18), 
	.A1(n296));
   AO22CHD U5010 (.O(n3585), 
	.B2(n432), 
	.B1(\ram[187][11] ), 
	.A2(n19), 
	.A1(n296));
   AO22CHD U5011 (.O(n3586), 
	.B2(n432), 
	.B1(\ram[187][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n296));
   AO22CHD U5012 (.O(n3587), 
	.B2(n432), 
	.B1(\ram[187][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n296));
   AO22CHD U5013 (.O(n3588), 
	.B2(n432), 
	.B1(\ram[187][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n296));
   AO22CHD U5014 (.O(n3589), 
	.B2(n432), 
	.B1(\ram[187][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n296));
   AO22CHD U5015 (.O(n3590), 
	.B2(n434), 
	.B1(\ram[188][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n298));
   AO22CHD U5016 (.O(n3591), 
	.B2(n434), 
	.B1(\ram[188][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n298));
   AO22CHD U5017 (.O(n3592), 
	.B2(n434), 
	.B1(\ram[188][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n298));
   AO22CHD U5018 (.O(n3593), 
	.B2(n434), 
	.B1(\ram[188][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n298));
   AO22CHD U5019 (.O(n3594), 
	.B2(n434), 
	.B1(\ram[188][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n298));
   AO22CHD U5020 (.O(n3595), 
	.B2(n434), 
	.B1(\ram[188][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n298));
   AO22CHD U5021 (.O(n3596), 
	.B2(n434), 
	.B1(\ram[188][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n298));
   AO22CHD U5022 (.O(n3597), 
	.B2(n434), 
	.B1(\ram[188][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n298));
   AO22CHD U5023 (.O(n3598), 
	.B2(n434), 
	.B1(\ram[188][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n298));
   AO22CHD U5024 (.O(n3599), 
	.B2(n434), 
	.B1(\ram[188][9] ), 
	.A2(n17), 
	.A1(n298));
   AO22CHD U5025 (.O(n3600), 
	.B2(n434), 
	.B1(\ram[188][10] ), 
	.A2(n18), 
	.A1(n298));
   AO22CHD U5026 (.O(n3601), 
	.B2(n434), 
	.B1(\ram[188][11] ), 
	.A2(n19), 
	.A1(n298));
   AO22CHD U5027 (.O(n3602), 
	.B2(n434), 
	.B1(\ram[188][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n298));
   AO22CHD U5028 (.O(n3603), 
	.B2(n434), 
	.B1(\ram[188][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n298));
   AO22CHD U5029 (.O(n3604), 
	.B2(n434), 
	.B1(\ram[188][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n298));
   AO22CHD U5030 (.O(n3605), 
	.B2(n434), 
	.B1(\ram[188][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n298));
   AO22CHD U5031 (.O(n3606), 
	.B2(n436), 
	.B1(\ram[189][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n300));
   AO22CHD U5032 (.O(n3607), 
	.B2(n436), 
	.B1(\ram[189][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n300));
   AO22CHD U5033 (.O(n3608), 
	.B2(n436), 
	.B1(\ram[189][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n300));
   AO22CHD U5034 (.O(n3609), 
	.B2(n436), 
	.B1(\ram[189][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n300));
   AO22CHD U5035 (.O(n3610), 
	.B2(n436), 
	.B1(\ram[189][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n300));
   AO22CHD U5036 (.O(n3611), 
	.B2(n436), 
	.B1(\ram[189][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n300));
   AO22CHD U5037 (.O(n3612), 
	.B2(n436), 
	.B1(\ram[189][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n300));
   AO22CHD U5038 (.O(n3613), 
	.B2(n436), 
	.B1(\ram[189][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n300));
   AO22CHD U5039 (.O(n3614), 
	.B2(n436), 
	.B1(\ram[189][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n300));
   AO22CHD U5040 (.O(n3615), 
	.B2(n436), 
	.B1(\ram[189][9] ), 
	.A2(n17), 
	.A1(n300));
   AO22CHD U5041 (.O(n3616), 
	.B2(n436), 
	.B1(\ram[189][10] ), 
	.A2(n18), 
	.A1(n300));
   AO22CHD U5042 (.O(n3617), 
	.B2(n436), 
	.B1(\ram[189][11] ), 
	.A2(n19), 
	.A1(n300));
   AO22CHD U5043 (.O(n3618), 
	.B2(n436), 
	.B1(\ram[189][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n300));
   AO22CHD U5044 (.O(n3619), 
	.B2(n436), 
	.B1(\ram[189][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n300));
   AO22CHD U5045 (.O(n3620), 
	.B2(n436), 
	.B1(\ram[189][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n300));
   AO22CHD U5046 (.O(n3621), 
	.B2(n436), 
	.B1(\ram[189][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n300));
   AO22CHD U5047 (.O(n3622), 
	.B2(n438), 
	.B1(\ram[190][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n302));
   AO22CHD U5048 (.O(n3623), 
	.B2(n438), 
	.B1(\ram[190][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n302));
   AO22CHD U5049 (.O(n3624), 
	.B2(n438), 
	.B1(\ram[190][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n302));
   AO22CHD U5050 (.O(n3625), 
	.B2(n438), 
	.B1(\ram[190][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n302));
   AO22CHD U5051 (.O(n3626), 
	.B2(n438), 
	.B1(\ram[190][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n302));
   AO22CHD U5052 (.O(n3627), 
	.B2(n438), 
	.B1(\ram[190][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n302));
   AO22CHD U5053 (.O(n3628), 
	.B2(n438), 
	.B1(\ram[190][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n302));
   AO22CHD U5054 (.O(n3629), 
	.B2(n438), 
	.B1(\ram[190][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n302));
   AO22CHD U5055 (.O(n3630), 
	.B2(n438), 
	.B1(\ram[190][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n302));
   AO22CHD U5056 (.O(n3631), 
	.B2(n438), 
	.B1(\ram[190][9] ), 
	.A2(n17), 
	.A1(n302));
   AO22CHD U5057 (.O(n3632), 
	.B2(n438), 
	.B1(\ram[190][10] ), 
	.A2(n18), 
	.A1(n302));
   AO22CHD U5058 (.O(n3633), 
	.B2(n438), 
	.B1(\ram[190][11] ), 
	.A2(n19), 
	.A1(n302));
   AO22CHD U5059 (.O(n3634), 
	.B2(n438), 
	.B1(\ram[190][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n302));
   AO22CHD U5060 (.O(n3635), 
	.B2(n438), 
	.B1(\ram[190][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n302));
   AO22CHD U5061 (.O(n3636), 
	.B2(n438), 
	.B1(\ram[190][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n302));
   AO22CHD U5062 (.O(n3637), 
	.B2(n438), 
	.B1(\ram[190][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n302));
   AO22CHD U5063 (.O(n3638), 
	.B2(n440), 
	.B1(\ram[191][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n304));
   AO22CHD U5064 (.O(n3639), 
	.B2(n440), 
	.B1(\ram[191][1] ), 
	.A2(FE_OFN46_n9), 
	.A1(n304));
   AO22CHD U5065 (.O(n3640), 
	.B2(n440), 
	.B1(\ram[191][2] ), 
	.A2(FE_OFN49_n10), 
	.A1(n304));
   AO22CHD U5066 (.O(n3641), 
	.B2(n440), 
	.B1(\ram[191][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n304));
   AO22CHD U5067 (.O(n3642), 
	.B2(n440), 
	.B1(\ram[191][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n304));
   AO22CHD U5068 (.O(n3643), 
	.B2(n440), 
	.B1(\ram[191][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n304));
   AO22CHD U5069 (.O(n3644), 
	.B2(n440), 
	.B1(\ram[191][6] ), 
	.A2(FE_OFN61_n14), 
	.A1(n304));
   AO22CHD U5070 (.O(n3645), 
	.B2(n440), 
	.B1(\ram[191][7] ), 
	.A2(FE_OFN63_n15), 
	.A1(n304));
   AO22CHD U5071 (.O(n3646), 
	.B2(n440), 
	.B1(\ram[191][8] ), 
	.A2(FE_OFN68_n16), 
	.A1(n304));
   AO22CHD U5072 (.O(n3647), 
	.B2(n440), 
	.B1(\ram[191][9] ), 
	.A2(n17), 
	.A1(n304));
   AO22CHD U5073 (.O(n3648), 
	.B2(n440), 
	.B1(\ram[191][10] ), 
	.A2(n18), 
	.A1(n304));
   AO22CHD U5074 (.O(n3649), 
	.B2(n440), 
	.B1(\ram[191][11] ), 
	.A2(n19), 
	.A1(n304));
   AO22CHD U5075 (.O(n3650), 
	.B2(n440), 
	.B1(\ram[191][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n304));
   AO22CHD U5076 (.O(n3651), 
	.B2(n440), 
	.B1(\ram[191][13] ), 
	.A2(FE_OFN85_n21), 
	.A1(n304));
   AO22CHD U5077 (.O(n3652), 
	.B2(n440), 
	.B1(\ram[191][14] ), 
	.A2(FE_OFN88_n22), 
	.A1(n304));
   AO22CHD U5078 (.O(n3653), 
	.B2(n440), 
	.B1(\ram[191][15] ), 
	.A2(FE_OFN91_n23), 
	.A1(n304));
   AO22CHD U5079 (.O(n3654), 
	.B2(n442), 
	.B1(\ram[192][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n306));
   AO22CHD U5080 (.O(n3655), 
	.B2(n442), 
	.B1(\ram[192][1] ), 
	.A2(n9), 
	.A1(n306));
   AO22CHD U5081 (.O(n3656), 
	.B2(n442), 
	.B1(\ram[192][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n306));
   AO22CHD U5082 (.O(n3657), 
	.B2(n442), 
	.B1(\ram[192][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n306));
   AO22CHD U5083 (.O(n3658), 
	.B2(n442), 
	.B1(\ram[192][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n306));
   AO22CHD U5084 (.O(n3659), 
	.B2(n442), 
	.B1(\ram[192][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n306));
   AO22CHD U5085 (.O(n3660), 
	.B2(n442), 
	.B1(\ram[192][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n306));
   AO22CHD U5086 (.O(n3661), 
	.B2(n442), 
	.B1(\ram[192][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n306));
   AO22CHD U5087 (.O(n3662), 
	.B2(n442), 
	.B1(\ram[192][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n306));
   AO22CHD U5088 (.O(n3663), 
	.B2(n442), 
	.B1(\ram[192][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n306));
   AO22CHD U5089 (.O(n3664), 
	.B2(n442), 
	.B1(\ram[192][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n306));
   AO22CHD U5090 (.O(n3665), 
	.B2(n442), 
	.B1(\ram[192][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n306));
   AO22CHD U5091 (.O(n3666), 
	.B2(n442), 
	.B1(\ram[192][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n306));
   AO22CHD U5092 (.O(n3667), 
	.B2(n442), 
	.B1(\ram[192][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n306));
   AO22CHD U5093 (.O(n3668), 
	.B2(n442), 
	.B1(\ram[192][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n306));
   AO22CHD U5094 (.O(n3669), 
	.B2(n442), 
	.B1(\ram[192][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n306));
   AO22CHD U5095 (.O(n3670), 
	.B2(n445), 
	.B1(\ram[193][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n308));
   AO22CHD U5096 (.O(n3671), 
	.B2(n445), 
	.B1(\ram[193][1] ), 
	.A2(n9), 
	.A1(n308));
   AO22CHD U5097 (.O(n3672), 
	.B2(n445), 
	.B1(\ram[193][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n308));
   AO22CHD U5098 (.O(n3673), 
	.B2(n445), 
	.B1(\ram[193][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n308));
   AO22CHD U5099 (.O(n3674), 
	.B2(n445), 
	.B1(\ram[193][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n308));
   AO22CHD U5100 (.O(n3675), 
	.B2(n445), 
	.B1(\ram[193][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n308));
   AO22CHD U5101 (.O(n3676), 
	.B2(n445), 
	.B1(\ram[193][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n308));
   AO22CHD U5102 (.O(n3677), 
	.B2(n445), 
	.B1(\ram[193][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n308));
   AO22CHD U5103 (.O(n3678), 
	.B2(n445), 
	.B1(\ram[193][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n308));
   AO22CHD U5104 (.O(n3679), 
	.B2(n445), 
	.B1(\ram[193][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n308));
   AO22CHD U5105 (.O(n3680), 
	.B2(n445), 
	.B1(\ram[193][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n308));
   AO22CHD U5106 (.O(n3681), 
	.B2(n445), 
	.B1(\ram[193][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n308));
   AO22CHD U5107 (.O(n3682), 
	.B2(n445), 
	.B1(\ram[193][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n308));
   AO22CHD U5108 (.O(n3683), 
	.B2(n445), 
	.B1(\ram[193][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n308));
   AO22CHD U5109 (.O(n3684), 
	.B2(n445), 
	.B1(\ram[193][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n308));
   AO22CHD U5110 (.O(n3685), 
	.B2(n445), 
	.B1(\ram[193][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n308));
   AO22CHD U5111 (.O(n3686), 
	.B2(n447), 
	.B1(\ram[194][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n310));
   AO22CHD U5112 (.O(n3687), 
	.B2(n447), 
	.B1(\ram[194][1] ), 
	.A2(n9), 
	.A1(n310));
   AO22CHD U5113 (.O(n3688), 
	.B2(n447), 
	.B1(\ram[194][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n310));
   AO22CHD U5114 (.O(n3689), 
	.B2(n447), 
	.B1(\ram[194][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n310));
   AO22CHD U5115 (.O(n3690), 
	.B2(n447), 
	.B1(\ram[194][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n310));
   AO22CHD U5116 (.O(n3691), 
	.B2(n447), 
	.B1(\ram[194][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n310));
   AO22CHD U5117 (.O(n3692), 
	.B2(n447), 
	.B1(\ram[194][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n310));
   AO22CHD U5118 (.O(n3693), 
	.B2(n447), 
	.B1(\ram[194][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n310));
   AO22CHD U5119 (.O(n3694), 
	.B2(n447), 
	.B1(\ram[194][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n310));
   AO22CHD U5120 (.O(n3695), 
	.B2(n447), 
	.B1(\ram[194][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n310));
   AO22CHD U5121 (.O(n3696), 
	.B2(n447), 
	.B1(\ram[194][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n310));
   AO22CHD U5122 (.O(n3697), 
	.B2(n447), 
	.B1(\ram[194][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n310));
   AO22CHD U5123 (.O(n3698), 
	.B2(n447), 
	.B1(\ram[194][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n310));
   AO22CHD U5124 (.O(n3699), 
	.B2(n447), 
	.B1(\ram[194][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n310));
   AO22CHD U5125 (.O(n3700), 
	.B2(n447), 
	.B1(\ram[194][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n310));
   AO22CHD U5126 (.O(n3701), 
	.B2(n447), 
	.B1(\ram[194][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n310));
   AO22CHD U5127 (.O(n3702), 
	.B2(n449), 
	.B1(\ram[195][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n311));
   AO22CHD U5128 (.O(n3703), 
	.B2(n449), 
	.B1(\ram[195][1] ), 
	.A2(n9), 
	.A1(n311));
   AO22CHD U5129 (.O(n3704), 
	.B2(n449), 
	.B1(\ram[195][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n311));
   AO22CHD U5130 (.O(n3705), 
	.B2(n449), 
	.B1(\ram[195][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n311));
   AO22CHD U5131 (.O(n3706), 
	.B2(n449), 
	.B1(\ram[195][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n311));
   AO22CHD U5132 (.O(n3707), 
	.B2(n449), 
	.B1(\ram[195][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n311));
   AO22CHD U5133 (.O(n3708), 
	.B2(n449), 
	.B1(\ram[195][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n311));
   AO22CHD U5134 (.O(n3709), 
	.B2(n449), 
	.B1(\ram[195][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n311));
   AO22CHD U5135 (.O(n3710), 
	.B2(n449), 
	.B1(\ram[195][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n311));
   AO22CHD U5136 (.O(n3711), 
	.B2(n449), 
	.B1(\ram[195][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n311));
   AO22CHD U5137 (.O(n3712), 
	.B2(n449), 
	.B1(\ram[195][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n311));
   AO22CHD U5138 (.O(n3713), 
	.B2(n449), 
	.B1(\ram[195][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n311));
   AO22CHD U5139 (.O(n3714), 
	.B2(n449), 
	.B1(\ram[195][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n311));
   AO22CHD U5140 (.O(n3715), 
	.B2(n449), 
	.B1(\ram[195][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n311));
   AO22CHD U5141 (.O(n3716), 
	.B2(n449), 
	.B1(\ram[195][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n311));
   AO22CHD U5142 (.O(n3717), 
	.B2(n449), 
	.B1(\ram[195][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n311));
   AO22CHD U5143 (.O(n3718), 
	.B2(n451), 
	.B1(\ram[196][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n313));
   AO22CHD U5144 (.O(n3719), 
	.B2(n451), 
	.B1(\ram[196][1] ), 
	.A2(n9), 
	.A1(n313));
   AO22CHD U5145 (.O(n3720), 
	.B2(n451), 
	.B1(\ram[196][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n313));
   AO22CHD U5146 (.O(n3721), 
	.B2(n451), 
	.B1(\ram[196][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n313));
   AO22CHD U5147 (.O(n3722), 
	.B2(n451), 
	.B1(\ram[196][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n313));
   AO22CHD U5148 (.O(n3723), 
	.B2(n451), 
	.B1(\ram[196][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n313));
   AO22CHD U5149 (.O(n3724), 
	.B2(n451), 
	.B1(\ram[196][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n313));
   AO22CHD U5150 (.O(n3725), 
	.B2(n451), 
	.B1(\ram[196][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n313));
   AO22CHD U5151 (.O(n3726), 
	.B2(n451), 
	.B1(\ram[196][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n313));
   AO22CHD U5152 (.O(n3727), 
	.B2(n451), 
	.B1(\ram[196][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n313));
   AO22CHD U5153 (.O(n3728), 
	.B2(n451), 
	.B1(\ram[196][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n313));
   AO22CHD U5154 (.O(n3729), 
	.B2(n451), 
	.B1(\ram[196][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n313));
   AO22CHD U5155 (.O(n3730), 
	.B2(n451), 
	.B1(\ram[196][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n313));
   AO22CHD U5156 (.O(n3731), 
	.B2(n451), 
	.B1(\ram[196][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n313));
   AO22CHD U5157 (.O(n3732), 
	.B2(n451), 
	.B1(\ram[196][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n313));
   AO22CHD U5158 (.O(n3733), 
	.B2(n451), 
	.B1(\ram[196][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n313));
   AO22CHD U5159 (.O(n3734), 
	.B2(n453), 
	.B1(\ram[197][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n315));
   AO22CHD U5160 (.O(n3735), 
	.B2(n453), 
	.B1(\ram[197][1] ), 
	.A2(n9), 
	.A1(n315));
   AO22CHD U5161 (.O(n3736), 
	.B2(n453), 
	.B1(\ram[197][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n315));
   AO22CHD U5162 (.O(n3737), 
	.B2(n453), 
	.B1(\ram[197][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n315));
   AO22CHD U5163 (.O(n3738), 
	.B2(n453), 
	.B1(\ram[197][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n315));
   AO22CHD U5164 (.O(n3739), 
	.B2(n453), 
	.B1(\ram[197][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n315));
   AO22CHD U5165 (.O(n3740), 
	.B2(n453), 
	.B1(\ram[197][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n315));
   AO22CHD U5166 (.O(n3741), 
	.B2(n453), 
	.B1(\ram[197][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n315));
   AO22CHD U5167 (.O(n3742), 
	.B2(n453), 
	.B1(\ram[197][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n315));
   AO22CHD U5168 (.O(n3743), 
	.B2(n453), 
	.B1(\ram[197][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n315));
   AO22CHD U5169 (.O(n3744), 
	.B2(n453), 
	.B1(\ram[197][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n315));
   AO22CHD U5170 (.O(n3745), 
	.B2(n453), 
	.B1(\ram[197][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n315));
   AO22CHD U5171 (.O(n3746), 
	.B2(n453), 
	.B1(\ram[197][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n315));
   AO22CHD U5172 (.O(n3747), 
	.B2(n453), 
	.B1(\ram[197][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n315));
   AO22CHD U5173 (.O(n3748), 
	.B2(n453), 
	.B1(\ram[197][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n315));
   AO22CHD U5174 (.O(n3749), 
	.B2(n453), 
	.B1(\ram[197][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n315));
   AO22CHD U5175 (.O(n3750), 
	.B2(n455), 
	.B1(\ram[198][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n317));
   AO22CHD U5176 (.O(n3751), 
	.B2(n455), 
	.B1(\ram[198][1] ), 
	.A2(n9), 
	.A1(n317));
   AO22CHD U5177 (.O(n3752), 
	.B2(n455), 
	.B1(\ram[198][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n317));
   AO22CHD U5178 (.O(n3753), 
	.B2(n455), 
	.B1(\ram[198][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n317));
   AO22CHD U5179 (.O(n3754), 
	.B2(n455), 
	.B1(\ram[198][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n317));
   AO22CHD U5180 (.O(n3755), 
	.B2(n455), 
	.B1(\ram[198][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n317));
   AO22CHD U5181 (.O(n3756), 
	.B2(n455), 
	.B1(\ram[198][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n317));
   AO22CHD U5182 (.O(n3757), 
	.B2(n455), 
	.B1(\ram[198][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n317));
   AO22CHD U5183 (.O(n3758), 
	.B2(n455), 
	.B1(\ram[198][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n317));
   AO22CHD U5184 (.O(n3759), 
	.B2(n455), 
	.B1(\ram[198][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n317));
   AO22CHD U5185 (.O(n3760), 
	.B2(n455), 
	.B1(\ram[198][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n317));
   AO22CHD U5186 (.O(n3761), 
	.B2(n455), 
	.B1(\ram[198][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n317));
   AO22CHD U5187 (.O(n3762), 
	.B2(n455), 
	.B1(\ram[198][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n317));
   AO22CHD U5188 (.O(n3763), 
	.B2(n455), 
	.B1(\ram[198][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n317));
   AO22CHD U5189 (.O(n3764), 
	.B2(n455), 
	.B1(\ram[198][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n317));
   AO22CHD U5190 (.O(n3765), 
	.B2(n455), 
	.B1(\ram[198][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n317));
   AO22CHD U5191 (.O(n3766), 
	.B2(n457), 
	.B1(\ram[199][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n319));
   AO22CHD U5192 (.O(n3767), 
	.B2(n457), 
	.B1(\ram[199][1] ), 
	.A2(n9), 
	.A1(n319));
   AO22CHD U5193 (.O(n3768), 
	.B2(n457), 
	.B1(\ram[199][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n319));
   AO22CHD U5194 (.O(n3769), 
	.B2(n457), 
	.B1(\ram[199][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n319));
   AO22CHD U5195 (.O(n3770), 
	.B2(n457), 
	.B1(\ram[199][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n319));
   AO22CHD U5196 (.O(n3771), 
	.B2(n457), 
	.B1(FE_PHN2195_ram_199__5_), 
	.A2(FE_OFN56_n13), 
	.A1(n319));
   AO22CHD U5197 (.O(n3772), 
	.B2(n457), 
	.B1(\ram[199][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n319));
   AO22CHD U5198 (.O(n3773), 
	.B2(n457), 
	.B1(\ram[199][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n319));
   AO22CHD U5199 (.O(n3774), 
	.B2(n457), 
	.B1(\ram[199][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n319));
   AO22CHD U5200 (.O(n3775), 
	.B2(n457), 
	.B1(\ram[199][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n319));
   AO22CHD U5201 (.O(n3776), 
	.B2(n457), 
	.B1(\ram[199][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n319));
   AO22CHD U5202 (.O(n3777), 
	.B2(n457), 
	.B1(\ram[199][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n319));
   AO22CHD U5203 (.O(n3778), 
	.B2(n457), 
	.B1(\ram[199][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n319));
   AO22CHD U5204 (.O(n3779), 
	.B2(n457), 
	.B1(\ram[199][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n319));
   AO22CHD U5205 (.O(n3780), 
	.B2(n457), 
	.B1(\ram[199][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n319));
   AO22CHD U5206 (.O(n3781), 
	.B2(n457), 
	.B1(\ram[199][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n319));
   AO22CHD U5207 (.O(n3782), 
	.B2(n459), 
	.B1(\ram[200][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n321));
   AO22CHD U5208 (.O(n3783), 
	.B2(n459), 
	.B1(\ram[200][1] ), 
	.A2(n9), 
	.A1(n321));
   AO22CHD U5209 (.O(n3784), 
	.B2(n459), 
	.B1(\ram[200][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n321));
   AO22CHD U5210 (.O(n3785), 
	.B2(n459), 
	.B1(\ram[200][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n321));
   AO22CHD U5211 (.O(n3786), 
	.B2(n459), 
	.B1(\ram[200][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n321));
   AO22CHD U5212 (.O(n3787), 
	.B2(n459), 
	.B1(\ram[200][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n321));
   AO22CHD U5213 (.O(n3788), 
	.B2(n459), 
	.B1(\ram[200][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n321));
   AO22CHD U5214 (.O(n3789), 
	.B2(n459), 
	.B1(\ram[200][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n321));
   AO22CHD U5215 (.O(n3790), 
	.B2(n459), 
	.B1(\ram[200][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n321));
   AO22CHD U5216 (.O(n3791), 
	.B2(n459), 
	.B1(\ram[200][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n321));
   AO22CHD U5217 (.O(n3792), 
	.B2(n459), 
	.B1(\ram[200][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n321));
   AO22CHD U5218 (.O(n3793), 
	.B2(n459), 
	.B1(\ram[200][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n321));
   AO22CHD U5219 (.O(n3794), 
	.B2(n459), 
	.B1(\ram[200][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n321));
   AO22CHD U5220 (.O(n3795), 
	.B2(n459), 
	.B1(\ram[200][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n321));
   AO22CHD U5221 (.O(n3796), 
	.B2(n459), 
	.B1(\ram[200][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n321));
   AO22CHD U5222 (.O(n3797), 
	.B2(n459), 
	.B1(\ram[200][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n321));
   AO22CHD U5223 (.O(n3798), 
	.B2(n461), 
	.B1(\ram[201][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n323));
   AO22CHD U5224 (.O(n3799), 
	.B2(n461), 
	.B1(\ram[201][1] ), 
	.A2(n9), 
	.A1(n323));
   AO22CHD U5225 (.O(n3800), 
	.B2(n461), 
	.B1(\ram[201][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n323));
   AO22CHD U5226 (.O(n3801), 
	.B2(n461), 
	.B1(\ram[201][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n323));
   AO22CHD U5227 (.O(n3802), 
	.B2(n461), 
	.B1(\ram[201][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n323));
   AO22CHD U5228 (.O(n3803), 
	.B2(n461), 
	.B1(FE_PHN1058_ram_201__5_), 
	.A2(FE_OFN56_n13), 
	.A1(n323));
   AO22CHD U5229 (.O(n3804), 
	.B2(n461), 
	.B1(\ram[201][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n323));
   AO22CHD U5230 (.O(n3805), 
	.B2(n461), 
	.B1(\ram[201][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n323));
   AO22CHD U5231 (.O(n3806), 
	.B2(n461), 
	.B1(\ram[201][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n323));
   AO22CHD U5232 (.O(n3807), 
	.B2(n461), 
	.B1(\ram[201][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n323));
   AO22CHD U5233 (.O(n3808), 
	.B2(n461), 
	.B1(\ram[201][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n323));
   AO22CHD U5234 (.O(n3809), 
	.B2(n461), 
	.B1(\ram[201][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n323));
   AO22CHD U5235 (.O(n3810), 
	.B2(n461), 
	.B1(\ram[201][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n323));
   AO22CHD U5236 (.O(n3811), 
	.B2(n461), 
	.B1(\ram[201][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n323));
   AO22CHD U5237 (.O(n3812), 
	.B2(n461), 
	.B1(\ram[201][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n323));
   AO22CHD U5238 (.O(n3813), 
	.B2(n461), 
	.B1(\ram[201][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n323));
   AO22CHD U5239 (.O(n3814), 
	.B2(n463), 
	.B1(\ram[202][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n325));
   AO22CHD U5240 (.O(n3815), 
	.B2(n463), 
	.B1(\ram[202][1] ), 
	.A2(n9), 
	.A1(n325));
   AO22CHD U5241 (.O(n3816), 
	.B2(n463), 
	.B1(\ram[202][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n325));
   AO22CHD U5242 (.O(n3817), 
	.B2(n463), 
	.B1(\ram[202][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n325));
   AO22CHD U5243 (.O(n3818), 
	.B2(n463), 
	.B1(\ram[202][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n325));
   AO22CHD U5244 (.O(n3819), 
	.B2(n463), 
	.B1(\ram[202][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n325));
   AO22CHD U5245 (.O(n3820), 
	.B2(n463), 
	.B1(\ram[202][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n325));
   AO22CHD U5246 (.O(n3821), 
	.B2(n463), 
	.B1(\ram[202][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n325));
   AO22CHD U5247 (.O(n3822), 
	.B2(n463), 
	.B1(\ram[202][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n325));
   AO22CHD U5248 (.O(n3823), 
	.B2(n463), 
	.B1(\ram[202][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n325));
   AO22CHD U5249 (.O(n3824), 
	.B2(n463), 
	.B1(\ram[202][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n325));
   AO22CHD U5250 (.O(n3825), 
	.B2(n463), 
	.B1(\ram[202][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n325));
   AO22CHD U5251 (.O(n3826), 
	.B2(n463), 
	.B1(\ram[202][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n325));
   AO22CHD U5252 (.O(n3827), 
	.B2(n463), 
	.B1(FE_PHN2005_ram_202__13_), 
	.A2(FE_OFN83_n21), 
	.A1(n325));
   AO22CHD U5253 (.O(n3828), 
	.B2(n463), 
	.B1(\ram[202][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n325));
   AO22CHD U5254 (.O(n3829), 
	.B2(n463), 
	.B1(\ram[202][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n325));
   AO22CHD U5255 (.O(n3830), 
	.B2(n465), 
	.B1(\ram[203][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n327));
   AO22CHD U5256 (.O(n3831), 
	.B2(n465), 
	.B1(\ram[203][1] ), 
	.A2(n9), 
	.A1(n327));
   AO22CHD U5257 (.O(n3832), 
	.B2(n465), 
	.B1(\ram[203][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n327));
   AO22CHD U5258 (.O(n3833), 
	.B2(n465), 
	.B1(\ram[203][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n327));
   AO22CHD U5259 (.O(n3834), 
	.B2(n465), 
	.B1(\ram[203][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n327));
   AO22CHD U5260 (.O(n3835), 
	.B2(n465), 
	.B1(\ram[203][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n327));
   AO22CHD U5261 (.O(n3836), 
	.B2(n465), 
	.B1(\ram[203][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n327));
   AO22CHD U5262 (.O(n3837), 
	.B2(n465), 
	.B1(\ram[203][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n327));
   AO22CHD U5263 (.O(n3838), 
	.B2(n465), 
	.B1(\ram[203][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n327));
   AO22CHD U5264 (.O(n3839), 
	.B2(n465), 
	.B1(\ram[203][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n327));
   AO22CHD U5265 (.O(n3840), 
	.B2(n465), 
	.B1(\ram[203][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n327));
   AO22CHD U5266 (.O(n3841), 
	.B2(n465), 
	.B1(\ram[203][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n327));
   AO22CHD U5267 (.O(n3842), 
	.B2(n465), 
	.B1(\ram[203][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n327));
   AO22CHD U5268 (.O(n3843), 
	.B2(n465), 
	.B1(\ram[203][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n327));
   AO22CHD U5269 (.O(n3844), 
	.B2(n465), 
	.B1(\ram[203][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n327));
   AO22CHD U5270 (.O(n3845), 
	.B2(n465), 
	.B1(\ram[203][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n327));
   AO22CHD U5271 (.O(n3846), 
	.B2(n467), 
	.B1(\ram[204][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n329));
   AO22CHD U5272 (.O(n3847), 
	.B2(n467), 
	.B1(\ram[204][1] ), 
	.A2(n9), 
	.A1(n329));
   AO22CHD U5273 (.O(n3848), 
	.B2(n467), 
	.B1(\ram[204][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n329));
   AO22CHD U5274 (.O(n3849), 
	.B2(n467), 
	.B1(\ram[204][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n329));
   AO22CHD U5275 (.O(n3850), 
	.B2(n467), 
	.B1(\ram[204][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n329));
   AO22CHD U5276 (.O(n3851), 
	.B2(n467), 
	.B1(\ram[204][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n329));
   AO22CHD U5277 (.O(n3852), 
	.B2(n467), 
	.B1(\ram[204][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n329));
   AO22CHD U5278 (.O(n3853), 
	.B2(n467), 
	.B1(\ram[204][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n329));
   AO22CHD U5279 (.O(n3854), 
	.B2(n467), 
	.B1(\ram[204][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n329));
   AO22CHD U5280 (.O(n3855), 
	.B2(n467), 
	.B1(\ram[204][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n329));
   AO22CHD U5281 (.O(n3856), 
	.B2(n467), 
	.B1(\ram[204][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n329));
   AO22CHD U5282 (.O(n3857), 
	.B2(n467), 
	.B1(\ram[204][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n329));
   AO22CHD U5283 (.O(n3858), 
	.B2(n467), 
	.B1(\ram[204][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n329));
   AO22CHD U5284 (.O(n3859), 
	.B2(n467), 
	.B1(\ram[204][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n329));
   AO22CHD U5285 (.O(n3860), 
	.B2(n467), 
	.B1(\ram[204][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n329));
   AO22CHD U5286 (.O(n3861), 
	.B2(n467), 
	.B1(\ram[204][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n329));
   AO22CHD U5287 (.O(n3862), 
	.B2(n469), 
	.B1(\ram[205][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n331));
   AO22CHD U5288 (.O(n3863), 
	.B2(n469), 
	.B1(\ram[205][1] ), 
	.A2(n9), 
	.A1(n331));
   AO22CHD U5289 (.O(n3864), 
	.B2(n469), 
	.B1(\ram[205][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n331));
   AO22CHD U5290 (.O(n3865), 
	.B2(n469), 
	.B1(\ram[205][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n331));
   AO22CHD U5291 (.O(n3866), 
	.B2(n469), 
	.B1(\ram[205][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n331));
   AO22CHD U5292 (.O(n3867), 
	.B2(n469), 
	.B1(\ram[205][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n331));
   AO22CHD U5293 (.O(n3868), 
	.B2(n469), 
	.B1(\ram[205][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n331));
   AO22CHD U5294 (.O(n3869), 
	.B2(n469), 
	.B1(\ram[205][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n331));
   AO22CHD U5295 (.O(n3870), 
	.B2(n469), 
	.B1(\ram[205][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n331));
   AO22CHD U5296 (.O(n3871), 
	.B2(n469), 
	.B1(\ram[205][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n331));
   AO22CHD U5297 (.O(n3872), 
	.B2(n469), 
	.B1(\ram[205][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n331));
   AO22CHD U5298 (.O(n3873), 
	.B2(n469), 
	.B1(\ram[205][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n331));
   AO22CHD U5299 (.O(n3874), 
	.B2(n469), 
	.B1(\ram[205][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n331));
   AO22CHD U5300 (.O(n3875), 
	.B2(n469), 
	.B1(\ram[205][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n331));
   AO22CHD U5301 (.O(n3876), 
	.B2(n469), 
	.B1(\ram[205][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n331));
   AO22CHD U5302 (.O(n3877), 
	.B2(n469), 
	.B1(\ram[205][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n331));
   AO22CHD U5303 (.O(n3878), 
	.B2(n471), 
	.B1(\ram[206][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n333));
   AO22CHD U5304 (.O(n3879), 
	.B2(n471), 
	.B1(\ram[206][1] ), 
	.A2(n9), 
	.A1(n333));
   AO22CHD U5305 (.O(n3880), 
	.B2(n471), 
	.B1(\ram[206][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n333));
   AO22CHD U5306 (.O(n3881), 
	.B2(n471), 
	.B1(\ram[206][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n333));
   AO22CHD U5307 (.O(n3882), 
	.B2(n471), 
	.B1(\ram[206][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n333));
   AO22CHD U5308 (.O(n3883), 
	.B2(n471), 
	.B1(\ram[206][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n333));
   AO22CHD U5309 (.O(n3884), 
	.B2(n471), 
	.B1(\ram[206][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n333));
   AO22CHD U5310 (.O(n3885), 
	.B2(n471), 
	.B1(\ram[206][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n333));
   AO22CHD U5311 (.O(n3886), 
	.B2(n471), 
	.B1(\ram[206][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n333));
   AO22CHD U5312 (.O(n3887), 
	.B2(n471), 
	.B1(\ram[206][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n333));
   AO22CHD U5313 (.O(n3888), 
	.B2(n471), 
	.B1(\ram[206][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n333));
   AO22CHD U5314 (.O(n3889), 
	.B2(n471), 
	.B1(\ram[206][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n333));
   AO22CHD U5315 (.O(n3890), 
	.B2(n471), 
	.B1(\ram[206][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n333));
   AO22CHD U5316 (.O(n3891), 
	.B2(n471), 
	.B1(\ram[206][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n333));
   AO22CHD U5317 (.O(n3892), 
	.B2(n471), 
	.B1(\ram[206][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n333));
   AO22CHD U5318 (.O(n3893), 
	.B2(n471), 
	.B1(\ram[206][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n333));
   AO22CHD U5319 (.O(n3894), 
	.B2(n473), 
	.B1(\ram[207][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n335));
   AO22CHD U5320 (.O(n3895), 
	.B2(n473), 
	.B1(\ram[207][1] ), 
	.A2(n9), 
	.A1(n335));
   AO22CHD U5321 (.O(n3896), 
	.B2(n473), 
	.B1(\ram[207][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n335));
   AO22CHD U5322 (.O(n3897), 
	.B2(n473), 
	.B1(\ram[207][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n335));
   AO22CHD U5323 (.O(n3898), 
	.B2(n473), 
	.B1(\ram[207][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n335));
   AO22CHD U5324 (.O(n3899), 
	.B2(n473), 
	.B1(\ram[207][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n335));
   AO22CHD U5325 (.O(n3900), 
	.B2(n473), 
	.B1(\ram[207][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n335));
   AO22CHD U5326 (.O(n3901), 
	.B2(n473), 
	.B1(\ram[207][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n335));
   AO22CHD U5327 (.O(n3902), 
	.B2(n473), 
	.B1(\ram[207][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n335));
   AO22CHD U5328 (.O(n3903), 
	.B2(n473), 
	.B1(\ram[207][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n335));
   AO22CHD U5329 (.O(n3904), 
	.B2(n473), 
	.B1(\ram[207][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n335));
   AO22CHD U5330 (.O(n3905), 
	.B2(n473), 
	.B1(\ram[207][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n335));
   AO22CHD U5331 (.O(n3906), 
	.B2(n473), 
	.B1(\ram[207][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n335));
   AO22CHD U5332 (.O(n3907), 
	.B2(n473), 
	.B1(\ram[207][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n335));
   AO22CHD U5333 (.O(n3908), 
	.B2(n473), 
	.B1(\ram[207][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n335));
   AO22CHD U5334 (.O(n3909), 
	.B2(n473), 
	.B1(\ram[207][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n335));
   AO22CHD U5335 (.O(n3910), 
	.B2(n476), 
	.B1(\ram[208][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n337));
   AO22CHD U5336 (.O(n3911), 
	.B2(n476), 
	.B1(\ram[208][1] ), 
	.A2(n9), 
	.A1(n337));
   AO22CHD U5337 (.O(n3912), 
	.B2(n476), 
	.B1(\ram[208][2] ), 
	.A2(n10), 
	.A1(n337));
   AO22CHD U5338 (.O(n3913), 
	.B2(n476), 
	.B1(\ram[208][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n337));
   AO22CHD U5339 (.O(n3914), 
	.B2(n476), 
	.B1(\ram[208][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n337));
   AO22CHD U5340 (.O(n3915), 
	.B2(n476), 
	.B1(\ram[208][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n337));
   AO22CHD U5341 (.O(n3916), 
	.B2(n476), 
	.B1(\ram[208][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n337));
   AO22CHD U5342 (.O(n3917), 
	.B2(n476), 
	.B1(\ram[208][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n337));
   AO22CHD U5343 (.O(n3918), 
	.B2(n476), 
	.B1(\ram[208][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n337));
   AO22CHD U5344 (.O(n3919), 
	.B2(n476), 
	.B1(\ram[208][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n337));
   AO22CHD U5345 (.O(n3920), 
	.B2(n476), 
	.B1(\ram[208][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n337));
   AO22CHD U5346 (.O(n3921), 
	.B2(n476), 
	.B1(\ram[208][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n337));
   AO22CHD U5347 (.O(n3922), 
	.B2(n476), 
	.B1(\ram[208][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n337));
   AO22CHD U5348 (.O(n3923), 
	.B2(n476), 
	.B1(\ram[208][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n337));
   AO22CHD U5349 (.O(n3924), 
	.B2(n476), 
	.B1(\ram[208][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n337));
   AO22CHD U5350 (.O(n3925), 
	.B2(n476), 
	.B1(\ram[208][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n337));
   AO22CHD U5351 (.O(n3926), 
	.B2(n479), 
	.B1(\ram[209][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n339));
   AO22CHD U5352 (.O(n3927), 
	.B2(n479), 
	.B1(\ram[209][1] ), 
	.A2(n9), 
	.A1(n339));
   AO22CHD U5353 (.O(n3928), 
	.B2(n479), 
	.B1(\ram[209][2] ), 
	.A2(n10), 
	.A1(n339));
   AO22CHD U5354 (.O(n3929), 
	.B2(n479), 
	.B1(\ram[209][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n339));
   AO22CHD U5355 (.O(n3930), 
	.B2(n479), 
	.B1(\ram[209][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n339));
   AO22CHD U5356 (.O(n3931), 
	.B2(n479), 
	.B1(\ram[209][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n339));
   AO22CHD U5357 (.O(n3932), 
	.B2(n479), 
	.B1(\ram[209][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n339));
   AO22CHD U5358 (.O(n3933), 
	.B2(n479), 
	.B1(\ram[209][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n339));
   AO22CHD U5359 (.O(n3934), 
	.B2(n479), 
	.B1(\ram[209][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n339));
   AO22CHD U5360 (.O(n3935), 
	.B2(n479), 
	.B1(\ram[209][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n339));
   AO22CHD U5361 (.O(n3936), 
	.B2(n479), 
	.B1(\ram[209][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n339));
   AO22CHD U5362 (.O(n3937), 
	.B2(n479), 
	.B1(\ram[209][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n339));
   AO22CHD U5363 (.O(n3938), 
	.B2(n479), 
	.B1(\ram[209][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n339));
   AO22CHD U5364 (.O(n3939), 
	.B2(n479), 
	.B1(\ram[209][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n339));
   AO22CHD U5365 (.O(n3940), 
	.B2(n479), 
	.B1(\ram[209][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n339));
   AO22CHD U5366 (.O(n3941), 
	.B2(n479), 
	.B1(\ram[209][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n339));
   AO22CHD U5367 (.O(n3942), 
	.B2(n481), 
	.B1(\ram[210][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n342));
   AO22CHD U5368 (.O(n3943), 
	.B2(n481), 
	.B1(\ram[210][1] ), 
	.A2(n9), 
	.A1(n342));
   AO22CHD U5369 (.O(n3944), 
	.B2(n481), 
	.B1(\ram[210][2] ), 
	.A2(n10), 
	.A1(n342));
   AO22CHD U5370 (.O(n3945), 
	.B2(n481), 
	.B1(\ram[210][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n342));
   AO22CHD U5371 (.O(n3946), 
	.B2(n481), 
	.B1(\ram[210][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n342));
   AO22CHD U5372 (.O(n3947), 
	.B2(n481), 
	.B1(\ram[210][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n342));
   AO22CHD U5373 (.O(n3948), 
	.B2(n481), 
	.B1(\ram[210][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n342));
   AO22CHD U5374 (.O(n3949), 
	.B2(n481), 
	.B1(\ram[210][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n342));
   AO22CHD U5375 (.O(n3950), 
	.B2(n481), 
	.B1(\ram[210][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n342));
   AO22CHD U5376 (.O(n3951), 
	.B2(n481), 
	.B1(\ram[210][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n342));
   AO22CHD U5377 (.O(n3952), 
	.B2(n481), 
	.B1(\ram[210][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n342));
   AO22CHD U5378 (.O(n3953), 
	.B2(n481), 
	.B1(\ram[210][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n342));
   AO22CHD U5379 (.O(n3954), 
	.B2(n481), 
	.B1(\ram[210][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n342));
   AO22CHD U5380 (.O(n3955), 
	.B2(n481), 
	.B1(\ram[210][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n342));
   AO22CHD U5381 (.O(n3956), 
	.B2(n481), 
	.B1(\ram[210][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n342));
   AO22CHD U5382 (.O(n3957), 
	.B2(n481), 
	.B1(\ram[210][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n342));
   AO22CHD U5383 (.O(n3958), 
	.B2(n483), 
	.B1(\ram[211][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n344));
   AO22CHD U5384 (.O(n3959), 
	.B2(n483), 
	.B1(\ram[211][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n344));
   AO22CHD U5385 (.O(n3960), 
	.B2(n483), 
	.B1(\ram[211][2] ), 
	.A2(n10), 
	.A1(n344));
   AO22CHD U5386 (.O(n3961), 
	.B2(n483), 
	.B1(\ram[211][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n344));
   AO22CHD U5387 (.O(n3962), 
	.B2(n483), 
	.B1(\ram[211][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n344));
   AO22CHD U5388 (.O(n3963), 
	.B2(n483), 
	.B1(\ram[211][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n344));
   AO22CHD U5389 (.O(FE_PHN7453_n3964), 
	.B2(n483), 
	.B1(\ram[211][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n344));
   AO22CHD U5390 (.O(n3965), 
	.B2(n483), 
	.B1(\ram[211][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n344));
   AO22CHD U5391 (.O(n3966), 
	.B2(n483), 
	.B1(\ram[211][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n344));
   AO22CHD U5392 (.O(n3967), 
	.B2(n483), 
	.B1(\ram[211][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n344));
   AO22CHD U5393 (.O(n3968), 
	.B2(n483), 
	.B1(\ram[211][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n344));
   AO22CHD U5394 (.O(n3969), 
	.B2(n483), 
	.B1(\ram[211][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n344));
   AO22CHD U5395 (.O(n3970), 
	.B2(n483), 
	.B1(\ram[211][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n344));
   AO22CHD U5396 (.O(n3971), 
	.B2(n483), 
	.B1(\ram[211][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n344));
   AO22CHD U5397 (.O(n3972), 
	.B2(n483), 
	.B1(\ram[211][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n344));
   AO22CHD U5398 (.O(n3973), 
	.B2(n483), 
	.B1(\ram[211][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n344));
   AO22CHD U5399 (.O(n3974), 
	.B2(n485), 
	.B1(\ram[212][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n345));
   AO22CHD U5400 (.O(n3975), 
	.B2(n485), 
	.B1(\ram[212][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n345));
   AO22CHD U5401 (.O(n3976), 
	.B2(n485), 
	.B1(\ram[212][2] ), 
	.A2(n10), 
	.A1(n345));
   AO22CHD U5402 (.O(n3977), 
	.B2(n485), 
	.B1(\ram[212][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n345));
   AO22CHD U5403 (.O(n3978), 
	.B2(n485), 
	.B1(\ram[212][4] ), 
	.A2(n12), 
	.A1(n345));
   AO22CHD U5404 (.O(n3979), 
	.B2(n485), 
	.B1(\ram[212][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n345));
   AO22CHD U5405 (.O(n3980), 
	.B2(n485), 
	.B1(\ram[212][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n345));
   AO22CHD U5406 (.O(n3981), 
	.B2(n485), 
	.B1(\ram[212][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n345));
   AO22CHD U5407 (.O(n3982), 
	.B2(n485), 
	.B1(\ram[212][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n345));
   AO22CHD U5408 (.O(n3983), 
	.B2(n485), 
	.B1(\ram[212][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n345));
   AO22CHD U5409 (.O(n3984), 
	.B2(n485), 
	.B1(\ram[212][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n345));
   AO22CHD U5410 (.O(n3985), 
	.B2(n485), 
	.B1(\ram[212][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n345));
   AO22CHD U5411 (.O(n3986), 
	.B2(n485), 
	.B1(\ram[212][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n345));
   AO22CHD U5412 (.O(n3987), 
	.B2(n485), 
	.B1(\ram[212][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n345));
   AO22CHD U5413 (.O(n3988), 
	.B2(n485), 
	.B1(\ram[212][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n345));
   AO22CHD U5414 (.O(n3989), 
	.B2(n485), 
	.B1(\ram[212][15] ), 
	.A2(n23), 
	.A1(n345));
   AO22CHD U5415 (.O(n3990), 
	.B2(n487), 
	.B1(\ram[213][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n347));
   AO22CHD U5416 (.O(n3991), 
	.B2(n487), 
	.B1(\ram[213][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n347));
   AO22CHD U5417 (.O(n3992), 
	.B2(n487), 
	.B1(\ram[213][2] ), 
	.A2(n10), 
	.A1(n347));
   AO22CHD U5418 (.O(n3993), 
	.B2(n487), 
	.B1(\ram[213][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n347));
   AO22CHD U5419 (.O(n3994), 
	.B2(n487), 
	.B1(\ram[213][4] ), 
	.A2(n12), 
	.A1(n347));
   AO22CHD U5420 (.O(n3995), 
	.B2(n487), 
	.B1(\ram[213][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n347));
   AO22CHD U5421 (.O(n3996), 
	.B2(n487), 
	.B1(\ram[213][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n347));
   AO22CHD U5422 (.O(n3997), 
	.B2(n487), 
	.B1(\ram[213][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n347));
   AO22CHD U5423 (.O(n3998), 
	.B2(n487), 
	.B1(\ram[213][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n347));
   AO22CHD U5424 (.O(n3999), 
	.B2(n487), 
	.B1(\ram[213][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n347));
   AO22CHD U5425 (.O(n4000), 
	.B2(n487), 
	.B1(\ram[213][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n347));
   AO22CHD U5426 (.O(n4001), 
	.B2(n487), 
	.B1(\ram[213][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n347));
   AO22CHD U5427 (.O(n4002), 
	.B2(n487), 
	.B1(\ram[213][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n347));
   AO22CHD U5428 (.O(n4003), 
	.B2(n487), 
	.B1(\ram[213][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n347));
   AO22CHD U5429 (.O(n4004), 
	.B2(n487), 
	.B1(\ram[213][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n347));
   AO22CHD U5430 (.O(n4005), 
	.B2(n487), 
	.B1(\ram[213][15] ), 
	.A2(n23), 
	.A1(n347));
   AO22CHD U5431 (.O(n4006), 
	.B2(n489), 
	.B1(\ram[214][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n349));
   AO22CHD U5432 (.O(n4007), 
	.B2(n489), 
	.B1(\ram[214][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n349));
   AO22CHD U5433 (.O(n4008), 
	.B2(n489), 
	.B1(\ram[214][2] ), 
	.A2(n10), 
	.A1(n349));
   AO22CHD U5434 (.O(n4009), 
	.B2(n489), 
	.B1(\ram[214][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n349));
   AO22CHD U5435 (.O(n4010), 
	.B2(n489), 
	.B1(\ram[214][4] ), 
	.A2(n12), 
	.A1(n349));
   AO22CHD U5436 (.O(n4011), 
	.B2(n489), 
	.B1(\ram[214][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n349));
   AO22CHD U5437 (.O(n4012), 
	.B2(n489), 
	.B1(\ram[214][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n349));
   AO22CHD U5438 (.O(n4013), 
	.B2(n489), 
	.B1(\ram[214][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n349));
   AO22CHD U5439 (.O(n4014), 
	.B2(n489), 
	.B1(\ram[214][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n349));
   AO22CHD U5440 (.O(n4015), 
	.B2(n489), 
	.B1(\ram[214][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n349));
   AO22CHD U5441 (.O(n4016), 
	.B2(n489), 
	.B1(\ram[214][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n349));
   AO22CHD U5442 (.O(n4017), 
	.B2(n489), 
	.B1(\ram[214][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n349));
   AO22CHD U5443 (.O(n4018), 
	.B2(n489), 
	.B1(\ram[214][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n349));
   AO22CHD U5444 (.O(n4019), 
	.B2(n489), 
	.B1(FE_PHN5476_ram_214__13_), 
	.A2(FE_OFN83_n21), 
	.A1(n349));
   AO22CHD U5445 (.O(n4020), 
	.B2(n489), 
	.B1(\ram[214][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n349));
   AO22CHD U5446 (.O(n4021), 
	.B2(n489), 
	.B1(\ram[214][15] ), 
	.A2(n23), 
	.A1(n349));
   AO22CHD U5447 (.O(n4022), 
	.B2(n491), 
	.B1(\ram[215][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n351));
   AO22CHD U5448 (.O(n4023), 
	.B2(n491), 
	.B1(\ram[215][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n351));
   AO22CHD U5449 (.O(n4024), 
	.B2(n491), 
	.B1(\ram[215][2] ), 
	.A2(n10), 
	.A1(n351));
   AO22CHD U5450 (.O(n4025), 
	.B2(n491), 
	.B1(\ram[215][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n351));
   AO22CHD U5451 (.O(n4026), 
	.B2(n491), 
	.B1(\ram[215][4] ), 
	.A2(n12), 
	.A1(n351));
   AO22CHD U5452 (.O(n4027), 
	.B2(n491), 
	.B1(\ram[215][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n351));
   AO22CHD U5453 (.O(n4028), 
	.B2(n491), 
	.B1(\ram[215][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n351));
   AO22CHD U5454 (.O(n4029), 
	.B2(n491), 
	.B1(\ram[215][7] ), 
	.A2(FE_OFN64_n15), 
	.A1(n351));
   AO22CHD U5455 (.O(n4030), 
	.B2(n491), 
	.B1(\ram[215][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n351));
   AO22CHD U5456 (.O(n4031), 
	.B2(n491), 
	.B1(\ram[215][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n351));
   AO22CHD U5457 (.O(n4032), 
	.B2(n491), 
	.B1(\ram[215][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n351));
   AO22CHD U5458 (.O(n4033), 
	.B2(n491), 
	.B1(\ram[215][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n351));
   AO22CHD U5459 (.O(n4034), 
	.B2(n491), 
	.B1(\ram[215][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n351));
   AO22CHD U5460 (.O(n4035), 
	.B2(n491), 
	.B1(\ram[215][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n351));
   AO22CHD U5461 (.O(n4036), 
	.B2(n491), 
	.B1(\ram[215][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n351));
   AO22CHD U5462 (.O(n4037), 
	.B2(n491), 
	.B1(\ram[215][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n351));
   AO22CHD U5463 (.O(n4038), 
	.B2(n493), 
	.B1(\ram[216][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n353));
   AO22CHD U5464 (.O(n4039), 
	.B2(n493), 
	.B1(\ram[216][1] ), 
	.A2(n9), 
	.A1(n353));
   AO22CHD U5465 (.O(n4040), 
	.B2(n493), 
	.B1(\ram[216][2] ), 
	.A2(n10), 
	.A1(n353));
   AO22CHD U5466 (.O(n4041), 
	.B2(n493), 
	.B1(\ram[216][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n353));
   AO22CHD U5467 (.O(n4042), 
	.B2(n493), 
	.B1(\ram[216][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n353));
   AO22CHD U5468 (.O(n4043), 
	.B2(n493), 
	.B1(\ram[216][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n353));
   AO22CHD U5469 (.O(n4044), 
	.B2(n493), 
	.B1(\ram[216][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n353));
   AO22CHD U5470 (.O(n4045), 
	.B2(n493), 
	.B1(\ram[216][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n353));
   AO22CHD U5471 (.O(n4046), 
	.B2(n493), 
	.B1(\ram[216][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n353));
   AO22CHD U5472 (.O(n4047), 
	.B2(n493), 
	.B1(\ram[216][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n353));
   AO22CHD U5473 (.O(n4048), 
	.B2(n493), 
	.B1(\ram[216][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n353));
   AO22CHD U5474 (.O(n4049), 
	.B2(n493), 
	.B1(\ram[216][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n353));
   AO22CHD U5475 (.O(n4050), 
	.B2(n493), 
	.B1(\ram[216][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n353));
   AO22CHD U5476 (.O(n4051), 
	.B2(n493), 
	.B1(\ram[216][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n353));
   AO22CHD U5477 (.O(n4052), 
	.B2(n493), 
	.B1(\ram[216][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n353));
   AO22CHD U5478 (.O(n4053), 
	.B2(n493), 
	.B1(\ram[216][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n353));
   AO22CHD U5479 (.O(n4054), 
	.B2(n495), 
	.B1(\ram[217][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n355));
   AO22CHD U5480 (.O(n4055), 
	.B2(n495), 
	.B1(\ram[217][1] ), 
	.A2(n9), 
	.A1(n355));
   AO22CHD U5481 (.O(n4056), 
	.B2(n495), 
	.B1(\ram[217][2] ), 
	.A2(n10), 
	.A1(n355));
   AO22CHD U5482 (.O(n4057), 
	.B2(n495), 
	.B1(FE_PHN2286_ram_217__3_), 
	.A2(FE_OFN50_n11), 
	.A1(n355));
   AO22CHD U5483 (.O(n4058), 
	.B2(n495), 
	.B1(\ram[217][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n355));
   AO22CHD U5484 (.O(n4059), 
	.B2(n495), 
	.B1(\ram[217][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n355));
   AO22CHD U5485 (.O(n4060), 
	.B2(n495), 
	.B1(\ram[217][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n355));
   AO22CHD U5486 (.O(n4061), 
	.B2(n495), 
	.B1(\ram[217][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n355));
   AO22CHD U5487 (.O(n4062), 
	.B2(n495), 
	.B1(\ram[217][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n355));
   AO22CHD U5488 (.O(n4063), 
	.B2(n495), 
	.B1(\ram[217][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n355));
   AO22CHD U5489 (.O(n4064), 
	.B2(n495), 
	.B1(\ram[217][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n355));
   AO22CHD U5490 (.O(n4065), 
	.B2(n495), 
	.B1(\ram[217][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n355));
   AO22CHD U5491 (.O(n4066), 
	.B2(n495), 
	.B1(\ram[217][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n355));
   AO22CHD U5492 (.O(n4067), 
	.B2(n495), 
	.B1(\ram[217][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n355));
   AO22CHD U5493 (.O(n4068), 
	.B2(n495), 
	.B1(\ram[217][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n355));
   AO22CHD U5494 (.O(n4069), 
	.B2(n495), 
	.B1(\ram[217][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n355));
   AO22CHD U5495 (.O(n4070), 
	.B2(n497), 
	.B1(\ram[218][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n357));
   AO22CHD U5496 (.O(n4071), 
	.B2(n497), 
	.B1(\ram[218][1] ), 
	.A2(n9), 
	.A1(n357));
   AO22CHD U5497 (.O(n4072), 
	.B2(n497), 
	.B1(\ram[218][2] ), 
	.A2(n10), 
	.A1(n357));
   AO22CHD U5498 (.O(n4073), 
	.B2(n497), 
	.B1(\ram[218][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n357));
   AO22CHD U5499 (.O(n4074), 
	.B2(n497), 
	.B1(\ram[218][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n357));
   AO22CHD U5500 (.O(n4075), 
	.B2(n497), 
	.B1(\ram[218][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n357));
   AO22CHD U5501 (.O(n4076), 
	.B2(n497), 
	.B1(\ram[218][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n357));
   AO22CHD U5502 (.O(n4077), 
	.B2(n497), 
	.B1(\ram[218][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n357));
   AO22CHD U5503 (.O(n4078), 
	.B2(n497), 
	.B1(\ram[218][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n357));
   AO22CHD U5504 (.O(n4079), 
	.B2(n497), 
	.B1(\ram[218][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n357));
   AO22CHD U5505 (.O(n4080), 
	.B2(n497), 
	.B1(\ram[218][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n357));
   AO22CHD U5506 (.O(n4081), 
	.B2(n497), 
	.B1(\ram[218][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n357));
   AO22CHD U5507 (.O(n4082), 
	.B2(n497), 
	.B1(\ram[218][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n357));
   AO22CHD U5508 (.O(n4083), 
	.B2(n497), 
	.B1(\ram[218][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n357));
   AO22CHD U5509 (.O(n4084), 
	.B2(n497), 
	.B1(\ram[218][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n357));
   AO22CHD U5510 (.O(n4085), 
	.B2(n497), 
	.B1(\ram[218][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n357));
   AO22CHD U5511 (.O(n4086), 
	.B2(n499), 
	.B1(\ram[219][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n359));
   AO22CHD U5512 (.O(n4087), 
	.B2(n499), 
	.B1(\ram[219][1] ), 
	.A2(n9), 
	.A1(n359));
   AO22CHD U5513 (.O(n4088), 
	.B2(n499), 
	.B1(\ram[219][2] ), 
	.A2(n10), 
	.A1(n359));
   AO22CHD U5514 (.O(n4089), 
	.B2(n499), 
	.B1(\ram[219][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n359));
   AO22CHD U5515 (.O(n4090), 
	.B2(n499), 
	.B1(\ram[219][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n359));
   AO22CHD U5516 (.O(n4091), 
	.B2(n499), 
	.B1(\ram[219][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n359));
   AO22CHD U5517 (.O(n4092), 
	.B2(n499), 
	.B1(\ram[219][6] ), 
	.A2(FE_OFN60_n14), 
	.A1(n359));
   AO22CHD U5518 (.O(n4093), 
	.B2(n499), 
	.B1(\ram[219][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n359));
   AO22CHD U5519 (.O(n4094), 
	.B2(n499), 
	.B1(\ram[219][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n359));
   AO22CHD U5520 (.O(n4095), 
	.B2(n499), 
	.B1(\ram[219][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n359));
   AO22CHD U5521 (.O(n4096), 
	.B2(n499), 
	.B1(\ram[219][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n359));
   AO22CHD U5522 (.O(n4097), 
	.B2(n499), 
	.B1(\ram[219][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n359));
   AO22CHD U5523 (.O(n4098), 
	.B2(n499), 
	.B1(\ram[219][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n359));
   AO22CHD U5524 (.O(n4099), 
	.B2(n499), 
	.B1(\ram[219][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n359));
   AO22CHD U5525 (.O(n4100), 
	.B2(n499), 
	.B1(\ram[219][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n359));
   AO22CHD U5526 (.O(n4101), 
	.B2(n499), 
	.B1(\ram[219][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n359));
   AO22CHD U5527 (.O(n4102), 
	.B2(n501), 
	.B1(\ram[220][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n361));
   AO22CHD U5528 (.O(n4103), 
	.B2(n501), 
	.B1(\ram[220][1] ), 
	.A2(n9), 
	.A1(n361));
   AO22CHD U5529 (.O(n4104), 
	.B2(n501), 
	.B1(\ram[220][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n361));
   AO22CHD U5530 (.O(n4105), 
	.B2(n501), 
	.B1(\ram[220][3] ), 
	.A2(n11), 
	.A1(n361));
   AO22CHD U5531 (.O(n4106), 
	.B2(n501), 
	.B1(\ram[220][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n361));
   AO22CHD U5532 (.O(n4107), 
	.B2(n501), 
	.B1(\ram[220][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n361));
   AO22CHD U5533 (.O(n4108), 
	.B2(n501), 
	.B1(\ram[220][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n361));
   AO22CHD U5534 (.O(n4109), 
	.B2(n501), 
	.B1(\ram[220][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n361));
   AO22CHD U5535 (.O(n4110), 
	.B2(n501), 
	.B1(\ram[220][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n361));
   AO22CHD U5536 (.O(n4111), 
	.B2(n501), 
	.B1(\ram[220][9] ), 
	.A2(FE_OFN71_n17), 
	.A1(n361));
   AO22CHD U5537 (.O(n4112), 
	.B2(n501), 
	.B1(\ram[220][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n361));
   AO22CHD U5538 (.O(n4113), 
	.B2(n501), 
	.B1(\ram[220][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n361));
   AO22CHD U5539 (.O(n4114), 
	.B2(n501), 
	.B1(\ram[220][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n361));
   AO22CHD U5540 (.O(n4115), 
	.B2(n501), 
	.B1(\ram[220][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n361));
   AO22CHD U5541 (.O(n4116), 
	.B2(n501), 
	.B1(\ram[220][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n361));
   AO22CHD U5542 (.O(n4117), 
	.B2(n501), 
	.B1(\ram[220][15] ), 
	.A2(n23), 
	.A1(n361));
   AO22CHD U5543 (.O(n4118), 
	.B2(n503), 
	.B1(\ram[221][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n363));
   AO22CHD U5544 (.O(n4119), 
	.B2(n503), 
	.B1(FE_PHN5513_ram_221__1_), 
	.A2(n9), 
	.A1(n363));
   AO22CHD U5545 (.O(n4120), 
	.B2(n503), 
	.B1(\ram[221][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n363));
   AO22CHD U5546 (.O(n4121), 
	.B2(n503), 
	.B1(\ram[221][3] ), 
	.A2(n11), 
	.A1(n363));
   AO22CHD U5547 (.O(n4122), 
	.B2(n503), 
	.B1(\ram[221][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n363));
   AO22CHD U5548 (.O(n4123), 
	.B2(n503), 
	.B1(\ram[221][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n363));
   AO22CHD U5549 (.O(n4124), 
	.B2(n503), 
	.B1(\ram[221][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n363));
   AO22CHD U5550 (.O(n4125), 
	.B2(n503), 
	.B1(\ram[221][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n363));
   AO22CHD U5551 (.O(n4126), 
	.B2(n503), 
	.B1(\ram[221][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n363));
   AO22CHD U5552 (.O(n4127), 
	.B2(n503), 
	.B1(\ram[221][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n363));
   AO22CHD U5553 (.O(n4128), 
	.B2(n503), 
	.B1(\ram[221][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n363));
   AO22CHD U5554 (.O(n4129), 
	.B2(n503), 
	.B1(\ram[221][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n363));
   AO22CHD U5555 (.O(n4130), 
	.B2(n503), 
	.B1(\ram[221][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n363));
   AO22CHD U5556 (.O(n4131), 
	.B2(n503), 
	.B1(\ram[221][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n363));
   AO22CHD U5557 (.O(n4132), 
	.B2(n503), 
	.B1(\ram[221][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n363));
   AO22CHD U5558 (.O(n4133), 
	.B2(n503), 
	.B1(\ram[221][15] ), 
	.A2(n23), 
	.A1(n363));
   AO22CHD U5559 (.O(n4134), 
	.B2(n505), 
	.B1(\ram[222][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n365));
   AO22CHD U5560 (.O(n4135), 
	.B2(n505), 
	.B1(\ram[222][1] ), 
	.A2(n9), 
	.A1(n365));
   AO22CHD U5561 (.O(n4136), 
	.B2(n505), 
	.B1(\ram[222][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n365));
   AO22CHD U5562 (.O(n4137), 
	.B2(n505), 
	.B1(\ram[222][3] ), 
	.A2(n11), 
	.A1(n365));
   AO22CHD U5563 (.O(n4138), 
	.B2(n505), 
	.B1(\ram[222][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n365));
   AO22CHD U5564 (.O(n4139), 
	.B2(n505), 
	.B1(\ram[222][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n365));
   AO22CHD U5565 (.O(n4140), 
	.B2(n505), 
	.B1(\ram[222][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n365));
   AO22CHD U5566 (.O(n4141), 
	.B2(n505), 
	.B1(\ram[222][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n365));
   AO22CHD U5567 (.O(n4142), 
	.B2(n505), 
	.B1(\ram[222][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n365));
   AO22CHD U5568 (.O(n4143), 
	.B2(n505), 
	.B1(\ram[222][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n365));
   AO22CHD U5569 (.O(n4144), 
	.B2(n505), 
	.B1(\ram[222][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n365));
   AO22CHD U5570 (.O(n4145), 
	.B2(n505), 
	.B1(\ram[222][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n365));
   AO22CHD U5571 (.O(n4146), 
	.B2(n505), 
	.B1(\ram[222][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n365));
   AO22CHD U5572 (.O(n4147), 
	.B2(n505), 
	.B1(\ram[222][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n365));
   AO22CHD U5573 (.O(n4148), 
	.B2(n505), 
	.B1(\ram[222][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n365));
   AO22CHD U5574 (.O(n4149), 
	.B2(n505), 
	.B1(\ram[222][15] ), 
	.A2(n23), 
	.A1(n365));
   AO22CHD U5575 (.O(n4150), 
	.B2(n507), 
	.B1(\ram[223][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n367));
   AO22CHD U5576 (.O(n4151), 
	.B2(n507), 
	.B1(\ram[223][1] ), 
	.A2(n9), 
	.A1(n367));
   AO22CHD U5577 (.O(n4152), 
	.B2(n507), 
	.B1(\ram[223][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n367));
   AO22CHD U5578 (.O(n4153), 
	.B2(n507), 
	.B1(\ram[223][3] ), 
	.A2(n11), 
	.A1(n367));
   AO22CHD U5579 (.O(n4154), 
	.B2(n507), 
	.B1(\ram[223][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n367));
   AO22CHD U5580 (.O(n4155), 
	.B2(n507), 
	.B1(\ram[223][5] ), 
	.A2(FE_OFN57_n13), 
	.A1(n367));
   AO22CHD U5581 (.O(n4156), 
	.B2(n507), 
	.B1(\ram[223][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n367));
   AO22CHD U5582 (.O(n4157), 
	.B2(n507), 
	.B1(\ram[223][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n367));
   AO22CHD U5583 (.O(n4158), 
	.B2(n507), 
	.B1(\ram[223][8] ), 
	.A2(FE_OFN67_n16), 
	.A1(n367));
   AO22CHD U5584 (.O(n4159), 
	.B2(n507), 
	.B1(\ram[223][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n367));
   AO22CHD U5585 (.O(n4160), 
	.B2(n507), 
	.B1(\ram[223][10] ), 
	.A2(FE_OFN74_n18), 
	.A1(n367));
   AO22CHD U5586 (.O(n4161), 
	.B2(n507), 
	.B1(\ram[223][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n367));
   AO22CHD U5587 (.O(n4162), 
	.B2(n507), 
	.B1(\ram[223][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n367));
   AO22CHD U5588 (.O(n4163), 
	.B2(n507), 
	.B1(\ram[223][13] ), 
	.A2(FE_OFN83_n21), 
	.A1(n367));
   AO22CHD U5589 (.O(n4164), 
	.B2(n507), 
	.B1(\ram[223][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n367));
   AO22CHD U5590 (.O(n4165), 
	.B2(n507), 
	.B1(\ram[223][15] ), 
	.A2(n23), 
	.A1(n367));
   AO22CHD U5591 (.O(n4166), 
	.B2(n509), 
	.B1(\ram[224][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n369));
   AO22CHD U5592 (.O(n4167), 
	.B2(n509), 
	.B1(\ram[224][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n369));
   AO22CHD U5593 (.O(n4168), 
	.B2(n509), 
	.B1(\ram[224][2] ), 
	.A2(n10), 
	.A1(n369));
   AO22CHD U5594 (.O(n4169), 
	.B2(n509), 
	.B1(\ram[224][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n369));
   AO22CHD U5595 (.O(n4170), 
	.B2(n509), 
	.B1(\ram[224][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n369));
   AO22CHD U5596 (.O(n4171), 
	.B2(n509), 
	.B1(\ram[224][5] ), 
	.A2(n13), 
	.A1(n369));
   AO22CHD U5597 (.O(n4172), 
	.B2(n509), 
	.B1(\ram[224][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n369));
   AO22CHD U5598 (.O(n4173), 
	.B2(n509), 
	.B1(\ram[224][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n369));
   AO22CHD U5599 (.O(n4174), 
	.B2(n509), 
	.B1(\ram[224][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n369));
   AO22CHD U5600 (.O(n4175), 
	.B2(n509), 
	.B1(\ram[224][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n369));
   AO22CHD U5601 (.O(n4176), 
	.B2(n509), 
	.B1(\ram[224][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n369));
   AO22CHD U5602 (.O(n4177), 
	.B2(n509), 
	.B1(\ram[224][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n369));
   AO22CHD U5603 (.O(n4178), 
	.B2(n509), 
	.B1(\ram[224][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n369));
   AO22CHD U5604 (.O(n4179), 
	.B2(n509), 
	.B1(\ram[224][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n369));
   AO22CHD U5605 (.O(n4180), 
	.B2(n509), 
	.B1(\ram[224][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n369));
   AO22CHD U5606 (.O(n4181), 
	.B2(n509), 
	.B1(\ram[224][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n369));
   AO22CHD U5607 (.O(n4182), 
	.B2(n512), 
	.B1(\ram[225][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n371));
   AO22CHD U5608 (.O(n4183), 
	.B2(n512), 
	.B1(\ram[225][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n371));
   AO22CHD U5609 (.O(n4184), 
	.B2(n512), 
	.B1(\ram[225][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n371));
   AO22CHD U5610 (.O(n4185), 
	.B2(n512), 
	.B1(\ram[225][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n371));
   AO22CHD U5611 (.O(n4186), 
	.B2(n512), 
	.B1(\ram[225][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n371));
   AO22CHD U5612 (.O(n4187), 
	.B2(n512), 
	.B1(\ram[225][5] ), 
	.A2(n13), 
	.A1(n371));
   AO22CHD U5613 (.O(n4188), 
	.B2(n512), 
	.B1(\ram[225][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n371));
   AO22CHD U5614 (.O(n4189), 
	.B2(n512), 
	.B1(\ram[225][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n371));
   AO22CHD U5615 (.O(n4190), 
	.B2(n512), 
	.B1(\ram[225][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n371));
   AO22CHD U5616 (.O(n4191), 
	.B2(n512), 
	.B1(\ram[225][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n371));
   AO22CHD U5617 (.O(n4192), 
	.B2(n512), 
	.B1(\ram[225][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n371));
   AO22CHD U5618 (.O(n4193), 
	.B2(n512), 
	.B1(\ram[225][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n371));
   AO22CHD U5619 (.O(n4194), 
	.B2(n512), 
	.B1(\ram[225][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n371));
   AO22CHD U5620 (.O(n4195), 
	.B2(n512), 
	.B1(\ram[225][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n371));
   AO22CHD U5621 (.O(n4196), 
	.B2(n512), 
	.B1(\ram[225][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n371));
   AO22CHD U5622 (.O(n4197), 
	.B2(n512), 
	.B1(\ram[225][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n371));
   AO22CHD U5623 (.O(n4198), 
	.B2(n514), 
	.B1(\ram[226][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n373));
   AO22CHD U5624 (.O(n4199), 
	.B2(n514), 
	.B1(\ram[226][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n373));
   AO22CHD U5625 (.O(n4200), 
	.B2(n514), 
	.B1(\ram[226][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n373));
   AO22CHD U5626 (.O(n4201), 
	.B2(n514), 
	.B1(\ram[226][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n373));
   AO22CHD U5627 (.O(n4202), 
	.B2(n514), 
	.B1(\ram[226][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n373));
   AO22CHD U5628 (.O(n4203), 
	.B2(n514), 
	.B1(\ram[226][5] ), 
	.A2(n13), 
	.A1(n373));
   AO22CHD U5629 (.O(n4204), 
	.B2(n514), 
	.B1(\ram[226][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n373));
   AO22CHD U5630 (.O(n4205), 
	.B2(n514), 
	.B1(\ram[226][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n373));
   AO22CHD U5631 (.O(n4206), 
	.B2(n514), 
	.B1(\ram[226][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n373));
   AO22CHD U5632 (.O(n4207), 
	.B2(n514), 
	.B1(\ram[226][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n373));
   AO22CHD U5633 (.O(n4208), 
	.B2(n514), 
	.B1(\ram[226][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n373));
   AO22CHD U5634 (.O(n4209), 
	.B2(n514), 
	.B1(\ram[226][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n373));
   AO22CHD U5635 (.O(n4210), 
	.B2(n514), 
	.B1(\ram[226][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n373));
   AO22CHD U5636 (.O(n4211), 
	.B2(n514), 
	.B1(\ram[226][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n373));
   AO22CHD U5637 (.O(n4212), 
	.B2(n514), 
	.B1(\ram[226][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n373));
   AO22CHD U5638 (.O(n4213), 
	.B2(n514), 
	.B1(\ram[226][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n373));
   AO22CHD U5639 (.O(n4214), 
	.B2(n516), 
	.B1(\ram[227][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n375));
   AO22CHD U5640 (.O(FE_PHN7456_n4215), 
	.B2(n516), 
	.B1(\ram[227][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n375));
   AO22CHD U5641 (.O(n4216), 
	.B2(n516), 
	.B1(\ram[227][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n375));
   AO22CHD U5642 (.O(n4217), 
	.B2(n516), 
	.B1(\ram[227][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n375));
   AO22CHD U5643 (.O(n4218), 
	.B2(n516), 
	.B1(\ram[227][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n375));
   AO22CHD U5644 (.O(n4219), 
	.B2(n516), 
	.B1(\ram[227][5] ), 
	.A2(n13), 
	.A1(n375));
   AO22CHD U5645 (.O(n4220), 
	.B2(n516), 
	.B1(\ram[227][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n375));
   AO22CHD U5646 (.O(n4221), 
	.B2(n516), 
	.B1(\ram[227][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n375));
   AO22CHD U5647 (.O(n4222), 
	.B2(n516), 
	.B1(\ram[227][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n375));
   AO22CHD U5648 (.O(n4223), 
	.B2(n516), 
	.B1(\ram[227][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n375));
   AO22CHD U5649 (.O(n4224), 
	.B2(n516), 
	.B1(\ram[227][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n375));
   AO22CHD U5650 (.O(n4225), 
	.B2(n516), 
	.B1(\ram[227][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n375));
   AO22CHD U5651 (.O(n4226), 
	.B2(n516), 
	.B1(\ram[227][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n375));
   AO22CHD U5652 (.O(n4227), 
	.B2(n516), 
	.B1(\ram[227][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n375));
   AO22CHD U5653 (.O(n4228), 
	.B2(n516), 
	.B1(\ram[227][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n375));
   AO22CHD U5654 (.O(FE_PHN7454_n4229), 
	.B2(n516), 
	.B1(\ram[227][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n375));
   AO22CHD U5655 (.O(n4230), 
	.B2(n518), 
	.B1(\ram[228][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n377));
   AO22CHD U5656 (.O(n4231), 
	.B2(n518), 
	.B1(\ram[228][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n377));
   AO22CHD U5657 (.O(n4232), 
	.B2(n518), 
	.B1(\ram[228][2] ), 
	.A2(n10), 
	.A1(n377));
   AO22CHD U5658 (.O(n4233), 
	.B2(n518), 
	.B1(\ram[228][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n377));
   AO22CHD U5659 (.O(n4234), 
	.B2(n518), 
	.B1(\ram[228][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n377));
   AO22CHD U5660 (.O(n4235), 
	.B2(n518), 
	.B1(\ram[228][5] ), 
	.A2(n13), 
	.A1(n377));
   AO22CHD U5661 (.O(n4236), 
	.B2(n518), 
	.B1(\ram[228][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n377));
   AO22CHD U5662 (.O(n4237), 
	.B2(n518), 
	.B1(\ram[228][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n377));
   AO22CHD U5663 (.O(n4238), 
	.B2(n518), 
	.B1(\ram[228][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n377));
   AO22CHD U5664 (.O(n4239), 
	.B2(n518), 
	.B1(\ram[228][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n377));
   AO22CHD U5665 (.O(n4240), 
	.B2(n518), 
	.B1(\ram[228][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n377));
   AO22CHD U5666 (.O(n4241), 
	.B2(n518), 
	.B1(\ram[228][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n377));
   AO22CHD U5667 (.O(n4242), 
	.B2(n518), 
	.B1(\ram[228][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n377));
   AO22CHD U5668 (.O(n4243), 
	.B2(n518), 
	.B1(\ram[228][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n377));
   AO22CHD U5669 (.O(n4244), 
	.B2(n518), 
	.B1(\ram[228][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n377));
   AO22CHD U5670 (.O(n4245), 
	.B2(n518), 
	.B1(\ram[228][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n377));
   AO22CHD U5671 (.O(n4246), 
	.B2(n520), 
	.B1(\ram[229][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n378));
   AO22CHD U5672 (.O(n4247), 
	.B2(n520), 
	.B1(\ram[229][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n378));
   AO22CHD U5673 (.O(n4248), 
	.B2(n520), 
	.B1(\ram[229][2] ), 
	.A2(n10), 
	.A1(n378));
   AO22CHD U5674 (.O(n4249), 
	.B2(n520), 
	.B1(FE_PHN4155_ram_229__3_), 
	.A2(FE_OFN50_n11), 
	.A1(n378));
   AO22CHD U5675 (.O(n4250), 
	.B2(n520), 
	.B1(\ram[229][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n378));
   AO22CHD U5676 (.O(n4251), 
	.B2(n520), 
	.B1(\ram[229][5] ), 
	.A2(n13), 
	.A1(n378));
   AO22CHD U5677 (.O(n4252), 
	.B2(n520), 
	.B1(\ram[229][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n378));
   AO22CHD U5678 (.O(n4253), 
	.B2(n520), 
	.B1(\ram[229][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n378));
   AO22CHD U5679 (.O(n4254), 
	.B2(n520), 
	.B1(\ram[229][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n378));
   AO22CHD U5680 (.O(n4255), 
	.B2(n520), 
	.B1(\ram[229][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n378));
   AO22CHD U5681 (.O(n4256), 
	.B2(n520), 
	.B1(\ram[229][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n378));
   AO22CHD U5682 (.O(n4257), 
	.B2(n520), 
	.B1(\ram[229][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n378));
   AO22CHD U5683 (.O(n4258), 
	.B2(n520), 
	.B1(FE_PHN4129_ram_229__12_), 
	.A2(FE_OFN81_n20), 
	.A1(n378));
   AO22CHD U5684 (.O(n4259), 
	.B2(n520), 
	.B1(\ram[229][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n378));
   AO22CHD U5685 (.O(n4260), 
	.B2(n520), 
	.B1(\ram[229][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n378));
   AO22CHD U5686 (.O(n4261), 
	.B2(n520), 
	.B1(\ram[229][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n378));
   AO22CHD U5687 (.O(n4262), 
	.B2(n522), 
	.B1(\ram[230][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n380));
   AO22CHD U5688 (.O(n4263), 
	.B2(n522), 
	.B1(\ram[230][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n380));
   AO22CHD U5689 (.O(n4264), 
	.B2(n522), 
	.B1(\ram[230][2] ), 
	.A2(n10), 
	.A1(n380));
   AO22CHD U5690 (.O(n4265), 
	.B2(n522), 
	.B1(\ram[230][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n380));
   AO22CHD U5691 (.O(n4266), 
	.B2(n522), 
	.B1(\ram[230][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n380));
   AO22CHD U5692 (.O(n4267), 
	.B2(n522), 
	.B1(\ram[230][5] ), 
	.A2(n13), 
	.A1(n380));
   AO22CHD U5693 (.O(n4268), 
	.B2(n522), 
	.B1(\ram[230][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n380));
   AO22CHD U5694 (.O(n4269), 
	.B2(n522), 
	.B1(\ram[230][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n380));
   AO22CHD U5695 (.O(n4270), 
	.B2(n522), 
	.B1(\ram[230][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n380));
   AO22CHD U5696 (.O(n4271), 
	.B2(n522), 
	.B1(\ram[230][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n380));
   AO22CHD U5697 (.O(n4272), 
	.B2(n522), 
	.B1(\ram[230][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n380));
   AO22CHD U5698 (.O(n4273), 
	.B2(n522), 
	.B1(\ram[230][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n380));
   AO22CHD U5699 (.O(n4274), 
	.B2(n522), 
	.B1(\ram[230][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n380));
   AO22CHD U5700 (.O(n4275), 
	.B2(n522), 
	.B1(\ram[230][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n380));
   AO22CHD U5701 (.O(n4276), 
	.B2(n522), 
	.B1(\ram[230][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n380));
   AO22CHD U5702 (.O(n4277), 
	.B2(n522), 
	.B1(\ram[230][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n380));
   AO22CHD U5703 (.O(n4278), 
	.B2(n524), 
	.B1(\ram[231][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n382));
   AO22CHD U5704 (.O(n4279), 
	.B2(n524), 
	.B1(\ram[231][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n382));
   AO22CHD U5705 (.O(n4280), 
	.B2(n524), 
	.B1(\ram[231][2] ), 
	.A2(n10), 
	.A1(n382));
   AO22CHD U5706 (.O(n4281), 
	.B2(n524), 
	.B1(\ram[231][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n382));
   AO22CHD U5707 (.O(n4282), 
	.B2(n524), 
	.B1(\ram[231][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n382));
   AO22CHD U5708 (.O(n4283), 
	.B2(n524), 
	.B1(\ram[231][5] ), 
	.A2(n13), 
	.A1(n382));
   AO22CHD U5709 (.O(n4284), 
	.B2(n524), 
	.B1(\ram[231][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n382));
   AO22CHD U5710 (.O(n4285), 
	.B2(n524), 
	.B1(\ram[231][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n382));
   AO22CHD U5711 (.O(n4286), 
	.B2(n524), 
	.B1(\ram[231][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n382));
   AO22CHD U5712 (.O(n4287), 
	.B2(n524), 
	.B1(\ram[231][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n382));
   AO22CHD U5713 (.O(n4288), 
	.B2(n524), 
	.B1(\ram[231][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n382));
   AO22CHD U5714 (.O(n4289), 
	.B2(n524), 
	.B1(\ram[231][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n382));
   AO22CHD U5715 (.O(n4290), 
	.B2(n524), 
	.B1(\ram[231][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n382));
   AO22CHD U5716 (.O(n4291), 
	.B2(n524), 
	.B1(\ram[231][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n382));
   AO22CHD U5717 (.O(n4292), 
	.B2(n524), 
	.B1(\ram[231][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n382));
   AO22CHD U5718 (.O(n4293), 
	.B2(n524), 
	.B1(\ram[231][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n382));
   AO22CHD U5719 (.O(n4294), 
	.B2(n526), 
	.B1(\ram[232][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n384));
   AO22CHD U5720 (.O(n4295), 
	.B2(n526), 
	.B1(\ram[232][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n384));
   AO22CHD U5721 (.O(n4296), 
	.B2(n526), 
	.B1(\ram[232][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n384));
   AO22CHD U5722 (.O(n4297), 
	.B2(n526), 
	.B1(\ram[232][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n384));
   AO22CHD U5723 (.O(n4298), 
	.B2(n526), 
	.B1(\ram[232][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n384));
   AO22CHD U5724 (.O(n4299), 
	.B2(n526), 
	.B1(\ram[232][5] ), 
	.A2(n13), 
	.A1(n384));
   AO22CHD U5725 (.O(n4300), 
	.B2(n526), 
	.B1(\ram[232][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n384));
   AO22CHD U5726 (.O(n4301), 
	.B2(n526), 
	.B1(\ram[232][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n384));
   AO22CHD U5727 (.O(n4302), 
	.B2(n526), 
	.B1(\ram[232][8] ), 
	.A2(n16), 
	.A1(n384));
   AO22CHD U5728 (.O(n4303), 
	.B2(n526), 
	.B1(\ram[232][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n384));
   AO22CHD U5729 (.O(n4304), 
	.B2(n526), 
	.B1(\ram[232][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n384));
   AO22CHD U5730 (.O(n4305), 
	.B2(n526), 
	.B1(\ram[232][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n384));
   AO22CHD U5731 (.O(n4306), 
	.B2(n526), 
	.B1(\ram[232][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n384));
   AO22CHD U5732 (.O(n4307), 
	.B2(n526), 
	.B1(\ram[232][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n384));
   AO22CHD U5733 (.O(n4308), 
	.B2(n526), 
	.B1(\ram[232][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n384));
   AO22CHD U5734 (.O(n4309), 
	.B2(n526), 
	.B1(\ram[232][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n384));
   AO22CHD U5735 (.O(n4310), 
	.B2(n528), 
	.B1(\ram[233][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n386));
   AO22CHD U5736 (.O(n4311), 
	.B2(n528), 
	.B1(\ram[233][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n386));
   AO22CHD U5737 (.O(n4312), 
	.B2(n528), 
	.B1(\ram[233][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n386));
   AO22CHD U5738 (.O(n4313), 
	.B2(n528), 
	.B1(\ram[233][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n386));
   AO22CHD U5739 (.O(n4314), 
	.B2(n528), 
	.B1(\ram[233][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n386));
   AO22CHD U5740 (.O(n4315), 
	.B2(n528), 
	.B1(\ram[233][5] ), 
	.A2(n13), 
	.A1(n386));
   AO22CHD U5741 (.O(n4316), 
	.B2(n528), 
	.B1(\ram[233][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n386));
   AO22CHD U5742 (.O(n4317), 
	.B2(n528), 
	.B1(\ram[233][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n386));
   AO22CHD U5743 (.O(n4318), 
	.B2(n528), 
	.B1(\ram[233][8] ), 
	.A2(n16), 
	.A1(n386));
   AO22CHD U5744 (.O(n4319), 
	.B2(n528), 
	.B1(\ram[233][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n386));
   AO22CHD U5745 (.O(n4320), 
	.B2(n528), 
	.B1(\ram[233][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n386));
   AO22CHD U5746 (.O(n4321), 
	.B2(n528), 
	.B1(\ram[233][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n386));
   AO22CHD U5747 (.O(n4322), 
	.B2(n528), 
	.B1(\ram[233][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n386));
   AO22CHD U5748 (.O(n4323), 
	.B2(n528), 
	.B1(\ram[233][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n386));
   AO22CHD U5749 (.O(n4324), 
	.B2(n528), 
	.B1(\ram[233][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n386));
   AO22CHD U5750 (.O(n4325), 
	.B2(n528), 
	.B1(\ram[233][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n386));
   AO22CHD U5751 (.O(n4326), 
	.B2(n530), 
	.B1(\ram[234][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n388));
   AO22CHD U5752 (.O(n4327), 
	.B2(n530), 
	.B1(\ram[234][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n388));
   AO22CHD U5753 (.O(n4328), 
	.B2(n530), 
	.B1(\ram[234][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n388));
   AO22CHD U5754 (.O(n4329), 
	.B2(n530), 
	.B1(\ram[234][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n388));
   AO22CHD U5755 (.O(n4330), 
	.B2(n530), 
	.B1(\ram[234][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n388));
   AO22CHD U5756 (.O(n4331), 
	.B2(n530), 
	.B1(\ram[234][5] ), 
	.A2(n13), 
	.A1(n388));
   AO22CHD U5757 (.O(n4332), 
	.B2(n530), 
	.B1(\ram[234][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n388));
   AO22CHD U5758 (.O(n4333), 
	.B2(n530), 
	.B1(\ram[234][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n388));
   AO22CHD U5759 (.O(n4334), 
	.B2(n530), 
	.B1(\ram[234][8] ), 
	.A2(n16), 
	.A1(n388));
   AO22CHD U5760 (.O(n4335), 
	.B2(n530), 
	.B1(\ram[234][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n388));
   AO22CHD U5761 (.O(n4336), 
	.B2(n530), 
	.B1(\ram[234][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n388));
   AO22CHD U5762 (.O(n4337), 
	.B2(n530), 
	.B1(\ram[234][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n388));
   AO22CHD U5763 (.O(n4338), 
	.B2(n530), 
	.B1(\ram[234][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n388));
   AO22CHD U5764 (.O(n4339), 
	.B2(n530), 
	.B1(\ram[234][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n388));
   AO22CHD U5765 (.O(n4340), 
	.B2(n530), 
	.B1(\ram[234][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n388));
   AO22CHD U5766 (.O(n4341), 
	.B2(n530), 
	.B1(\ram[234][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n388));
   AO22CHD U5767 (.O(n4342), 
	.B2(n532), 
	.B1(\ram[235][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n390));
   AO22CHD U5768 (.O(n4343), 
	.B2(n532), 
	.B1(\ram[235][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n390));
   AO22CHD U5769 (.O(n4344), 
	.B2(n532), 
	.B1(\ram[235][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n390));
   AO22CHD U5770 (.O(n4345), 
	.B2(n532), 
	.B1(\ram[235][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n390));
   AO22CHD U5771 (.O(n4346), 
	.B2(n532), 
	.B1(\ram[235][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n390));
   AO22CHD U5772 (.O(n4347), 
	.B2(n532), 
	.B1(\ram[235][5] ), 
	.A2(n13), 
	.A1(n390));
   AO22CHD U5773 (.O(n4348), 
	.B2(n532), 
	.B1(\ram[235][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n390));
   AO22CHD U5774 (.O(n4349), 
	.B2(n532), 
	.B1(\ram[235][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n390));
   AO22CHD U5775 (.O(n4350), 
	.B2(n532), 
	.B1(\ram[235][8] ), 
	.A2(n16), 
	.A1(n390));
   AO22CHD U5776 (.O(n4351), 
	.B2(n532), 
	.B1(\ram[235][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n390));
   AO22CHD U5777 (.O(n4352), 
	.B2(n532), 
	.B1(\ram[235][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n390));
   AO22CHD U5778 (.O(n4353), 
	.B2(n532), 
	.B1(\ram[235][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n390));
   AO22CHD U5779 (.O(n4354), 
	.B2(n532), 
	.B1(\ram[235][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n390));
   AO22CHD U5780 (.O(n4355), 
	.B2(n532), 
	.B1(\ram[235][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n390));
   AO22CHD U5781 (.O(n4356), 
	.B2(n532), 
	.B1(\ram[235][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n390));
   AO22CHD U5782 (.O(n4357), 
	.B2(n532), 
	.B1(\ram[235][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n390));
   AO22CHD U5783 (.O(n4358), 
	.B2(n534), 
	.B1(\ram[236][0] ), 
	.A2(n6), 
	.A1(n392));
   AO22CHD U5784 (.O(n4359), 
	.B2(n534), 
	.B1(\ram[236][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n392));
   AO22CHD U5785 (.O(n4360), 
	.B2(n534), 
	.B1(\ram[236][2] ), 
	.A2(n10), 
	.A1(n392));
   AO22CHD U5786 (.O(n4361), 
	.B2(n534), 
	.B1(\ram[236][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n392));
   AO22CHD U5787 (.O(n4362), 
	.B2(n534), 
	.B1(\ram[236][4] ), 
	.A2(n12), 
	.A1(n392));
   AO22CHD U5788 (.O(n4363), 
	.B2(n534), 
	.B1(\ram[236][5] ), 
	.A2(n13), 
	.A1(n392));
   AO22CHD U5789 (.O(n4364), 
	.B2(n534), 
	.B1(\ram[236][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n392));
   AO22CHD U5790 (.O(n4365), 
	.B2(n534), 
	.B1(\ram[236][7] ), 
	.A2(n15), 
	.A1(n392));
   AO22CHD U5791 (.O(n4366), 
	.B2(n534), 
	.B1(\ram[236][8] ), 
	.A2(n16), 
	.A1(n392));
   AO22CHD U5792 (.O(n4367), 
	.B2(n534), 
	.B1(\ram[236][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n392));
   AO22CHD U5793 (.O(n4368), 
	.B2(n534), 
	.B1(\ram[236][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n392));
   AO22CHD U5794 (.O(n4369), 
	.B2(n534), 
	.B1(\ram[236][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n392));
   AO22CHD U5795 (.O(n4370), 
	.B2(n534), 
	.B1(\ram[236][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n392));
   AO22CHD U5796 (.O(n4371), 
	.B2(n534), 
	.B1(\ram[236][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n392));
   AO22CHD U5797 (.O(n4372), 
	.B2(n534), 
	.B1(\ram[236][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n392));
   AO22CHD U5798 (.O(n4373), 
	.B2(n534), 
	.B1(\ram[236][15] ), 
	.A2(n23), 
	.A1(n392));
   AO22CHD U5799 (.O(n4374), 
	.B2(n536), 
	.B1(\ram[237][0] ), 
	.A2(n6), 
	.A1(n394));
   AO22CHD U5800 (.O(n4375), 
	.B2(n536), 
	.B1(\ram[237][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n394));
   AO22CHD U5801 (.O(n4376), 
	.B2(n536), 
	.B1(\ram[237][2] ), 
	.A2(n10), 
	.A1(n394));
   AO22CHD U5802 (.O(n4377), 
	.B2(n536), 
	.B1(\ram[237][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n394));
   AO22CHD U5803 (.O(n4378), 
	.B2(n536), 
	.B1(\ram[237][4] ), 
	.A2(n12), 
	.A1(n394));
   AO22CHD U5804 (.O(n4379), 
	.B2(n536), 
	.B1(\ram[237][5] ), 
	.A2(n13), 
	.A1(n394));
   AO22CHD U5805 (.O(n4380), 
	.B2(n536), 
	.B1(\ram[237][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n394));
   AO22CHD U5806 (.O(n4381), 
	.B2(n536), 
	.B1(FE_PHN4172_ram_237__7_), 
	.A2(n15), 
	.A1(n394));
   AO22CHD U5807 (.O(n4382), 
	.B2(n536), 
	.B1(\ram[237][8] ), 
	.A2(n16), 
	.A1(n394));
   AO22CHD U5808 (.O(n4383), 
	.B2(n536), 
	.B1(\ram[237][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n394));
   AO22CHD U5809 (.O(n4384), 
	.B2(n536), 
	.B1(\ram[237][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n394));
   AO22CHD U5810 (.O(n4385), 
	.B2(n536), 
	.B1(\ram[237][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n394));
   AO22CHD U5811 (.O(n4386), 
	.B2(n536), 
	.B1(\ram[237][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n394));
   AO22CHD U5812 (.O(n4387), 
	.B2(n536), 
	.B1(\ram[237][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n394));
   AO22CHD U5813 (.O(n4388), 
	.B2(n536), 
	.B1(\ram[237][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n394));
   AO22CHD U5814 (.O(n4389), 
	.B2(n536), 
	.B1(\ram[237][15] ), 
	.A2(n23), 
	.A1(n394));
   AO22CHD U5815 (.O(n4390), 
	.B2(n538), 
	.B1(FE_PHN4224_ram_238__0_), 
	.A2(n6), 
	.A1(n396));
   AO22CHD U5816 (.O(n4391), 
	.B2(n538), 
	.B1(\ram[238][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n396));
   AO22CHD U5817 (.O(n4392), 
	.B2(n538), 
	.B1(\ram[238][2] ), 
	.A2(n10), 
	.A1(n396));
   AO22CHD U5818 (.O(n4393), 
	.B2(n538), 
	.B1(\ram[238][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n396));
   AO22CHD U5819 (.O(n4394), 
	.B2(n538), 
	.B1(\ram[238][4] ), 
	.A2(n12), 
	.A1(n396));
   AO22CHD U5820 (.O(n4395), 
	.B2(n538), 
	.B1(\ram[238][5] ), 
	.A2(n13), 
	.A1(n396));
   AO22CHD U5821 (.O(n4396), 
	.B2(n538), 
	.B1(\ram[238][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n396));
   AO22CHD U5822 (.O(n4397), 
	.B2(n538), 
	.B1(\ram[238][7] ), 
	.A2(n15), 
	.A1(n396));
   AO22CHD U5823 (.O(n4398), 
	.B2(n538), 
	.B1(\ram[238][8] ), 
	.A2(n16), 
	.A1(n396));
   AO22CHD U5824 (.O(n4399), 
	.B2(n538), 
	.B1(\ram[238][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n396));
   AO22CHD U5825 (.O(n4400), 
	.B2(n538), 
	.B1(\ram[238][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n396));
   AO22CHD U5826 (.O(n4401), 
	.B2(n538), 
	.B1(\ram[238][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n396));
   AO22CHD U5827 (.O(n4402), 
	.B2(n538), 
	.B1(\ram[238][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n396));
   AO22CHD U5828 (.O(n4403), 
	.B2(n538), 
	.B1(\ram[238][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n396));
   AO22CHD U5829 (.O(n4404), 
	.B2(n538), 
	.B1(\ram[238][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n396));
   AO22CHD U5830 (.O(n4405), 
	.B2(n538), 
	.B1(\ram[238][15] ), 
	.A2(n23), 
	.A1(n396));
   AO22CHD U5831 (.O(n4406), 
	.B2(n540), 
	.B1(\ram[239][0] ), 
	.A2(n6), 
	.A1(n398));
   AO22CHD U5832 (.O(n4407), 
	.B2(n540), 
	.B1(\ram[239][1] ), 
	.A2(FE_OFN45_n9), 
	.A1(n398));
   AO22CHD U5833 (.O(n4408), 
	.B2(n540), 
	.B1(\ram[239][2] ), 
	.A2(n10), 
	.A1(n398));
   AO22CHD U5834 (.O(n4409), 
	.B2(n540), 
	.B1(\ram[239][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n398));
   AO22CHD U5835 (.O(n4410), 
	.B2(n540), 
	.B1(\ram[239][4] ), 
	.A2(n12), 
	.A1(n398));
   AO22CHD U5836 (.O(n4411), 
	.B2(n540), 
	.B1(\ram[239][5] ), 
	.A2(n13), 
	.A1(n398));
   AO22CHD U5837 (.O(n4412), 
	.B2(n540), 
	.B1(\ram[239][6] ), 
	.A2(FE_OFN59_n14), 
	.A1(n398));
   AO22CHD U5838 (.O(n4413), 
	.B2(n540), 
	.B1(\ram[239][7] ), 
	.A2(n15), 
	.A1(n398));
   AO22CHD U5839 (.O(n4414), 
	.B2(n540), 
	.B1(\ram[239][8] ), 
	.A2(n16), 
	.A1(n398));
   AO22CHD U5840 (.O(n4415), 
	.B2(n540), 
	.B1(\ram[239][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n398));
   AO22CHD U5841 (.O(n4416), 
	.B2(n540), 
	.B1(\ram[239][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n398));
   AO22CHD U5842 (.O(n4417), 
	.B2(n540), 
	.B1(\ram[239][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n398));
   AO22CHD U5843 (.O(n4418), 
	.B2(n540), 
	.B1(\ram[239][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n398));
   AO22CHD U5844 (.O(n4419), 
	.B2(n540), 
	.B1(\ram[239][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n398));
   AO22CHD U5845 (.O(n4420), 
	.B2(n540), 
	.B1(\ram[239][14] ), 
	.A2(FE_OFN86_n22), 
	.A1(n398));
   AO22CHD U5846 (.O(n4421), 
	.B2(n540), 
	.B1(\ram[239][15] ), 
	.A2(n23), 
	.A1(n398));
   AO22CHD U5847 (.O(n4422), 
	.B2(n542), 
	.B1(\ram[240][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n400));
   AO22CHD U5848 (.O(n4423), 
	.B2(n542), 
	.B1(\ram[240][1] ), 
	.A2(n9), 
	.A1(n400));
   AO22CHD U5849 (.O(n4424), 
	.B2(n542), 
	.B1(\ram[240][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n400));
   AO22CHD U5850 (.O(n4425), 
	.B2(n542), 
	.B1(\ram[240][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n400));
   AO22CHD U5851 (.O(n4426), 
	.B2(n542), 
	.B1(\ram[240][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n400));
   AO22CHD U5852 (.O(n4427), 
	.B2(n542), 
	.B1(\ram[240][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n400));
   AO22CHD U5853 (.O(n4428), 
	.B2(n542), 
	.B1(\ram[240][6] ), 
	.A2(n14), 
	.A1(n400));
   AO22CHD U5854 (.O(n4429), 
	.B2(n542), 
	.B1(\ram[240][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n400));
   AO22CHD U5855 (.O(n4430), 
	.B2(n542), 
	.B1(\ram[240][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n400));
   AO22CHD U5856 (.O(n4431), 
	.B2(n542), 
	.B1(\ram[240][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n400));
   AO22CHD U5857 (.O(n4432), 
	.B2(n542), 
	.B1(\ram[240][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n400));
   AO22CHD U5858 (.O(n4433), 
	.B2(n542), 
	.B1(\ram[240][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n400));
   AO22CHD U5859 (.O(n4434), 
	.B2(n542), 
	.B1(\ram[240][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n400));
   AO22CHD U5860 (.O(n4435), 
	.B2(n542), 
	.B1(\ram[240][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n400));
   AO22CHD U5861 (.O(n4436), 
	.B2(n542), 
	.B1(\ram[240][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n400));
   AO22CHD U5862 (.O(n4437), 
	.B2(n542), 
	.B1(\ram[240][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n400));
   AO22CHD U5863 (.O(n4438), 
	.B2(n547), 
	.B1(FE_PHN2371_ram_241__0_), 
	.A2(FE_OFN43_n6), 
	.A1(n402));
   AO22CHD U5864 (.O(n4439), 
	.B2(n547), 
	.B1(FE_PHN165_ram_241__1_), 
	.A2(n9), 
	.A1(n402));
   AO22CHD U5865 (.O(n4440), 
	.B2(n547), 
	.B1(\ram[241][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n402));
   AO22CHD U5866 (.O(n4441), 
	.B2(n547), 
	.B1(\ram[241][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n402));
   AO22CHD U5867 (.O(n4442), 
	.B2(n547), 
	.B1(\ram[241][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n402));
   AO22CHD U5868 (.O(n4443), 
	.B2(n547), 
	.B1(\ram[241][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n402));
   AO22CHD U5869 (.O(n4444), 
	.B2(n547), 
	.B1(\ram[241][6] ), 
	.A2(n14), 
	.A1(n402));
   AO22CHD U5870 (.O(n4445), 
	.B2(n547), 
	.B1(\ram[241][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n402));
   AO22CHD U5871 (.O(n4446), 
	.B2(n547), 
	.B1(\ram[241][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n402));
   AO22CHD U5872 (.O(n4447), 
	.B2(n547), 
	.B1(\ram[241][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n402));
   AO22CHD U5873 (.O(n4448), 
	.B2(n547), 
	.B1(\ram[241][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n402));
   AO22CHD U5874 (.O(n4449), 
	.B2(n547), 
	.B1(\ram[241][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n402));
   AO22CHD U5875 (.O(n4450), 
	.B2(n547), 
	.B1(\ram[241][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n402));
   AO22CHD U5876 (.O(n4451), 
	.B2(n547), 
	.B1(\ram[241][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n402));
   AO22CHD U5877 (.O(n4452), 
	.B2(n547), 
	.B1(\ram[241][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n402));
   AO22CHD U5878 (.O(n4453), 
	.B2(n547), 
	.B1(\ram[241][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n402));
   AO22CHD U5879 (.O(n4454), 
	.B2(n550), 
	.B1(\ram[242][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n404));
   AO22CHD U5880 (.O(n4455), 
	.B2(n550), 
	.B1(\ram[242][1] ), 
	.A2(n9), 
	.A1(n404));
   AO22CHD U5881 (.O(n4456), 
	.B2(n550), 
	.B1(\ram[242][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n404));
   AO22CHD U5882 (.O(n4457), 
	.B2(n550), 
	.B1(\ram[242][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n404));
   AO22CHD U5883 (.O(n4458), 
	.B2(n550), 
	.B1(\ram[242][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n404));
   AO22CHD U5884 (.O(n4459), 
	.B2(n550), 
	.B1(\ram[242][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n404));
   AO22CHD U5885 (.O(n4460), 
	.B2(n550), 
	.B1(\ram[242][6] ), 
	.A2(n14), 
	.A1(n404));
   AO22CHD U5886 (.O(n4461), 
	.B2(n550), 
	.B1(\ram[242][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n404));
   AO22CHD U5887 (.O(n4462), 
	.B2(n550), 
	.B1(\ram[242][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n404));
   AO22CHD U5888 (.O(n4463), 
	.B2(n550), 
	.B1(\ram[242][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n404));
   AO22CHD U5889 (.O(n4464), 
	.B2(n550), 
	.B1(\ram[242][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n404));
   AO22CHD U5890 (.O(n4465), 
	.B2(n550), 
	.B1(\ram[242][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n404));
   AO22CHD U5891 (.O(n4466), 
	.B2(n550), 
	.B1(\ram[242][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n404));
   AO22CHD U5892 (.O(n4467), 
	.B2(n550), 
	.B1(\ram[242][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n404));
   AO22CHD U5893 (.O(n4468), 
	.B2(n550), 
	.B1(\ram[242][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n404));
   AO22CHD U5894 (.O(n4469), 
	.B2(n550), 
	.B1(\ram[242][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n404));
   AO22CHD U5895 (.O(n4470), 
	.B2(n553), 
	.B1(\ram[243][0] ), 
	.A2(FE_OFN43_n6), 
	.A1(n406));
   AO22CHD U5896 (.O(n4471), 
	.B2(n553), 
	.B1(\ram[243][1] ), 
	.A2(n9), 
	.A1(n406));
   AO22CHD U5897 (.O(n4472), 
	.B2(n553), 
	.B1(\ram[243][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n406));
   AO22CHD U5898 (.O(n4473), 
	.B2(n553), 
	.B1(\ram[243][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n406));
   AO22CHD U5899 (.O(n4474), 
	.B2(n553), 
	.B1(\ram[243][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n406));
   AO22CHD U5900 (.O(n4475), 
	.B2(n553), 
	.B1(\ram[243][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n406));
   AO22CHD U5901 (.O(n4476), 
	.B2(n553), 
	.B1(\ram[243][6] ), 
	.A2(n14), 
	.A1(n406));
   AO22CHD U5902 (.O(n4477), 
	.B2(n553), 
	.B1(\ram[243][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n406));
   AO22CHD U5903 (.O(n4478), 
	.B2(n553), 
	.B1(\ram[243][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n406));
   AO22CHD U5904 (.O(n4479), 
	.B2(n553), 
	.B1(\ram[243][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n406));
   AO22CHD U5905 (.O(n4480), 
	.B2(n553), 
	.B1(\ram[243][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n406));
   AO22CHD U5906 (.O(n4481), 
	.B2(n553), 
	.B1(\ram[243][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n406));
   AO22CHD U5907 (.O(n4482), 
	.B2(n553), 
	.B1(\ram[243][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n406));
   AO22CHD U5908 (.O(n4483), 
	.B2(n553), 
	.B1(\ram[243][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n406));
   AO22CHD U5909 (.O(n4484), 
	.B2(n553), 
	.B1(\ram[243][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n406));
   AO22CHD U5910 (.O(n4485), 
	.B2(n553), 
	.B1(\ram[243][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n406));
   AO22CHD U5911 (.O(n4486), 
	.B2(n556), 
	.B1(\ram[244][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n408));
   AO22CHD U5912 (.O(n4487), 
	.B2(n556), 
	.B1(\ram[244][1] ), 
	.A2(n9), 
	.A1(n408));
   AO22CHD U5913 (.O(n4488), 
	.B2(n556), 
	.B1(\ram[244][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n408));
   AO22CHD U5914 (.O(n4489), 
	.B2(n556), 
	.B1(\ram[244][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n408));
   AO22CHD U5915 (.O(n4490), 
	.B2(n556), 
	.B1(\ram[244][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n408));
   AO22CHD U5916 (.O(n4491), 
	.B2(n556), 
	.B1(\ram[244][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n408));
   AO22CHD U5917 (.O(n4492), 
	.B2(n556), 
	.B1(\ram[244][6] ), 
	.A2(n14), 
	.A1(n408));
   AO22CHD U5918 (.O(n4493), 
	.B2(n556), 
	.B1(\ram[244][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n408));
   AO22CHD U5919 (.O(n4494), 
	.B2(n556), 
	.B1(\ram[244][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n408));
   AO22CHD U5920 (.O(n4495), 
	.B2(n556), 
	.B1(\ram[244][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n408));
   AO22CHD U5921 (.O(n4496), 
	.B2(n556), 
	.B1(FE_PHN3013_ram_244__10_), 
	.A2(FE_OFN75_n18), 
	.A1(n408));
   AO22CHD U5922 (.O(n4497), 
	.B2(n556), 
	.B1(\ram[244][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n408));
   AO22CHD U5923 (.O(n4498), 
	.B2(n556), 
	.B1(\ram[244][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n408));
   AO22CHD U5924 (.O(n4499), 
	.B2(n556), 
	.B1(\ram[244][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n408));
   AO22CHD U5925 (.O(n4500), 
	.B2(n556), 
	.B1(\ram[244][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n408));
   AO22CHD U5926 (.O(n4501), 
	.B2(n556), 
	.B1(\ram[244][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n408));
   AO22CHD U5927 (.O(n4502), 
	.B2(n559), 
	.B1(\ram[245][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n410));
   AO22CHD U5928 (.O(n4503), 
	.B2(n559), 
	.B1(\ram[245][1] ), 
	.A2(n9), 
	.A1(n410));
   AO22CHD U5929 (.O(n4504), 
	.B2(n559), 
	.B1(\ram[245][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n410));
   AO22CHD U5930 (.O(n4505), 
	.B2(n559), 
	.B1(\ram[245][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n410));
   AO22CHD U5931 (.O(n4506), 
	.B2(n559), 
	.B1(\ram[245][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n410));
   AO22CHD U5932 (.O(n4507), 
	.B2(n559), 
	.B1(\ram[245][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n410));
   AO22CHD U5933 (.O(n4508), 
	.B2(n559), 
	.B1(\ram[245][6] ), 
	.A2(n14), 
	.A1(n410));
   AO22CHD U5934 (.O(n4509), 
	.B2(n559), 
	.B1(\ram[245][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n410));
   AO22CHD U5935 (.O(n4510), 
	.B2(n559), 
	.B1(\ram[245][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n410));
   AO22CHD U5936 (.O(n4511), 
	.B2(n559), 
	.B1(\ram[245][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n410));
   AO22CHD U5937 (.O(n4512), 
	.B2(n559), 
	.B1(\ram[245][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n410));
   AO22CHD U5938 (.O(n4513), 
	.B2(n559), 
	.B1(\ram[245][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n410));
   AO22CHD U5939 (.O(n4514), 
	.B2(n559), 
	.B1(\ram[245][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n410));
   AO22CHD U5940 (.O(n4515), 
	.B2(n559), 
	.B1(\ram[245][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n410));
   AO22CHD U5941 (.O(n4516), 
	.B2(n559), 
	.B1(\ram[245][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n410));
   AO22CHD U5942 (.O(n4517), 
	.B2(n559), 
	.B1(\ram[245][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n410));
   AO22CHD U5943 (.O(n4518), 
	.B2(n561), 
	.B1(\ram[246][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n411));
   AO22CHD U5944 (.O(n4519), 
	.B2(n561), 
	.B1(\ram[246][1] ), 
	.A2(n9), 
	.A1(n411));
   AO22CHD U5945 (.O(n4520), 
	.B2(n561), 
	.B1(\ram[246][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n411));
   AO22CHD U5946 (.O(n4521), 
	.B2(n561), 
	.B1(\ram[246][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n411));
   AO22CHD U5947 (.O(n4522), 
	.B2(n561), 
	.B1(\ram[246][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n411));
   AO22CHD U5948 (.O(n4523), 
	.B2(n561), 
	.B1(\ram[246][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n411));
   AO22CHD U5949 (.O(n4524), 
	.B2(n561), 
	.B1(\ram[246][6] ), 
	.A2(n14), 
	.A1(n411));
   AO22CHD U5950 (.O(n4525), 
	.B2(n561), 
	.B1(\ram[246][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n411));
   AO22CHD U5951 (.O(n4526), 
	.B2(n561), 
	.B1(\ram[246][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n411));
   AO22CHD U5952 (.O(n4527), 
	.B2(n561), 
	.B1(\ram[246][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n411));
   AO22CHD U5953 (.O(n4528), 
	.B2(n561), 
	.B1(\ram[246][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n411));
   AO22CHD U5954 (.O(n4529), 
	.B2(n561), 
	.B1(\ram[246][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n411));
   AO22CHD U5955 (.O(n4530), 
	.B2(n561), 
	.B1(\ram[246][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n411));
   AO22CHD U5956 (.O(n4531), 
	.B2(n561), 
	.B1(\ram[246][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n411));
   AO22CHD U5957 (.O(n4532), 
	.B2(n561), 
	.B1(\ram[246][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n411));
   AO22CHD U5958 (.O(n4533), 
	.B2(n561), 
	.B1(\ram[246][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n411));
   AO22CHD U5959 (.O(n4534), 
	.B2(n563), 
	.B1(\ram[247][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n413));
   AO22CHD U5960 (.O(n4535), 
	.B2(n563), 
	.B1(\ram[247][1] ), 
	.A2(n9), 
	.A1(n413));
   AO22CHD U5961 (.O(n4536), 
	.B2(n563), 
	.B1(\ram[247][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n413));
   AO22CHD U5962 (.O(n4537), 
	.B2(n563), 
	.B1(\ram[247][3] ), 
	.A2(FE_OFN51_n11), 
	.A1(n413));
   AO22CHD U5963 (.O(n4538), 
	.B2(n563), 
	.B1(\ram[247][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n413));
   AO22CHD U5964 (.O(n4539), 
	.B2(n563), 
	.B1(\ram[247][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n413));
   AO22CHD U5965 (.O(n4540), 
	.B2(n563), 
	.B1(\ram[247][6] ), 
	.A2(n14), 
	.A1(n413));
   AO22CHD U5966 (.O(n4541), 
	.B2(n563), 
	.B1(\ram[247][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n413));
   AO22CHD U5967 (.O(n4542), 
	.B2(n563), 
	.B1(\ram[247][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n413));
   AO22CHD U5968 (.O(n4543), 
	.B2(n563), 
	.B1(\ram[247][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n413));
   AO22CHD U5969 (.O(n4544), 
	.B2(n563), 
	.B1(\ram[247][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n413));
   AO22CHD U5970 (.O(n4545), 
	.B2(n563), 
	.B1(\ram[247][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n413));
   AO22CHD U5971 (.O(n4546), 
	.B2(n563), 
	.B1(\ram[247][12] ), 
	.A2(FE_OFN82_n20), 
	.A1(n413));
   AO22CHD U5972 (.O(n4547), 
	.B2(n563), 
	.B1(\ram[247][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n413));
   AO22CHD U5973 (.O(n4548), 
	.B2(n563), 
	.B1(\ram[247][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n413));
   AO22CHD U5974 (.O(n4549), 
	.B2(n563), 
	.B1(\ram[247][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n413));
   AO22CHD U5975 (.O(n4550), 
	.B2(n565), 
	.B1(\ram[248][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n415));
   AO22CHD U5976 (.O(n4551), 
	.B2(n565), 
	.B1(\ram[248][1] ), 
	.A2(n9), 
	.A1(n415));
   AO22CHD U5977 (.O(n4552), 
	.B2(n565), 
	.B1(\ram[248][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n415));
   AO22CHD U5978 (.O(n4553), 
	.B2(n565), 
	.B1(\ram[248][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n415));
   AO22CHD U5979 (.O(n4554), 
	.B2(n565), 
	.B1(\ram[248][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n415));
   AO22CHD U5980 (.O(n4555), 
	.B2(n565), 
	.B1(\ram[248][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n415));
   AO22CHD U5981 (.O(n4556), 
	.B2(n565), 
	.B1(\ram[248][6] ), 
	.A2(n14), 
	.A1(n415));
   AO22CHD U5982 (.O(n4557), 
	.B2(n565), 
	.B1(\ram[248][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n415));
   AO22CHD U5983 (.O(n4558), 
	.B2(n565), 
	.B1(\ram[248][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n415));
   AO22CHD U5984 (.O(n4559), 
	.B2(n565), 
	.B1(\ram[248][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n415));
   AO22CHD U5985 (.O(n4560), 
	.B2(n565), 
	.B1(\ram[248][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n415));
   AO22CHD U5986 (.O(n4561), 
	.B2(n565), 
	.B1(\ram[248][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n415));
   AO22CHD U5987 (.O(n4562), 
	.B2(n565), 
	.B1(\ram[248][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n415));
   AO22CHD U5988 (.O(n4563), 
	.B2(n565), 
	.B1(\ram[248][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n415));
   AO22CHD U5989 (.O(n4564), 
	.B2(n565), 
	.B1(\ram[248][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n415));
   AO22CHD U5990 (.O(n4565), 
	.B2(n565), 
	.B1(\ram[248][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n415));
   AO22CHD U5991 (.O(n4566), 
	.B2(n568), 
	.B1(\ram[249][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n417));
   AO22CHD U5992 (.O(n4567), 
	.B2(n568), 
	.B1(\ram[249][1] ), 
	.A2(n9), 
	.A1(n417));
   AO22CHD U5993 (.O(n4568), 
	.B2(n568), 
	.B1(\ram[249][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n417));
   AO22CHD U5994 (.O(n4569), 
	.B2(n568), 
	.B1(\ram[249][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n417));
   AO22CHD U5995 (.O(n4570), 
	.B2(n568), 
	.B1(\ram[249][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n417));
   AO22CHD U5996 (.O(n4571), 
	.B2(n568), 
	.B1(\ram[249][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n417));
   AO22CHD U5997 (.O(n4572), 
	.B2(n568), 
	.B1(\ram[249][6] ), 
	.A2(n14), 
	.A1(n417));
   AO22CHD U5998 (.O(n4573), 
	.B2(n568), 
	.B1(\ram[249][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n417));
   AO22CHD U5999 (.O(n4574), 
	.B2(n568), 
	.B1(\ram[249][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n417));
   AO22CHD U6000 (.O(n4575), 
	.B2(n568), 
	.B1(\ram[249][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n417));
   AO22CHD U6001 (.O(n4576), 
	.B2(n568), 
	.B1(\ram[249][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n417));
   AO22CHD U6002 (.O(n4577), 
	.B2(n568), 
	.B1(\ram[249][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n417));
   AO22CHD U6003 (.O(n4578), 
	.B2(n568), 
	.B1(FE_PHN871_ram_249__12_), 
	.A2(FE_OFN81_n20), 
	.A1(n417));
   AO22CHD U6004 (.O(n4579), 
	.B2(n568), 
	.B1(\ram[249][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n417));
   AO22CHD U6005 (.O(n4580), 
	.B2(n568), 
	.B1(\ram[249][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n417));
   AO22CHD U6006 (.O(n4581), 
	.B2(n568), 
	.B1(\ram[249][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n417));
   AO22CHD U6007 (.O(n4582), 
	.B2(n570), 
	.B1(\ram[250][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n419));
   AO22CHD U6008 (.O(n4583), 
	.B2(n570), 
	.B1(FE_PHN2995_ram_250__1_), 
	.A2(n9), 
	.A1(n419));
   AO22CHD U6009 (.O(n4584), 
	.B2(n570), 
	.B1(\ram[250][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n419));
   AO22CHD U6010 (.O(n4585), 
	.B2(n570), 
	.B1(\ram[250][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n419));
   AO22CHD U6011 (.O(n4586), 
	.B2(n570), 
	.B1(\ram[250][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n419));
   AO22CHD U6012 (.O(n4587), 
	.B2(n570), 
	.B1(\ram[250][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n419));
   AO22CHD U6013 (.O(n4588), 
	.B2(n570), 
	.B1(\ram[250][6] ), 
	.A2(n14), 
	.A1(n419));
   AO22CHD U6014 (.O(n4589), 
	.B2(n570), 
	.B1(\ram[250][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n419));
   AO22CHD U6015 (.O(n4590), 
	.B2(n570), 
	.B1(\ram[250][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n419));
   AO22CHD U6016 (.O(n4591), 
	.B2(n570), 
	.B1(\ram[250][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n419));
   AO22CHD U6017 (.O(n4592), 
	.B2(n570), 
	.B1(\ram[250][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n419));
   AO22CHD U6018 (.O(n4593), 
	.B2(n570), 
	.B1(\ram[250][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n419));
   AO22CHD U6019 (.O(n4594), 
	.B2(n570), 
	.B1(\ram[250][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n419));
   AO22CHD U6020 (.O(n4595), 
	.B2(n570), 
	.B1(\ram[250][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n419));
   AO22CHD U6021 (.O(n4596), 
	.B2(n570), 
	.B1(\ram[250][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n419));
   AO22CHD U6022 (.O(n4597), 
	.B2(n570), 
	.B1(\ram[250][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n419));
   AO22CHD U6023 (.O(n4598), 
	.B2(n572), 
	.B1(\ram[251][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n421));
   AO22CHD U6024 (.O(n4599), 
	.B2(n572), 
	.B1(\ram[251][1] ), 
	.A2(n9), 
	.A1(n421));
   AO22CHD U6025 (.O(n4600), 
	.B2(n572), 
	.B1(\ram[251][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n421));
   AO22CHD U6026 (.O(n4601), 
	.B2(n572), 
	.B1(\ram[251][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n421));
   AO22CHD U6027 (.O(n4602), 
	.B2(n572), 
	.B1(\ram[251][4] ), 
	.A2(FE_OFN53_n12), 
	.A1(n421));
   AO22CHD U6028 (.O(n4603), 
	.B2(n572), 
	.B1(\ram[251][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n421));
   AO22CHD U6029 (.O(n4604), 
	.B2(n572), 
	.B1(\ram[251][6] ), 
	.A2(n14), 
	.A1(n421));
   AO22CHD U6030 (.O(n4605), 
	.B2(n572), 
	.B1(\ram[251][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n421));
   AO22CHD U6031 (.O(n4606), 
	.B2(n572), 
	.B1(\ram[251][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n421));
   AO22CHD U6032 (.O(n4607), 
	.B2(n572), 
	.B1(\ram[251][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n421));
   AO22CHD U6033 (.O(n4608), 
	.B2(n572), 
	.B1(\ram[251][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n421));
   AO22CHD U6034 (.O(n4609), 
	.B2(n572), 
	.B1(\ram[251][11] ), 
	.A2(FE_OFN77_n19), 
	.A1(n421));
   AO22CHD U6035 (.O(n4610), 
	.B2(n572), 
	.B1(\ram[251][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n421));
   AO22CHD U6036 (.O(n4611), 
	.B2(n572), 
	.B1(\ram[251][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n421));
   AO22CHD U6037 (.O(n4612), 
	.B2(n572), 
	.B1(\ram[251][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n421));
   AO22CHD U6038 (.O(n4613), 
	.B2(n572), 
	.B1(\ram[251][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n421));
   AO22CHD U6039 (.O(n4614), 
	.B2(n574), 
	.B1(\ram[252][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n423));
   AO22CHD U6040 (.O(n4615), 
	.B2(n574), 
	.B1(\ram[252][1] ), 
	.A2(n9), 
	.A1(n423));
   AO22CHD U6041 (.O(n4616), 
	.B2(n574), 
	.B1(\ram[252][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n423));
   AO22CHD U6042 (.O(n4617), 
	.B2(n574), 
	.B1(\ram[252][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n423));
   AO22CHD U6043 (.O(n4618), 
	.B2(n574), 
	.B1(\ram[252][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n423));
   AO22CHD U6044 (.O(n4619), 
	.B2(n574), 
	.B1(\ram[252][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n423));
   AO22CHD U6045 (.O(n4620), 
	.B2(n574), 
	.B1(\ram[252][6] ), 
	.A2(n14), 
	.A1(n423));
   AO22CHD U6046 (.O(n4621), 
	.B2(n574), 
	.B1(\ram[252][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n423));
   AO22CHD U6047 (.O(n4622), 
	.B2(n574), 
	.B1(\ram[252][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n423));
   AO22CHD U6048 (.O(n4623), 
	.B2(n574), 
	.B1(\ram[252][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n423));
   AO22CHD U6049 (.O(n4624), 
	.B2(n574), 
	.B1(\ram[252][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n423));
   AO22CHD U6050 (.O(n4625), 
	.B2(n574), 
	.B1(\ram[252][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n423));
   AO22CHD U6051 (.O(n4626), 
	.B2(n574), 
	.B1(\ram[252][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n423));
   AO22CHD U6052 (.O(n4627), 
	.B2(n574), 
	.B1(\ram[252][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n423));
   AO22CHD U6053 (.O(n4628), 
	.B2(n574), 
	.B1(\ram[252][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n423));
   AO22CHD U6054 (.O(n4629), 
	.B2(n574), 
	.B1(\ram[252][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n423));
   AO22CHD U6055 (.O(n4630), 
	.B2(n577), 
	.B1(\ram[253][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n425));
   AO22CHD U6056 (.O(n4631), 
	.B2(n577), 
	.B1(\ram[253][1] ), 
	.A2(n9), 
	.A1(n425));
   AO22CHD U6057 (.O(n4632), 
	.B2(n577), 
	.B1(\ram[253][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n425));
   AO22CHD U6058 (.O(n4633), 
	.B2(n577), 
	.B1(\ram[253][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n425));
   AO22CHD U6059 (.O(n4634), 
	.B2(n577), 
	.B1(\ram[253][4] ), 
	.A2(n12), 
	.A1(n425));
   AO22CHD U6060 (.O(n4635), 
	.B2(n577), 
	.B1(\ram[253][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n425));
   AO22CHD U6061 (.O(n4636), 
	.B2(n577), 
	.B1(\ram[253][6] ), 
	.A2(n14), 
	.A1(n425));
   AO22CHD U6062 (.O(n4637), 
	.B2(n577), 
	.B1(\ram[253][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n425));
   AO22CHD U6063 (.O(n4638), 
	.B2(n577), 
	.B1(\ram[253][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n425));
   AO22CHD U6064 (.O(n4639), 
	.B2(n577), 
	.B1(\ram[253][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n425));
   AO22CHD U6065 (.O(n4640), 
	.B2(n577), 
	.B1(\ram[253][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n425));
   AO22CHD U6066 (.O(n4641), 
	.B2(n577), 
	.B1(\ram[253][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n425));
   AO22CHD U6067 (.O(n4642), 
	.B2(n577), 
	.B1(\ram[253][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n425));
   AO22CHD U6068 (.O(n4643), 
	.B2(n577), 
	.B1(\ram[253][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n425));
   AO22CHD U6069 (.O(n4644), 
	.B2(n577), 
	.B1(\ram[253][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n425));
   AO22CHD U6070 (.O(n4645), 
	.B2(n577), 
	.B1(\ram[253][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n425));
   AO22CHD U6071 (.O(n4646), 
	.B2(n579), 
	.B1(\ram[254][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n427));
   AO22CHD U6072 (.O(n4647), 
	.B2(n579), 
	.B1(\ram[254][1] ), 
	.A2(n9), 
	.A1(n427));
   AO22CHD U6073 (.O(n4648), 
	.B2(n579), 
	.B1(\ram[254][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n427));
   AO22CHD U6074 (.O(n4649), 
	.B2(n579), 
	.B1(\ram[254][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n427));
   AO22CHD U6075 (.O(n4650), 
	.B2(n579), 
	.B1(\ram[254][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n427));
   AO22CHD U6076 (.O(n4651), 
	.B2(n579), 
	.B1(\ram[254][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n427));
   AO22CHD U6077 (.O(n4652), 
	.B2(n579), 
	.B1(\ram[254][6] ), 
	.A2(n14), 
	.A1(n427));
   AO22CHD U6078 (.O(n4653), 
	.B2(n579), 
	.B1(\ram[254][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n427));
   AO22CHD U6079 (.O(n4654), 
	.B2(n579), 
	.B1(\ram[254][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n427));
   AO22CHD U6080 (.O(n4655), 
	.B2(n579), 
	.B1(FE_PHN2943_ram_254__9_), 
	.A2(FE_OFN72_n17), 
	.A1(n427));
   AO22CHD U6081 (.O(n4656), 
	.B2(n579), 
	.B1(\ram[254][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n427));
   AO22CHD U6082 (.O(n4657), 
	.B2(n579), 
	.B1(\ram[254][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n427));
   AO22CHD U6083 (.O(n4658), 
	.B2(n579), 
	.B1(\ram[254][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n427));
   AO22CHD U6084 (.O(n4659), 
	.B2(n579), 
	.B1(\ram[254][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n427));
   AO22CHD U6085 (.O(n4660), 
	.B2(n579), 
	.B1(\ram[254][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n427));
   AO22CHD U6086 (.O(n4661), 
	.B2(n579), 
	.B1(\ram[254][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n427));
   AO22CHD U6087 (.O(n4662), 
	.B2(n581), 
	.B1(\ram[255][0] ), 
	.A2(FE_OFN42_n6), 
	.A1(n429));
   AO22CHD U6088 (.O(n4663), 
	.B2(n581), 
	.B1(\ram[255][1] ), 
	.A2(n9), 
	.A1(n429));
   AO22CHD U6089 (.O(n4664), 
	.B2(n581), 
	.B1(\ram[255][2] ), 
	.A2(FE_OFN48_n10), 
	.A1(n429));
   AO22CHD U6090 (.O(n4665), 
	.B2(n581), 
	.B1(\ram[255][3] ), 
	.A2(FE_OFN50_n11), 
	.A1(n429));
   AO22CHD U6091 (.O(n4666), 
	.B2(n581), 
	.B1(\ram[255][4] ), 
	.A2(FE_OFN54_n12), 
	.A1(n429));
   AO22CHD U6092 (.O(n4667), 
	.B2(n581), 
	.B1(\ram[255][5] ), 
	.A2(FE_OFN56_n13), 
	.A1(n429));
   AO22CHD U6093 (.O(n4668), 
	.B2(n581), 
	.B1(\ram[255][6] ), 
	.A2(n14), 
	.A1(n429));
   AO22CHD U6094 (.O(n4669), 
	.B2(n581), 
	.B1(\ram[255][7] ), 
	.A2(FE_OFN65_n15), 
	.A1(n429));
   AO22CHD U6095 (.O(n4670), 
	.B2(n581), 
	.B1(\ram[255][8] ), 
	.A2(FE_OFN66_n16), 
	.A1(n429));
   AO22CHD U6096 (.O(n4671), 
	.B2(n581), 
	.B1(\ram[255][9] ), 
	.A2(FE_OFN72_n17), 
	.A1(n429));
   AO22CHD U6097 (.O(n4672), 
	.B2(n581), 
	.B1(\ram[255][10] ), 
	.A2(FE_OFN75_n18), 
	.A1(n429));
   AO22CHD U6098 (.O(n4673), 
	.B2(n581), 
	.B1(\ram[255][11] ), 
	.A2(FE_OFN78_n19), 
	.A1(n429));
   AO22CHD U6099 (.O(n4674), 
	.B2(n581), 
	.B1(\ram[255][12] ), 
	.A2(FE_OFN81_n20), 
	.A1(n429));
   AO22CHD U6100 (.O(n4675), 
	.B2(n581), 
	.B1(\ram[255][13] ), 
	.A2(FE_OFN84_n21), 
	.A1(n429));
   AO22CHD U6101 (.O(n4676), 
	.B2(n581), 
	.B1(\ram[255][14] ), 
	.A2(FE_OFN87_n22), 
	.A1(n429));
   AO22CHD U6102 (.O(n4677), 
	.B2(n581), 
	.B1(\ram[255][15] ), 
	.A2(FE_OFN90_n23), 
	.A1(n429));
   AO22CHD U6103 (.O(n582), 
	.B2(n8), 
	.B1(\ram[0][0] ), 
	.A2(n433), 
	.A1(n6));
   AO22CHD U6104 (.O(n583), 
	.B2(n8), 
	.B1(\ram[0][1] ), 
	.A2(n433), 
	.A1(FE_OFN46_n9));
   AO22CHD U6105 (.O(n584), 
	.B2(n8), 
	.B1(\ram[0][2] ), 
	.A2(n433), 
	.A1(FE_OFN49_n10));
   AO22CHD U6106 (.O(n585), 
	.B2(n8), 
	.B1(\ram[0][3] ), 
	.A2(n433), 
	.A1(FE_OFN52_n11));
   AO22CHD U6107 (.O(n586), 
	.B2(n8), 
	.B1(\ram[0][4] ), 
	.A2(n433), 
	.A1(FE_OFN55_n12));
   AO22CHD U6108 (.O(n587), 
	.B2(n8), 
	.B1(\ram[0][5] ), 
	.A2(n433), 
	.A1(FE_OFN58_n13));
   AO22CHD U6109 (.O(n588), 
	.B2(n8), 
	.B1(\ram[0][6] ), 
	.A2(n433), 
	.A1(FE_OFN62_n14));
   AO22CHD U6110 (.O(n589), 
	.B2(n8), 
	.B1(\ram[0][7] ), 
	.A2(n433), 
	.A1(FE_OFN63_n15));
   AO22CHD U6111 (.O(n590), 
	.B2(n8), 
	.B1(\ram[0][8] ), 
	.A2(n433), 
	.A1(FE_OFN68_n16));
   AO22CHD U6112 (.O(n591), 
	.B2(n8), 
	.B1(\ram[0][9] ), 
	.A2(n433), 
	.A1(FE_OFN70_n17));
   AO22CHD U6113 (.O(n592), 
	.B2(n8), 
	.B1(\ram[0][10] ), 
	.A2(n433), 
	.A1(FE_OFN73_n18));
   AO22CHD U6114 (.O(n593), 
	.B2(n8), 
	.B1(\ram[0][11] ), 
	.A2(n433), 
	.A1(FE_OFN76_n19));
   AO22CHD U6115 (.O(n594), 
	.B2(n8), 
	.B1(\ram[0][12] ), 
	.A2(n433), 
	.A1(FE_OFN80_n20));
   AO22CHD U6116 (.O(n595), 
	.B2(n8), 
	.B1(\ram[0][13] ), 
	.A2(n433), 
	.A1(FE_OFN85_n21));
   AO22CHD U6117 (.O(n596), 
	.B2(n8), 
	.B1(\ram[0][14] ), 
	.A2(n433), 
	.A1(n22));
   AO22CHD U6118 (.O(n597), 
	.B2(n8), 
	.B1(\ram[0][15] ), 
	.A2(n433), 
	.A1(FE_OFN91_n23));
   MUX4EHD U6119 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n571), 
	.D(\ram[255][0] ), 
	.C(\ram[253][0] ), 
	.B(\ram[254][0] ), 
	.A(\ram[252][0] ));
   MUX4EHD U6120 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n573), 
	.D(\ram[251][0] ), 
	.C(\ram[249][0] ), 
	.B(\ram[250][0] ), 
	.A(\ram[248][0] ));
   MUX4EHD U6121 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n576), 
	.D(\ram[247][0] ), 
	.C(\ram[245][0] ), 
	.B(\ram[246][0] ), 
	.A(\ram[244][0] ));
   MUX4EHD U6122 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n578), 
	.D(\ram[243][0] ), 
	.C(\ram[241][0] ), 
	.B(\ram[242][0] ), 
	.A(\ram[240][0] ));
   MUX4EHD U6123 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n580), 
	.D(n571), 
	.C(n576), 
	.B(n573), 
	.A(n578));
   MUX4EHD U6124 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4678), 
	.D(\ram[239][0] ), 
	.C(\ram[237][0] ), 
	.B(\ram[238][0] ), 
	.A(\ram[236][0] ));
   MUX4EHD U6125 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4679), 
	.D(\ram[235][0] ), 
	.C(\ram[233][0] ), 
	.B(\ram[234][0] ), 
	.A(\ram[232][0] ));
   MUX4EHD U6126 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4680), 
	.D(\ram[231][0] ), 
	.C(\ram[229][0] ), 
	.B(\ram[230][0] ), 
	.A(\ram[228][0] ));
   MUX4EHD U6127 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4681), 
	.D(\ram[227][0] ), 
	.C(\ram[225][0] ), 
	.B(\ram[226][0] ), 
	.A(\ram[224][0] ));
   MUX4EHD U6128 (.S1(n6136), 
	.S0(n7442), 
	.O(n4682), 
	.D(n4678), 
	.C(n4680), 
	.B(n4679), 
	.A(n4681));
   MUX4EHD U6129 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4683), 
	.D(\ram[223][0] ), 
	.C(\ram[221][0] ), 
	.B(\ram[222][0] ), 
	.A(\ram[220][0] ));
   MUX4EHD U6130 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4684), 
	.D(\ram[219][0] ), 
	.C(\ram[217][0] ), 
	.B(\ram[218][0] ), 
	.A(\ram[216][0] ));
   MUX4EHD U6131 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4685), 
	.D(\ram[215][0] ), 
	.C(\ram[213][0] ), 
	.B(\ram[214][0] ), 
	.A(\ram[212][0] ));
   MUX4EHD U6132 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4686), 
	.D(\ram[211][0] ), 
	.C(\ram[209][0] ), 
	.B(\ram[210][0] ), 
	.A(\ram[208][0] ));
   MUX4EHD U6133 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4687), 
	.D(n4683), 
	.C(n4685), 
	.B(n4684), 
	.A(n4686));
   MUX4EHD U6134 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4688), 
	.D(\ram[207][0] ), 
	.C(\ram[205][0] ), 
	.B(\ram[206][0] ), 
	.A(\ram[204][0] ));
   MUX4EHD U6135 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4689), 
	.D(\ram[203][0] ), 
	.C(\ram[201][0] ), 
	.B(\ram[202][0] ), 
	.A(\ram[200][0] ));
   MUX4EHD U6136 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4690), 
	.D(\ram[199][0] ), 
	.C(\ram[197][0] ), 
	.B(\ram[198][0] ), 
	.A(\ram[196][0] ));
   MUX4EHD U6137 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4691), 
	.D(\ram[195][0] ), 
	.C(\ram[193][0] ), 
	.B(\ram[194][0] ), 
	.A(\ram[192][0] ));
   MUX4EHD U6138 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4692), 
	.D(n4688), 
	.C(n4690), 
	.B(n4689), 
	.A(n4691));
   MUX4EHD U6139 (.S1(n6038), 
	.S0(n7444), 
	.O(n4693), 
	.D(n580), 
	.C(n4687), 
	.B(n4682), 
	.A(n4692));
   MUX4EHD U6140 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4694), 
	.D(\ram[191][0] ), 
	.C(\ram[189][0] ), 
	.B(\ram[190][0] ), 
	.A(\ram[188][0] ));
   MUX4EHD U6141 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4695), 
	.D(\ram[187][0] ), 
	.C(\ram[185][0] ), 
	.B(\ram[186][0] ), 
	.A(\ram[184][0] ));
   MUX4EHD U6142 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4696), 
	.D(\ram[183][0] ), 
	.C(\ram[181][0] ), 
	.B(\ram[182][0] ), 
	.A(\ram[180][0] ));
   MUX4EHD U6143 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4697), 
	.D(\ram[179][0] ), 
	.C(\ram[177][0] ), 
	.B(\ram[178][0] ), 
	.A(\ram[176][0] ));
   MUX4EHD U6144 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4698), 
	.D(n4694), 
	.C(n4696), 
	.B(n4695), 
	.A(n4697));
   MUX4EHD U6145 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4699), 
	.D(\ram[175][0] ), 
	.C(\ram[173][0] ), 
	.B(\ram[174][0] ), 
	.A(\ram[172][0] ));
   MUX4EHD U6146 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4700), 
	.D(\ram[171][0] ), 
	.C(\ram[169][0] ), 
	.B(\ram[170][0] ), 
	.A(\ram[168][0] ));
   MUX4EHD U6147 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4701), 
	.D(\ram[167][0] ), 
	.C(\ram[165][0] ), 
	.B(\ram[166][0] ), 
	.A(\ram[164][0] ));
   MUX4EHD U6148 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4702), 
	.D(\ram[163][0] ), 
	.C(\ram[161][0] ), 
	.B(\ram[162][0] ), 
	.A(\ram[160][0] ));
   MUX4EHD U6149 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4703), 
	.D(n4699), 
	.C(n4701), 
	.B(n4700), 
	.A(n4702));
   MUX4EHD U6150 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4704), 
	.D(\ram[159][0] ), 
	.C(\ram[157][0] ), 
	.B(\ram[158][0] ), 
	.A(\ram[156][0] ));
   MUX4EHD U6151 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4705), 
	.D(\ram[155][0] ), 
	.C(\ram[153][0] ), 
	.B(\ram[154][0] ), 
	.A(\ram[152][0] ));
   MUX4EHD U6152 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4706), 
	.D(\ram[151][0] ), 
	.C(\ram[149][0] ), 
	.B(\ram[150][0] ), 
	.A(\ram[148][0] ));
   MUX4EHD U6153 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4707), 
	.D(\ram[147][0] ), 
	.C(\ram[145][0] ), 
	.B(\ram[146][0] ), 
	.A(\ram[144][0] ));
   MUX4EHD U6154 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4708), 
	.D(n4704), 
	.C(n4706), 
	.B(n4705), 
	.A(n4707));
   MUX4EHD U6155 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4709), 
	.D(\ram[143][0] ), 
	.C(\ram[141][0] ), 
	.B(\ram[142][0] ), 
	.A(\ram[140][0] ));
   MUX4EHD U6156 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4710), 
	.D(\ram[139][0] ), 
	.C(\ram[137][0] ), 
	.B(\ram[138][0] ), 
	.A(\ram[136][0] ));
   MUX4EHD U6157 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4711), 
	.D(\ram[135][0] ), 
	.C(\ram[133][0] ), 
	.B(\ram[134][0] ), 
	.A(\ram[132][0] ));
   MUX4EHD U6158 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4712), 
	.D(\ram[131][0] ), 
	.C(\ram[129][0] ), 
	.B(\ram[130][0] ), 
	.A(\ram[128][0] ));
   MUX4EHD U6159 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4713), 
	.D(n4709), 
	.C(n4711), 
	.B(n4710), 
	.A(n4712));
   MUX4EHD U6160 (.S1(n6038), 
	.S0(n7444), 
	.O(n4714), 
	.D(n4698), 
	.C(n4708), 
	.B(n4703), 
	.A(n4713));
   MUX4EHD U6161 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4715), 
	.D(\ram[127][0] ), 
	.C(\ram[125][0] ), 
	.B(\ram[126][0] ), 
	.A(\ram[124][0] ));
   MUX4EHD U6162 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4716), 
	.D(\ram[123][0] ), 
	.C(\ram[121][0] ), 
	.B(\ram[122][0] ), 
	.A(\ram[120][0] ));
   MUX4EHD U6163 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4717), 
	.D(\ram[119][0] ), 
	.C(\ram[117][0] ), 
	.B(\ram[118][0] ), 
	.A(\ram[116][0] ));
   MUX4EHD U6164 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4718), 
	.D(\ram[115][0] ), 
	.C(\ram[113][0] ), 
	.B(\ram[114][0] ), 
	.A(\ram[112][0] ));
   MUX4EHD U6165 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4719), 
	.D(n4715), 
	.C(n4717), 
	.B(n4716), 
	.A(n4718));
   MUX4EHD U6166 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4720), 
	.D(\ram[111][0] ), 
	.C(\ram[109][0] ), 
	.B(\ram[110][0] ), 
	.A(\ram[108][0] ));
   MUX4EHD U6167 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4721), 
	.D(\ram[107][0] ), 
	.C(\ram[105][0] ), 
	.B(\ram[106][0] ), 
	.A(\ram[104][0] ));
   MUX4EHD U6168 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4722), 
	.D(\ram[103][0] ), 
	.C(\ram[101][0] ), 
	.B(\ram[102][0] ), 
	.A(\ram[100][0] ));
   MUX4EHD U6169 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4723), 
	.D(\ram[99][0] ), 
	.C(\ram[97][0] ), 
	.B(\ram[98][0] ), 
	.A(\ram[96][0] ));
   MUX4EHD U6170 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4724), 
	.D(n4720), 
	.C(n4722), 
	.B(n4721), 
	.A(n4723));
   MUX4EHD U6171 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4725), 
	.D(\ram[95][0] ), 
	.C(\ram[93][0] ), 
	.B(\ram[94][0] ), 
	.A(\ram[92][0] ));
   MUX4EHD U6172 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4726), 
	.D(\ram[91][0] ), 
	.C(\ram[89][0] ), 
	.B(\ram[90][0] ), 
	.A(\ram[88][0] ));
   MUX4EHD U6173 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4727), 
	.D(\ram[87][0] ), 
	.C(\ram[85][0] ), 
	.B(\ram[86][0] ), 
	.A(\ram[84][0] ));
   MUX4EHD U6174 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4728), 
	.D(\ram[83][0] ), 
	.C(\ram[81][0] ), 
	.B(\ram[82][0] ), 
	.A(\ram[80][0] ));
   MUX4EHD U6175 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4729), 
	.D(n4725), 
	.C(n4727), 
	.B(n4726), 
	.A(n4728));
   MUX4EHD U6176 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4730), 
	.D(\ram[79][0] ), 
	.C(\ram[77][0] ), 
	.B(\ram[78][0] ), 
	.A(\ram[76][0] ));
   MUX4EHD U6177 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4731), 
	.D(\ram[75][0] ), 
	.C(\ram[73][0] ), 
	.B(\ram[74][0] ), 
	.A(\ram[72][0] ));
   MUX4EHD U6178 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4732), 
	.D(\ram[71][0] ), 
	.C(\ram[69][0] ), 
	.B(\ram[70][0] ), 
	.A(\ram[68][0] ));
   MUX4EHD U6179 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4733), 
	.D(\ram[67][0] ), 
	.C(\ram[65][0] ), 
	.B(\ram[66][0] ), 
	.A(\ram[64][0] ));
   MUX4EHD U6180 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4734), 
	.D(n4730), 
	.C(n4732), 
	.B(n4731), 
	.A(n4733));
   MUX4EHD U6181 (.S1(n6038), 
	.S0(n7444), 
	.O(n4735), 
	.D(n4719), 
	.C(n4729), 
	.B(n4724), 
	.A(n4734));
   MUX4EHD U6182 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4736), 
	.D(\ram[63][0] ), 
	.C(\ram[61][0] ), 
	.B(\ram[62][0] ), 
	.A(\ram[60][0] ));
   MUX4EHD U6183 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4737), 
	.D(\ram[59][0] ), 
	.C(\ram[57][0] ), 
	.B(\ram[58][0] ), 
	.A(\ram[56][0] ));
   MUX4EHD U6184 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4738), 
	.D(\ram[55][0] ), 
	.C(\ram[53][0] ), 
	.B(\ram[54][0] ), 
	.A(\ram[52][0] ));
   MUX4EHD U6185 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4739), 
	.D(\ram[51][0] ), 
	.C(\ram[49][0] ), 
	.B(\ram[50][0] ), 
	.A(\ram[48][0] ));
   MUX4EHD U6186 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4740), 
	.D(n4736), 
	.C(n4738), 
	.B(n4737), 
	.A(n4739));
   MUX4EHD U6187 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4741), 
	.D(\ram[47][0] ), 
	.C(\ram[45][0] ), 
	.B(\ram[46][0] ), 
	.A(\ram[44][0] ));
   MUX4EHD U6188 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4742), 
	.D(\ram[43][0] ), 
	.C(\ram[41][0] ), 
	.B(\ram[42][0] ), 
	.A(\ram[40][0] ));
   MUX4EHD U6189 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4743), 
	.D(\ram[39][0] ), 
	.C(\ram[37][0] ), 
	.B(\ram[38][0] ), 
	.A(\ram[36][0] ));
   MUX4EHD U6190 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4744), 
	.D(\ram[35][0] ), 
	.C(\ram[33][0] ), 
	.B(\ram[34][0] ), 
	.A(\ram[32][0] ));
   MUX4EHD U6191 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4745), 
	.D(n4741), 
	.C(n4743), 
	.B(n4742), 
	.A(n4744));
   MUX4EHD U6192 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4746), 
	.D(\ram[31][0] ), 
	.C(\ram[29][0] ), 
	.B(\ram[30][0] ), 
	.A(\ram[28][0] ));
   MUX4EHD U6193 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4747), 
	.D(\ram[27][0] ), 
	.C(\ram[25][0] ), 
	.B(\ram[26][0] ), 
	.A(\ram[24][0] ));
   MUX4EHD U6194 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4748), 
	.D(\ram[23][0] ), 
	.C(\ram[21][0] ), 
	.B(\ram[22][0] ), 
	.A(\ram[20][0] ));
   MUX4EHD U6195 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4749), 
	.D(\ram[19][0] ), 
	.C(\ram[17][0] ), 
	.B(\ram[18][0] ), 
	.A(\ram[16][0] ));
   MUX4EHD U6196 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4750), 
	.D(n4746), 
	.C(n4748), 
	.B(n4747), 
	.A(n4749));
   MUX4EHD U6197 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4751), 
	.D(\ram[15][0] ), 
	.C(\ram[13][0] ), 
	.B(\ram[14][0] ), 
	.A(\ram[12][0] ));
   MUX4EHD U6198 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4752), 
	.D(\ram[11][0] ), 
	.C(\ram[9][0] ), 
	.B(\ram[10][0] ), 
	.A(\ram[8][0] ));
   MUX4EHD U6199 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4753), 
	.D(\ram[7][0] ), 
	.C(\ram[5][0] ), 
	.B(\ram[6][0] ), 
	.A(\ram[4][0] ));
   MUX4EHD U6200 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4754), 
	.D(\ram[3][0] ), 
	.C(\ram[1][0] ), 
	.B(\ram[2][0] ), 
	.A(\ram[0][0] ));
   MUX4EHD U6201 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4755), 
	.D(n4751), 
	.C(n4753), 
	.B(n4752), 
	.A(n4754));
   MUX4EHD U6202 (.S1(n6038), 
	.S0(n7444), 
	.O(n4756), 
	.D(n4740), 
	.C(n4750), 
	.B(n4745), 
	.A(n4755));
   MUX4EHD U6203 (.S1(n6469), 
	.S0(n6470), 
	.O(N4141), 
	.D(n4693), 
	.C(n4735), 
	.B(n4714), 
	.A(n4756));
   MUX4EHD U6204 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4757), 
	.D(\ram[255][1] ), 
	.C(\ram[253][1] ), 
	.B(\ram[254][1] ), 
	.A(\ram[252][1] ));
   MUX4EHD U6205 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4758), 
	.D(\ram[251][1] ), 
	.C(\ram[249][1] ), 
	.B(\ram[250][1] ), 
	.A(\ram[248][1] ));
   MUX4EHD U6206 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4759), 
	.D(\ram[247][1] ), 
	.C(\ram[245][1] ), 
	.B(\ram[246][1] ), 
	.A(\ram[244][1] ));
   MUX4EHD U6207 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4760), 
	.D(\ram[243][1] ), 
	.C(\ram[241][1] ), 
	.B(\ram[242][1] ), 
	.A(\ram[240][1] ));
   MUX4EHD U6208 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4761), 
	.D(n4757), 
	.C(n4759), 
	.B(n4758), 
	.A(n4760));
   MUX4EHD U6209 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4762), 
	.D(\ram[239][1] ), 
	.C(\ram[237][1] ), 
	.B(\ram[238][1] ), 
	.A(\ram[236][1] ));
   MUX4EHD U6210 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4763), 
	.D(\ram[235][1] ), 
	.C(\ram[233][1] ), 
	.B(\ram[234][1] ), 
	.A(\ram[232][1] ));
   MUX4EHD U6211 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4764), 
	.D(\ram[231][1] ), 
	.C(\ram[229][1] ), 
	.B(\ram[230][1] ), 
	.A(\ram[228][1] ));
   MUX4EHD U6212 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4765), 
	.D(\ram[227][1] ), 
	.C(\ram[225][1] ), 
	.B(\ram[226][1] ), 
	.A(\ram[224][1] ));
   MUX4EHD U6213 (.S1(n6136), 
	.S0(n7442), 
	.O(n4766), 
	.D(n4762), 
	.C(n4764), 
	.B(n4763), 
	.A(n4765));
   MUX4EHD U6214 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4767), 
	.D(\ram[223][1] ), 
	.C(\ram[221][1] ), 
	.B(\ram[222][1] ), 
	.A(\ram[220][1] ));
   MUX4EHD U6215 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4768), 
	.D(\ram[219][1] ), 
	.C(\ram[217][1] ), 
	.B(\ram[218][1] ), 
	.A(\ram[216][1] ));
   MUX4EHD U6216 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4769), 
	.D(\ram[215][1] ), 
	.C(\ram[213][1] ), 
	.B(\ram[214][1] ), 
	.A(\ram[212][1] ));
   MUX4EHD U6217 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4770), 
	.D(\ram[211][1] ), 
	.C(\ram[209][1] ), 
	.B(\ram[210][1] ), 
	.A(\ram[208][1] ));
   MUX4EHD U6218 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4771), 
	.D(n4767), 
	.C(n4769), 
	.B(n4768), 
	.A(n4770));
   MUX4EHD U6219 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4772), 
	.D(\ram[207][1] ), 
	.C(\ram[205][1] ), 
	.B(\ram[206][1] ), 
	.A(\ram[204][1] ));
   MUX4EHD U6220 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4773), 
	.D(\ram[203][1] ), 
	.C(\ram[201][1] ), 
	.B(\ram[202][1] ), 
	.A(\ram[200][1] ));
   MUX4EHD U6221 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4774), 
	.D(\ram[199][1] ), 
	.C(\ram[197][1] ), 
	.B(\ram[198][1] ), 
	.A(\ram[196][1] ));
   MUX4EHD U6222 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4775), 
	.D(\ram[195][1] ), 
	.C(\ram[193][1] ), 
	.B(\ram[194][1] ), 
	.A(\ram[192][1] ));
   MUX4EHD U6223 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4776), 
	.D(n4772), 
	.C(n4774), 
	.B(n4773), 
	.A(n4775));
   MUX4EHD U6224 (.S1(n6038), 
	.S0(n7444), 
	.O(n4777), 
	.D(n4761), 
	.C(n4771), 
	.B(n4766), 
	.A(n4776));
   MUX4EHD U6225 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4778), 
	.D(\ram[191][1] ), 
	.C(\ram[189][1] ), 
	.B(\ram[190][1] ), 
	.A(\ram[188][1] ));
   MUX4EHD U6226 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4779), 
	.D(\ram[187][1] ), 
	.C(\ram[185][1] ), 
	.B(\ram[186][1] ), 
	.A(\ram[184][1] ));
   MUX4EHD U6227 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4780), 
	.D(\ram[183][1] ), 
	.C(\ram[181][1] ), 
	.B(\ram[182][1] ), 
	.A(\ram[180][1] ));
   MUX4EHD U6228 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4781), 
	.D(\ram[179][1] ), 
	.C(\ram[177][1] ), 
	.B(\ram[178][1] ), 
	.A(\ram[176][1] ));
   MUX4EHD U6229 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4782), 
	.D(n4778), 
	.C(n4780), 
	.B(n4779), 
	.A(n4781));
   MUX4EHD U6230 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4783), 
	.D(\ram[175][1] ), 
	.C(\ram[173][1] ), 
	.B(\ram[174][1] ), 
	.A(\ram[172][1] ));
   MUX4EHD U6231 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4784), 
	.D(\ram[171][1] ), 
	.C(\ram[169][1] ), 
	.B(\ram[170][1] ), 
	.A(\ram[168][1] ));
   MUX4EHD U6232 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4785), 
	.D(\ram[167][1] ), 
	.C(\ram[165][1] ), 
	.B(\ram[166][1] ), 
	.A(\ram[164][1] ));
   MUX4EHD U6233 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4786), 
	.D(\ram[163][1] ), 
	.C(\ram[161][1] ), 
	.B(\ram[162][1] ), 
	.A(\ram[160][1] ));
   MUX4EHD U6234 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4787), 
	.D(n4783), 
	.C(n4785), 
	.B(n4784), 
	.A(n4786));
   MUX4EHD U6235 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4788), 
	.D(\ram[159][1] ), 
	.C(\ram[157][1] ), 
	.B(\ram[158][1] ), 
	.A(\ram[156][1] ));
   MUX4EHD U6236 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4789), 
	.D(\ram[155][1] ), 
	.C(\ram[153][1] ), 
	.B(\ram[154][1] ), 
	.A(\ram[152][1] ));
   MUX4EHD U6237 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4790), 
	.D(\ram[151][1] ), 
	.C(\ram[149][1] ), 
	.B(\ram[150][1] ), 
	.A(\ram[148][1] ));
   MUX4EHD U6238 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4791), 
	.D(\ram[147][1] ), 
	.C(\ram[145][1] ), 
	.B(\ram[146][1] ), 
	.A(\ram[144][1] ));
   MUX4EHD U6239 (.S1(n6136), 
	.S0(n7442), 
	.O(n4792), 
	.D(n4788), 
	.C(n4790), 
	.B(n4789), 
	.A(n4791));
   MUX4EHD U6240 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4793), 
	.D(\ram[143][1] ), 
	.C(\ram[141][1] ), 
	.B(\ram[142][1] ), 
	.A(\ram[140][1] ));
   MUX4EHD U6241 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4794), 
	.D(\ram[139][1] ), 
	.C(\ram[137][1] ), 
	.B(\ram[138][1] ), 
	.A(\ram[136][1] ));
   MUX4EHD U6242 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4795), 
	.D(\ram[135][1] ), 
	.C(\ram[133][1] ), 
	.B(\ram[134][1] ), 
	.A(\ram[132][1] ));
   MUX4EHD U6243 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4796), 
	.D(\ram[131][1] ), 
	.C(\ram[129][1] ), 
	.B(\ram[130][1] ), 
	.A(\ram[128][1] ));
   MUX4EHD U6244 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4797), 
	.D(n4793), 
	.C(n4795), 
	.B(n4794), 
	.A(n4796));
   MUX4EHD U6245 (.S1(n6038), 
	.S0(n7444), 
	.O(n4798), 
	.D(n4782), 
	.C(n4792), 
	.B(n4787), 
	.A(n4797));
   MUX4EHD U6246 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4799), 
	.D(\ram[127][1] ), 
	.C(\ram[125][1] ), 
	.B(\ram[126][1] ), 
	.A(\ram[124][1] ));
   MUX4EHD U6247 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4800), 
	.D(\ram[123][1] ), 
	.C(\ram[121][1] ), 
	.B(\ram[122][1] ), 
	.A(\ram[120][1] ));
   MUX4EHD U6248 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4801), 
	.D(\ram[119][1] ), 
	.C(\ram[117][1] ), 
	.B(\ram[118][1] ), 
	.A(\ram[116][1] ));
   MUX4EHD U6249 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4802), 
	.D(\ram[115][1] ), 
	.C(\ram[113][1] ), 
	.B(\ram[114][1] ), 
	.A(\ram[112][1] ));
   MUX4EHD U6250 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4803), 
	.D(n4799), 
	.C(n4801), 
	.B(n4800), 
	.A(n4802));
   MUX4EHD U6251 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4804), 
	.D(\ram[111][1] ), 
	.C(\ram[109][1] ), 
	.B(\ram[110][1] ), 
	.A(\ram[108][1] ));
   MUX4EHD U6252 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4805), 
	.D(\ram[107][1] ), 
	.C(\ram[105][1] ), 
	.B(\ram[106][1] ), 
	.A(\ram[104][1] ));
   MUX4EHD U6253 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4806), 
	.D(\ram[103][1] ), 
	.C(\ram[101][1] ), 
	.B(\ram[102][1] ), 
	.A(\ram[100][1] ));
   MUX4EHD U6254 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4807), 
	.D(\ram[99][1] ), 
	.C(\ram[97][1] ), 
	.B(\ram[98][1] ), 
	.A(\ram[96][1] ));
   MUX4EHD U6255 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4808), 
	.D(n4804), 
	.C(n4806), 
	.B(n4805), 
	.A(n4807));
   MUX4EHD U6256 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4809), 
	.D(\ram[95][1] ), 
	.C(\ram[93][1] ), 
	.B(\ram[94][1] ), 
	.A(\ram[92][1] ));
   MUX4EHD U6257 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4810), 
	.D(\ram[91][1] ), 
	.C(\ram[89][1] ), 
	.B(\ram[90][1] ), 
	.A(\ram[88][1] ));
   MUX4EHD U6258 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4811), 
	.D(\ram[87][1] ), 
	.C(\ram[85][1] ), 
	.B(\ram[86][1] ), 
	.A(\ram[84][1] ));
   MUX4EHD U6259 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4812), 
	.D(\ram[83][1] ), 
	.C(\ram[81][1] ), 
	.B(\ram[82][1] ), 
	.A(\ram[80][1] ));
   MUX4EHD U6260 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4813), 
	.D(n4809), 
	.C(n4811), 
	.B(n4810), 
	.A(n4812));
   MUX4EHD U6261 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4814), 
	.D(\ram[79][1] ), 
	.C(\ram[77][1] ), 
	.B(\ram[78][1] ), 
	.A(\ram[76][1] ));
   MUX4EHD U6262 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4815), 
	.D(\ram[75][1] ), 
	.C(\ram[73][1] ), 
	.B(\ram[74][1] ), 
	.A(\ram[72][1] ));
   MUX4EHD U6263 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4816), 
	.D(\ram[71][1] ), 
	.C(\ram[69][1] ), 
	.B(\ram[70][1] ), 
	.A(\ram[68][1] ));
   MUX4EHD U6264 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4817), 
	.D(\ram[67][1] ), 
	.C(\ram[65][1] ), 
	.B(\ram[66][1] ), 
	.A(\ram[64][1] ));
   MUX4EHD U6265 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4818), 
	.D(n4814), 
	.C(n4816), 
	.B(n4815), 
	.A(n4817));
   MUX4EHD U6266 (.S1(n6038), 
	.S0(n7444), 
	.O(n4819), 
	.D(n4803), 
	.C(n4813), 
	.B(n4808), 
	.A(n4818));
   MUX4EHD U6267 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4820), 
	.D(\ram[63][1] ), 
	.C(\ram[61][1] ), 
	.B(\ram[62][1] ), 
	.A(\ram[60][1] ));
   MUX4EHD U6268 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4821), 
	.D(\ram[59][1] ), 
	.C(\ram[57][1] ), 
	.B(\ram[58][1] ), 
	.A(\ram[56][1] ));
   MUX4EHD U6269 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4822), 
	.D(\ram[55][1] ), 
	.C(\ram[53][1] ), 
	.B(\ram[54][1] ), 
	.A(\ram[52][1] ));
   MUX4EHD U6270 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4823), 
	.D(\ram[51][1] ), 
	.C(\ram[49][1] ), 
	.B(\ram[50][1] ), 
	.A(\ram[48][1] ));
   MUX4EHD U6271 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4824), 
	.D(n4820), 
	.C(n4822), 
	.B(n4821), 
	.A(n4823));
   MUX4EHD U6272 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4825), 
	.D(\ram[47][1] ), 
	.C(\ram[45][1] ), 
	.B(\ram[46][1] ), 
	.A(\ram[44][1] ));
   MUX4EHD U6273 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4826), 
	.D(\ram[43][1] ), 
	.C(\ram[41][1] ), 
	.B(\ram[42][1] ), 
	.A(\ram[40][1] ));
   MUX4EHD U6274 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4827), 
	.D(\ram[39][1] ), 
	.C(\ram[37][1] ), 
	.B(\ram[38][1] ), 
	.A(\ram[36][1] ));
   MUX4EHD U6275 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4828), 
	.D(\ram[35][1] ), 
	.C(\ram[33][1] ), 
	.B(\ram[34][1] ), 
	.A(\ram[32][1] ));
   MUX4EHD U6276 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4829), 
	.D(n4825), 
	.C(n4827), 
	.B(n4826), 
	.A(n4828));
   MUX4EHD U6277 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4830), 
	.D(\ram[31][1] ), 
	.C(\ram[29][1] ), 
	.B(\ram[30][1] ), 
	.A(\ram[28][1] ));
   MUX4EHD U6278 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4831), 
	.D(\ram[27][1] ), 
	.C(\ram[25][1] ), 
	.B(\ram[26][1] ), 
	.A(\ram[24][1] ));
   MUX4EHD U6279 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4832), 
	.D(\ram[23][1] ), 
	.C(\ram[21][1] ), 
	.B(\ram[22][1] ), 
	.A(\ram[20][1] ));
   MUX4EHD U6280 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4833), 
	.D(\ram[19][1] ), 
	.C(\ram[17][1] ), 
	.B(\ram[18][1] ), 
	.A(\ram[16][1] ));
   MUX4EHD U6281 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4834), 
	.D(n4830), 
	.C(n4832), 
	.B(n4831), 
	.A(n4833));
   MUX4EHD U6282 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n4835), 
	.D(\ram[15][1] ), 
	.C(\ram[13][1] ), 
	.B(\ram[14][1] ), 
	.A(\ram[12][1] ));
   MUX4EHD U6283 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n4836), 
	.D(\ram[11][1] ), 
	.C(\ram[9][1] ), 
	.B(\ram[10][1] ), 
	.A(\ram[8][1] ));
   MUX4EHD U6284 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4837), 
	.D(\ram[7][1] ), 
	.C(\ram[5][1] ), 
	.B(\ram[6][1] ), 
	.A(\ram[4][1] ));
   MUX4EHD U6285 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n4838), 
	.D(\ram[3][1] ), 
	.C(\ram[1][1] ), 
	.B(\ram[2][1] ), 
	.A(\ram[0][1] ));
   MUX4EHD U6286 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4839), 
	.D(n4835), 
	.C(n4837), 
	.B(n4836), 
	.A(n4838));
   MUX4EHD U6287 (.S1(n6038), 
	.S0(n7444), 
	.O(n4840), 
	.D(n4824), 
	.C(n4834), 
	.B(n4829), 
	.A(n4839));
   MUX4EHD U6288 (.S1(n6469), 
	.S0(n6470), 
	.O(N4140), 
	.D(n4777), 
	.C(n4819), 
	.B(n4798), 
	.A(n4840));
   MUX4EHD U6289 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4841), 
	.D(\ram[255][2] ), 
	.C(\ram[253][2] ), 
	.B(\ram[254][2] ), 
	.A(\ram[252][2] ));
   MUX4EHD U6290 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4842), 
	.D(\ram[251][2] ), 
	.C(\ram[249][2] ), 
	.B(\ram[250][2] ), 
	.A(\ram[248][2] ));
   MUX4EHD U6291 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4843), 
	.D(\ram[247][2] ), 
	.C(\ram[245][2] ), 
	.B(\ram[246][2] ), 
	.A(\ram[244][2] ));
   MUX4EHD U6292 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4844), 
	.D(\ram[243][2] ), 
	.C(\ram[241][2] ), 
	.B(\ram[242][2] ), 
	.A(\ram[240][2] ));
   MUX4EHD U6293 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4845), 
	.D(n4841), 
	.C(n4843), 
	.B(n4842), 
	.A(n4844));
   MUX4EHD U6294 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4846), 
	.D(\ram[239][2] ), 
	.C(\ram[237][2] ), 
	.B(\ram[238][2] ), 
	.A(\ram[236][2] ));
   MUX4EHD U6295 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4847), 
	.D(\ram[235][2] ), 
	.C(\ram[233][2] ), 
	.B(\ram[234][2] ), 
	.A(\ram[232][2] ));
   MUX4EHD U6296 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4848), 
	.D(\ram[231][2] ), 
	.C(\ram[229][2] ), 
	.B(\ram[230][2] ), 
	.A(\ram[228][2] ));
   MUX4EHD U6297 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4849), 
	.D(\ram[227][2] ), 
	.C(\ram[225][2] ), 
	.B(\ram[226][2] ), 
	.A(\ram[224][2] ));
   MUX4EHD U6298 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4850), 
	.D(n4846), 
	.C(n4848), 
	.B(n4847), 
	.A(n4849));
   MUX4EHD U6299 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4851), 
	.D(\ram[223][2] ), 
	.C(\ram[221][2] ), 
	.B(\ram[222][2] ), 
	.A(\ram[220][2] ));
   MUX4EHD U6300 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4852), 
	.D(\ram[219][2] ), 
	.C(\ram[217][2] ), 
	.B(\ram[218][2] ), 
	.A(\ram[216][2] ));
   MUX4EHD U6301 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4853), 
	.D(\ram[215][2] ), 
	.C(\ram[213][2] ), 
	.B(\ram[214][2] ), 
	.A(\ram[212][2] ));
   MUX4EHD U6302 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4854), 
	.D(\ram[211][2] ), 
	.C(\ram[209][2] ), 
	.B(\ram[210][2] ), 
	.A(\ram[208][2] ));
   MUX4EHD U6303 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4855), 
	.D(n4851), 
	.C(n4853), 
	.B(n4852), 
	.A(n4854));
   MUX4EHD U6304 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4856), 
	.D(\ram[207][2] ), 
	.C(\ram[205][2] ), 
	.B(\ram[206][2] ), 
	.A(\ram[204][2] ));
   MUX4EHD U6305 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4857), 
	.D(\ram[203][2] ), 
	.C(\ram[201][2] ), 
	.B(\ram[202][2] ), 
	.A(\ram[200][2] ));
   MUX4EHD U6306 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4858), 
	.D(\ram[199][2] ), 
	.C(\ram[197][2] ), 
	.B(\ram[198][2] ), 
	.A(\ram[196][2] ));
   MUX4EHD U6307 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4859), 
	.D(\ram[195][2] ), 
	.C(\ram[193][2] ), 
	.B(\ram[194][2] ), 
	.A(\ram[192][2] ));
   MUX4EHD U6308 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4860), 
	.D(n4856), 
	.C(n4858), 
	.B(n4857), 
	.A(n4859));
   MUX4EHD U6309 (.S1(n6038), 
	.S0(n7444), 
	.O(n4861), 
	.D(n4845), 
	.C(n4855), 
	.B(n4850), 
	.A(n4860));
   MUX4EHD U6310 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4862), 
	.D(\ram[191][2] ), 
	.C(\ram[189][2] ), 
	.B(\ram[190][2] ), 
	.A(\ram[188][2] ));
   MUX4EHD U6311 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4863), 
	.D(\ram[187][2] ), 
	.C(\ram[185][2] ), 
	.B(\ram[186][2] ), 
	.A(\ram[184][2] ));
   MUX4EHD U6312 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4864), 
	.D(\ram[183][2] ), 
	.C(\ram[181][2] ), 
	.B(\ram[182][2] ), 
	.A(\ram[180][2] ));
   MUX4EHD U6313 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4865), 
	.D(\ram[179][2] ), 
	.C(\ram[177][2] ), 
	.B(\ram[178][2] ), 
	.A(\ram[176][2] ));
   MUX4EHD U6314 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4866), 
	.D(n4862), 
	.C(n4864), 
	.B(n4863), 
	.A(n4865));
   MUX4EHD U6315 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4867), 
	.D(\ram[175][2] ), 
	.C(\ram[173][2] ), 
	.B(\ram[174][2] ), 
	.A(\ram[172][2] ));
   MUX4EHD U6316 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4868), 
	.D(\ram[171][2] ), 
	.C(\ram[169][2] ), 
	.B(\ram[170][2] ), 
	.A(\ram[168][2] ));
   MUX4EHD U6317 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4869), 
	.D(\ram[167][2] ), 
	.C(\ram[165][2] ), 
	.B(\ram[166][2] ), 
	.A(\ram[164][2] ));
   MUX4EHD U6318 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4870), 
	.D(\ram[163][2] ), 
	.C(\ram[161][2] ), 
	.B(\ram[162][2] ), 
	.A(\ram[160][2] ));
   MUX4EHD U6319 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4871), 
	.D(n4867), 
	.C(n4869), 
	.B(n4868), 
	.A(n4870));
   MUX4EHD U6320 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4872), 
	.D(\ram[159][2] ), 
	.C(\ram[157][2] ), 
	.B(\ram[158][2] ), 
	.A(\ram[156][2] ));
   MUX4EHD U6321 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4873), 
	.D(\ram[155][2] ), 
	.C(\ram[153][2] ), 
	.B(\ram[154][2] ), 
	.A(\ram[152][2] ));
   MUX4EHD U6322 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n4874), 
	.D(\ram[151][2] ), 
	.C(\ram[149][2] ), 
	.B(\ram[150][2] ), 
	.A(\ram[148][2] ));
   MUX4EHD U6323 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4875), 
	.D(\ram[147][2] ), 
	.C(\ram[145][2] ), 
	.B(\ram[146][2] ), 
	.A(\ram[144][2] ));
   MUX4EHD U6324 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4876), 
	.D(n4872), 
	.C(n4874), 
	.B(n4873), 
	.A(n4875));
   MUX4EHD U6325 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4877), 
	.D(\ram[143][2] ), 
	.C(\ram[141][2] ), 
	.B(\ram[142][2] ), 
	.A(\ram[140][2] ));
   MUX4EHD U6326 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4878), 
	.D(\ram[139][2] ), 
	.C(\ram[137][2] ), 
	.B(\ram[138][2] ), 
	.A(\ram[136][2] ));
   MUX4EHD U6327 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4879), 
	.D(\ram[135][2] ), 
	.C(\ram[133][2] ), 
	.B(\ram[134][2] ), 
	.A(\ram[132][2] ));
   MUX4EHD U6328 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4880), 
	.D(\ram[131][2] ), 
	.C(\ram[129][2] ), 
	.B(\ram[130][2] ), 
	.A(\ram[128][2] ));
   MUX4EHD U6329 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4881), 
	.D(n4877), 
	.C(n4879), 
	.B(n4878), 
	.A(n4880));
   MUX4EHD U6330 (.S1(n6038), 
	.S0(n7444), 
	.O(n4882), 
	.D(n4866), 
	.C(n4876), 
	.B(n4871), 
	.A(n4881));
   MUX4EHD U6331 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4883), 
	.D(\ram[127][2] ), 
	.C(\ram[125][2] ), 
	.B(\ram[126][2] ), 
	.A(\ram[124][2] ));
   MUX4EHD U6332 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4884), 
	.D(\ram[123][2] ), 
	.C(\ram[121][2] ), 
	.B(\ram[122][2] ), 
	.A(\ram[120][2] ));
   MUX4EHD U6333 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4885), 
	.D(\ram[119][2] ), 
	.C(\ram[117][2] ), 
	.B(\ram[118][2] ), 
	.A(\ram[116][2] ));
   MUX4EHD U6334 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4886), 
	.D(\ram[115][2] ), 
	.C(\ram[113][2] ), 
	.B(\ram[114][2] ), 
	.A(\ram[112][2] ));
   MUX4EHD U6335 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4887), 
	.D(n4883), 
	.C(n4885), 
	.B(n4884), 
	.A(n4886));
   MUX4EHD U6336 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4888), 
	.D(\ram[111][2] ), 
	.C(\ram[109][2] ), 
	.B(\ram[110][2] ), 
	.A(\ram[108][2] ));
   MUX4EHD U6337 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4889), 
	.D(\ram[107][2] ), 
	.C(\ram[105][2] ), 
	.B(\ram[106][2] ), 
	.A(\ram[104][2] ));
   MUX4EHD U6338 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4890), 
	.D(\ram[103][2] ), 
	.C(\ram[101][2] ), 
	.B(\ram[102][2] ), 
	.A(\ram[100][2] ));
   MUX4EHD U6339 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4891), 
	.D(\ram[99][2] ), 
	.C(\ram[97][2] ), 
	.B(\ram[98][2] ), 
	.A(\ram[96][2] ));
   MUX4EHD U6340 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4892), 
	.D(n4888), 
	.C(n4890), 
	.B(n4889), 
	.A(n4891));
   MUX4EHD U6341 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4893), 
	.D(\ram[95][2] ), 
	.C(\ram[93][2] ), 
	.B(\ram[94][2] ), 
	.A(\ram[92][2] ));
   MUX4EHD U6342 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4894), 
	.D(\ram[91][2] ), 
	.C(\ram[89][2] ), 
	.B(\ram[90][2] ), 
	.A(\ram[88][2] ));
   MUX4EHD U6343 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4895), 
	.D(\ram[87][2] ), 
	.C(\ram[85][2] ), 
	.B(\ram[86][2] ), 
	.A(\ram[84][2] ));
   MUX4EHD U6344 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4896), 
	.D(\ram[83][2] ), 
	.C(\ram[81][2] ), 
	.B(\ram[82][2] ), 
	.A(\ram[80][2] ));
   MUX4EHD U6345 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4897), 
	.D(n4893), 
	.C(n4895), 
	.B(n4894), 
	.A(n4896));
   MUX4EHD U6346 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4898), 
	.D(\ram[79][2] ), 
	.C(\ram[77][2] ), 
	.B(\ram[78][2] ), 
	.A(\ram[76][2] ));
   MUX4EHD U6347 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4899), 
	.D(\ram[75][2] ), 
	.C(\ram[73][2] ), 
	.B(\ram[74][2] ), 
	.A(\ram[72][2] ));
   MUX4EHD U6348 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4900), 
	.D(\ram[71][2] ), 
	.C(\ram[69][2] ), 
	.B(\ram[70][2] ), 
	.A(\ram[68][2] ));
   MUX4EHD U6349 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4901), 
	.D(\ram[67][2] ), 
	.C(\ram[65][2] ), 
	.B(\ram[66][2] ), 
	.A(\ram[64][2] ));
   MUX4EHD U6350 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4902), 
	.D(n4898), 
	.C(n4900), 
	.B(n4899), 
	.A(n4901));
   MUX4EHD U6351 (.S1(n6038), 
	.S0(n7444), 
	.O(n4903), 
	.D(n4887), 
	.C(n4897), 
	.B(n4892), 
	.A(n4902));
   MUX4EHD U6352 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4904), 
	.D(\ram[63][2] ), 
	.C(\ram[61][2] ), 
	.B(\ram[62][2] ), 
	.A(\ram[60][2] ));
   MUX4EHD U6353 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4905), 
	.D(\ram[59][2] ), 
	.C(\ram[57][2] ), 
	.B(\ram[58][2] ), 
	.A(\ram[56][2] ));
   MUX4EHD U6354 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4906), 
	.D(\ram[55][2] ), 
	.C(\ram[53][2] ), 
	.B(\ram[54][2] ), 
	.A(\ram[52][2] ));
   MUX4EHD U6355 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4907), 
	.D(\ram[51][2] ), 
	.C(\ram[49][2] ), 
	.B(\ram[50][2] ), 
	.A(\ram[48][2] ));
   MUX4EHD U6356 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4908), 
	.D(n4904), 
	.C(n4906), 
	.B(n4905), 
	.A(n4907));
   MUX4EHD U6357 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4909), 
	.D(\ram[47][2] ), 
	.C(\ram[45][2] ), 
	.B(\ram[46][2] ), 
	.A(\ram[44][2] ));
   MUX4EHD U6358 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4910), 
	.D(\ram[43][2] ), 
	.C(\ram[41][2] ), 
	.B(\ram[42][2] ), 
	.A(\ram[40][2] ));
   MUX4EHD U6359 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4911), 
	.D(\ram[39][2] ), 
	.C(\ram[37][2] ), 
	.B(\ram[38][2] ), 
	.A(\ram[36][2] ));
   MUX4EHD U6360 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4912), 
	.D(\ram[35][2] ), 
	.C(\ram[33][2] ), 
	.B(\ram[34][2] ), 
	.A(\ram[32][2] ));
   MUX4EHD U6361 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4913), 
	.D(n4909), 
	.C(n4911), 
	.B(n4910), 
	.A(n4912));
   MUX4EHD U6362 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4914), 
	.D(\ram[31][2] ), 
	.C(\ram[29][2] ), 
	.B(\ram[30][2] ), 
	.A(\ram[28][2] ));
   MUX4EHD U6363 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4915), 
	.D(\ram[27][2] ), 
	.C(\ram[25][2] ), 
	.B(\ram[26][2] ), 
	.A(\ram[24][2] ));
   MUX4EHD U6364 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4916), 
	.D(\ram[23][2] ), 
	.C(\ram[21][2] ), 
	.B(\ram[22][2] ), 
	.A(\ram[20][2] ));
   MUX4EHD U6365 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4917), 
	.D(\ram[19][2] ), 
	.C(\ram[17][2] ), 
	.B(\ram[18][2] ), 
	.A(\ram[16][2] ));
   MUX4EHD U6366 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4918), 
	.D(n4914), 
	.C(n4916), 
	.B(n4915), 
	.A(n4917));
   MUX4EHD U6367 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4919), 
	.D(\ram[15][2] ), 
	.C(\ram[13][2] ), 
	.B(\ram[14][2] ), 
	.A(\ram[12][2] ));
   MUX4EHD U6368 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4920), 
	.D(\ram[11][2] ), 
	.C(\ram[9][2] ), 
	.B(\ram[10][2] ), 
	.A(\ram[8][2] ));
   MUX4EHD U6369 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4921), 
	.D(\ram[7][2] ), 
	.C(\ram[5][2] ), 
	.B(\ram[6][2] ), 
	.A(\ram[4][2] ));
   MUX4EHD U6370 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n4922), 
	.D(\ram[3][2] ), 
	.C(\ram[1][2] ), 
	.B(\ram[2][2] ), 
	.A(\ram[0][2] ));
   MUX4EHD U6371 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4923), 
	.D(n4919), 
	.C(n4921), 
	.B(n4920), 
	.A(n4922));
   MUX4EHD U6372 (.S1(n6038), 
	.S0(n7444), 
	.O(n4924), 
	.D(n4908), 
	.C(n4918), 
	.B(n4913), 
	.A(n4923));
   MUX4EHD U6373 (.S1(n6469), 
	.S0(n6470), 
	.O(N4139), 
	.D(n4861), 
	.C(n4903), 
	.B(n4882), 
	.A(n4924));
   MUX4EHD U6374 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4925), 
	.D(\ram[255][3] ), 
	.C(\ram[253][3] ), 
	.B(\ram[254][3] ), 
	.A(\ram[252][3] ));
   MUX4EHD U6375 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4926), 
	.D(\ram[251][3] ), 
	.C(\ram[249][3] ), 
	.B(\ram[250][3] ), 
	.A(\ram[248][3] ));
   MUX4EHD U6376 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4927), 
	.D(\ram[247][3] ), 
	.C(\ram[245][3] ), 
	.B(\ram[246][3] ), 
	.A(\ram[244][3] ));
   MUX4EHD U6377 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4928), 
	.D(\ram[243][3] ), 
	.C(\ram[241][3] ), 
	.B(\ram[242][3] ), 
	.A(\ram[240][3] ));
   MUX4EHD U6378 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4929), 
	.D(n4925), 
	.C(n4927), 
	.B(n4926), 
	.A(n4928));
   MUX4EHD U6379 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4930), 
	.D(\ram[239][3] ), 
	.C(\ram[237][3] ), 
	.B(\ram[238][3] ), 
	.A(\ram[236][3] ));
   MUX4EHD U6380 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4931), 
	.D(\ram[235][3] ), 
	.C(\ram[233][3] ), 
	.B(\ram[234][3] ), 
	.A(\ram[232][3] ));
   MUX4EHD U6381 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4932), 
	.D(\ram[231][3] ), 
	.C(\ram[229][3] ), 
	.B(\ram[230][3] ), 
	.A(\ram[228][3] ));
   MUX4EHD U6382 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4933), 
	.D(\ram[227][3] ), 
	.C(\ram[225][3] ), 
	.B(\ram[226][3] ), 
	.A(\ram[224][3] ));
   MUX4EHD U6383 (.S1(n6136), 
	.S0(n7442), 
	.O(n4934), 
	.D(n4930), 
	.C(n4932), 
	.B(n4931), 
	.A(n4933));
   MUX4EHD U6384 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4935), 
	.D(\ram[223][3] ), 
	.C(\ram[221][3] ), 
	.B(\ram[222][3] ), 
	.A(\ram[220][3] ));
   MUX4EHD U6385 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4936), 
	.D(\ram[219][3] ), 
	.C(\ram[217][3] ), 
	.B(\ram[218][3] ), 
	.A(\ram[216][3] ));
   MUX4EHD U6386 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4937), 
	.D(\ram[215][3] ), 
	.C(\ram[213][3] ), 
	.B(\ram[214][3] ), 
	.A(\ram[212][3] ));
   MUX4EHD U6387 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n4938), 
	.D(\ram[211][3] ), 
	.C(\ram[209][3] ), 
	.B(\ram[210][3] ), 
	.A(\ram[208][3] ));
   MUX4EHD U6388 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n4939), 
	.D(n4935), 
	.C(n4937), 
	.B(n4936), 
	.A(n4938));
   MUX4EHD U6389 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4940), 
	.D(\ram[207][3] ), 
	.C(\ram[205][3] ), 
	.B(\ram[206][3] ), 
	.A(\ram[204][3] ));
   MUX4EHD U6390 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4941), 
	.D(\ram[203][3] ), 
	.C(\ram[201][3] ), 
	.B(\ram[202][3] ), 
	.A(\ram[200][3] ));
   MUX4EHD U6391 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4942), 
	.D(\ram[199][3] ), 
	.C(\ram[197][3] ), 
	.B(\ram[198][3] ), 
	.A(\ram[196][3] ));
   MUX4EHD U6392 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n4943), 
	.D(\ram[195][3] ), 
	.C(\ram[193][3] ), 
	.B(\ram[194][3] ), 
	.A(\ram[192][3] ));
   MUX4EHD U6393 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4944), 
	.D(n4940), 
	.C(n4942), 
	.B(n4941), 
	.A(n4943));
   MUX4EHD U6394 (.S1(n6038), 
	.S0(n7444), 
	.O(n4945), 
	.D(n4929), 
	.C(n4939), 
	.B(n4934), 
	.A(n4944));
   MUX4EHD U6395 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4946), 
	.D(\ram[191][3] ), 
	.C(\ram[189][3] ), 
	.B(\ram[190][3] ), 
	.A(\ram[188][3] ));
   MUX4EHD U6396 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4947), 
	.D(\ram[187][3] ), 
	.C(\ram[185][3] ), 
	.B(\ram[186][3] ), 
	.A(\ram[184][3] ));
   MUX4EHD U6397 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n4948), 
	.D(\ram[183][3] ), 
	.C(\ram[181][3] ), 
	.B(\ram[182][3] ), 
	.A(\ram[180][3] ));
   MUX4EHD U6398 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n4949), 
	.D(\ram[179][3] ), 
	.C(\ram[177][3] ), 
	.B(\ram[178][3] ), 
	.A(\ram[176][3] ));
   MUX4EHD U6399 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n4950), 
	.D(n4946), 
	.C(n4948), 
	.B(n4947), 
	.A(n4949));
   MUX4EHD U6400 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n4951), 
	.D(\ram[175][3] ), 
	.C(\ram[173][3] ), 
	.B(\ram[174][3] ), 
	.A(\ram[172][3] ));
   MUX4EHD U6401 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4952), 
	.D(\ram[171][3] ), 
	.C(\ram[169][3] ), 
	.B(\ram[170][3] ), 
	.A(\ram[168][3] ));
   MUX4EHD U6402 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4953), 
	.D(\ram[167][3] ), 
	.C(\ram[165][3] ), 
	.B(\ram[166][3] ), 
	.A(\ram[164][3] ));
   MUX4EHD U6403 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4954), 
	.D(\ram[163][3] ), 
	.C(\ram[161][3] ), 
	.B(\ram[162][3] ), 
	.A(\ram[160][3] ));
   MUX4EHD U6404 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4955), 
	.D(n4951), 
	.C(n4953), 
	.B(n4952), 
	.A(n4954));
   MUX4EHD U6405 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4956), 
	.D(\ram[159][3] ), 
	.C(\ram[157][3] ), 
	.B(\ram[158][3] ), 
	.A(\ram[156][3] ));
   MUX4EHD U6406 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4957), 
	.D(\ram[155][3] ), 
	.C(\ram[153][3] ), 
	.B(\ram[154][3] ), 
	.A(\ram[152][3] ));
   MUX4EHD U6407 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n4958), 
	.D(\ram[151][3] ), 
	.C(\ram[149][3] ), 
	.B(\ram[150][3] ), 
	.A(\ram[148][3] ));
   MUX4EHD U6408 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4959), 
	.D(\ram[147][3] ), 
	.C(\ram[145][3] ), 
	.B(\ram[146][3] ), 
	.A(\ram[144][3] ));
   MUX4EHD U6409 (.S1(n6136), 
	.S0(n7442), 
	.O(n4960), 
	.D(n4956), 
	.C(n4958), 
	.B(n4957), 
	.A(n4959));
   MUX4EHD U6410 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4961), 
	.D(\ram[143][3] ), 
	.C(\ram[141][3] ), 
	.B(\ram[142][3] ), 
	.A(\ram[140][3] ));
   MUX4EHD U6411 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4962), 
	.D(\ram[139][3] ), 
	.C(\ram[137][3] ), 
	.B(\ram[138][3] ), 
	.A(\ram[136][3] ));
   MUX4EHD U6412 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n4963), 
	.D(\ram[135][3] ), 
	.C(\ram[133][3] ), 
	.B(\ram[134][3] ), 
	.A(\ram[132][3] ));
   MUX4EHD U6413 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n4964), 
	.D(\ram[131][3] ), 
	.C(\ram[129][3] ), 
	.B(\ram[130][3] ), 
	.A(\ram[128][3] ));
   MUX4EHD U6414 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n4965), 
	.D(n4961), 
	.C(n4963), 
	.B(n4962), 
	.A(n4964));
   MUX4EHD U6415 (.S1(n6038), 
	.S0(n7444), 
	.O(n4966), 
	.D(n4950), 
	.C(n4960), 
	.B(n4955), 
	.A(n4965));
   MUX4EHD U6416 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4967), 
	.D(\ram[127][3] ), 
	.C(\ram[125][3] ), 
	.B(\ram[126][3] ), 
	.A(\ram[124][3] ));
   MUX4EHD U6417 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4968), 
	.D(\ram[123][3] ), 
	.C(\ram[121][3] ), 
	.B(\ram[122][3] ), 
	.A(\ram[120][3] ));
   MUX4EHD U6418 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4969), 
	.D(\ram[119][3] ), 
	.C(\ram[117][3] ), 
	.B(\ram[118][3] ), 
	.A(\ram[116][3] ));
   MUX4EHD U6419 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4970), 
	.D(\ram[115][3] ), 
	.C(\ram[113][3] ), 
	.B(\ram[114][3] ), 
	.A(\ram[112][3] ));
   MUX4EHD U6420 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4971), 
	.D(n4967), 
	.C(n4969), 
	.B(n4968), 
	.A(n4970));
   MUX4EHD U6421 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n4972), 
	.D(\ram[111][3] ), 
	.C(\ram[109][3] ), 
	.B(\ram[110][3] ), 
	.A(\ram[108][3] ));
   MUX4EHD U6422 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4973), 
	.D(\ram[107][3] ), 
	.C(\ram[105][3] ), 
	.B(\ram[106][3] ), 
	.A(\ram[104][3] ));
   MUX4EHD U6423 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n4974), 
	.D(\ram[103][3] ), 
	.C(\ram[101][3] ), 
	.B(\ram[102][3] ), 
	.A(\ram[100][3] ));
   MUX4EHD U6424 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n4975), 
	.D(\ram[99][3] ), 
	.C(\ram[97][3] ), 
	.B(\ram[98][3] ), 
	.A(\ram[96][3] ));
   MUX4EHD U6425 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4976), 
	.D(n4972), 
	.C(n4974), 
	.B(n4973), 
	.A(n4975));
   MUX4EHD U6426 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4977), 
	.D(\ram[95][3] ), 
	.C(\ram[93][3] ), 
	.B(\ram[94][3] ), 
	.A(\ram[92][3] ));
   MUX4EHD U6427 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4978), 
	.D(\ram[91][3] ), 
	.C(\ram[89][3] ), 
	.B(\ram[90][3] ), 
	.A(\ram[88][3] ));
   MUX4EHD U6428 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n4979), 
	.D(\ram[87][3] ), 
	.C(\ram[85][3] ), 
	.B(\ram[86][3] ), 
	.A(\ram[84][3] ));
   MUX4EHD U6429 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n4980), 
	.D(\ram[83][3] ), 
	.C(\ram[81][3] ), 
	.B(\ram[82][3] ), 
	.A(\ram[80][3] ));
   MUX4EHD U6430 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n4981), 
	.D(n4977), 
	.C(n4979), 
	.B(n4978), 
	.A(n4980));
   MUX4EHD U6431 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4982), 
	.D(\ram[79][3] ), 
	.C(\ram[77][3] ), 
	.B(\ram[78][3] ), 
	.A(\ram[76][3] ));
   MUX4EHD U6432 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4983), 
	.D(\ram[75][3] ), 
	.C(\ram[73][3] ), 
	.B(\ram[74][3] ), 
	.A(\ram[72][3] ));
   MUX4EHD U6433 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4984), 
	.D(\ram[71][3] ), 
	.C(\ram[69][3] ), 
	.B(\ram[70][3] ), 
	.A(\ram[68][3] ));
   MUX4EHD U6434 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n4985), 
	.D(\ram[67][3] ), 
	.C(\ram[65][3] ), 
	.B(\ram[66][3] ), 
	.A(\ram[64][3] ));
   MUX4EHD U6435 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n4986), 
	.D(n4982), 
	.C(n4984), 
	.B(n4983), 
	.A(n4985));
   MUX4EHD U6436 (.S1(n6038), 
	.S0(n7444), 
	.O(n4987), 
	.D(n4971), 
	.C(n4981), 
	.B(n4976), 
	.A(n4986));
   MUX4EHD U6437 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4988), 
	.D(\ram[63][3] ), 
	.C(\ram[61][3] ), 
	.B(\ram[62][3] ), 
	.A(\ram[60][3] ));
   MUX4EHD U6438 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4989), 
	.D(\ram[59][3] ), 
	.C(\ram[57][3] ), 
	.B(\ram[58][3] ), 
	.A(\ram[56][3] ));
   MUX4EHD U6439 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4990), 
	.D(\ram[55][3] ), 
	.C(\ram[53][3] ), 
	.B(\ram[54][3] ), 
	.A(\ram[52][3] ));
   MUX4EHD U6440 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n4991), 
	.D(\ram[51][3] ), 
	.C(\ram[49][3] ), 
	.B(\ram[50][3] ), 
	.A(\ram[48][3] ));
   MUX4EHD U6441 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4992), 
	.D(n4988), 
	.C(n4990), 
	.B(n4989), 
	.A(n4991));
   MUX4EHD U6442 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4993), 
	.D(\ram[47][3] ), 
	.C(\ram[45][3] ), 
	.B(\ram[46][3] ), 
	.A(\ram[44][3] ));
   MUX4EHD U6443 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4994), 
	.D(\ram[43][3] ), 
	.C(\ram[41][3] ), 
	.B(\ram[42][3] ), 
	.A(\ram[40][3] ));
   MUX4EHD U6444 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4995), 
	.D(\ram[39][3] ), 
	.C(\ram[37][3] ), 
	.B(\ram[38][3] ), 
	.A(\ram[36][3] ));
   MUX4EHD U6445 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n4996), 
	.D(\ram[35][3] ), 
	.C(\ram[33][3] ), 
	.B(\ram[34][3] ), 
	.A(\ram[32][3] ));
   MUX4EHD U6446 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n4997), 
	.D(n4993), 
	.C(n4995), 
	.B(n4994), 
	.A(n4996));
   MUX4EHD U6447 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n4998), 
	.D(\ram[31][3] ), 
	.C(\ram[29][3] ), 
	.B(\ram[30][3] ), 
	.A(\ram[28][3] ));
   MUX4EHD U6448 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n4999), 
	.D(\ram[27][3] ), 
	.C(\ram[25][3] ), 
	.B(\ram[26][3] ), 
	.A(\ram[24][3] ));
   MUX4EHD U6449 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5000), 
	.D(\ram[23][3] ), 
	.C(\ram[21][3] ), 
	.B(\ram[22][3] ), 
	.A(\ram[20][3] ));
   MUX4EHD U6450 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5001), 
	.D(\ram[19][3] ), 
	.C(\ram[17][3] ), 
	.B(\ram[18][3] ), 
	.A(\ram[16][3] ));
   MUX4EHD U6451 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5002), 
	.D(n4998), 
	.C(n5000), 
	.B(n4999), 
	.A(n5001));
   MUX4EHD U6452 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5003), 
	.D(\ram[15][3] ), 
	.C(\ram[13][3] ), 
	.B(\ram[14][3] ), 
	.A(\ram[12][3] ));
   MUX4EHD U6453 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5004), 
	.D(\ram[11][3] ), 
	.C(\ram[9][3] ), 
	.B(\ram[10][3] ), 
	.A(\ram[8][3] ));
   MUX4EHD U6454 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5005), 
	.D(\ram[7][3] ), 
	.C(\ram[5][3] ), 
	.B(\ram[6][3] ), 
	.A(\ram[4][3] ));
   MUX4EHD U6455 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5006), 
	.D(\ram[3][3] ), 
	.C(\ram[1][3] ), 
	.B(\ram[2][3] ), 
	.A(\ram[0][3] ));
   MUX4EHD U6456 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5007), 
	.D(n5003), 
	.C(n5005), 
	.B(n5004), 
	.A(n5006));
   MUX4EHD U6457 (.S1(n6038), 
	.S0(n7444), 
	.O(n5008), 
	.D(n4992), 
	.C(n5002), 
	.B(n4997), 
	.A(n5007));
   MUX4EHD U6458 (.S1(n6469), 
	.S0(n6470), 
	.O(N4138), 
	.D(n4945), 
	.C(n4987), 
	.B(n4966), 
	.A(n5008));
   MUX4EHD U6459 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5009), 
	.D(\ram[255][4] ), 
	.C(\ram[253][4] ), 
	.B(\ram[254][4] ), 
	.A(\ram[252][4] ));
   MUX4EHD U6460 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5010), 
	.D(\ram[251][4] ), 
	.C(\ram[249][4] ), 
	.B(\ram[250][4] ), 
	.A(\ram[248][4] ));
   MUX4EHD U6461 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5011), 
	.D(\ram[247][4] ), 
	.C(\ram[245][4] ), 
	.B(\ram[246][4] ), 
	.A(\ram[244][4] ));
   MUX4EHD U6462 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5012), 
	.D(\ram[243][4] ), 
	.C(\ram[241][4] ), 
	.B(\ram[242][4] ), 
	.A(\ram[240][4] ));
   MUX4EHD U6463 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5013), 
	.D(n5009), 
	.C(n5011), 
	.B(n5010), 
	.A(n5012));
   MUX4EHD U6464 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5014), 
	.D(\ram[239][4] ), 
	.C(\ram[237][4] ), 
	.B(\ram[238][4] ), 
	.A(\ram[236][4] ));
   MUX4EHD U6465 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5015), 
	.D(\ram[235][4] ), 
	.C(\ram[233][4] ), 
	.B(\ram[234][4] ), 
	.A(\ram[232][4] ));
   MUX4EHD U6466 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5016), 
	.D(\ram[231][4] ), 
	.C(\ram[229][4] ), 
	.B(\ram[230][4] ), 
	.A(\ram[228][4] ));
   MUX4EHD U6467 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5017), 
	.D(\ram[227][4] ), 
	.C(\ram[225][4] ), 
	.B(\ram[226][4] ), 
	.A(\ram[224][4] ));
   MUX4EHD U6468 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5018), 
	.D(n5014), 
	.C(n5016), 
	.B(n5015), 
	.A(n5017));
   MUX4EHD U6469 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5019), 
	.D(\ram[223][4] ), 
	.C(\ram[221][4] ), 
	.B(\ram[222][4] ), 
	.A(\ram[220][4] ));
   MUX4EHD U6470 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5020), 
	.D(\ram[219][4] ), 
	.C(\ram[217][4] ), 
	.B(\ram[218][4] ), 
	.A(\ram[216][4] ));
   MUX4EHD U6471 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5021), 
	.D(\ram[215][4] ), 
	.C(\ram[213][4] ), 
	.B(\ram[214][4] ), 
	.A(\ram[212][4] ));
   MUX4EHD U6472 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5022), 
	.D(\ram[211][4] ), 
	.C(\ram[209][4] ), 
	.B(\ram[210][4] ), 
	.A(\ram[208][4] ));
   MUX4EHD U6473 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5023), 
	.D(n5019), 
	.C(n5021), 
	.B(n5020), 
	.A(n5022));
   MUX4EHD U6474 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5024), 
	.D(\ram[207][4] ), 
	.C(\ram[205][4] ), 
	.B(\ram[206][4] ), 
	.A(\ram[204][4] ));
   MUX4EHD U6475 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5025), 
	.D(\ram[203][4] ), 
	.C(\ram[201][4] ), 
	.B(\ram[202][4] ), 
	.A(\ram[200][4] ));
   MUX4EHD U6476 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5026), 
	.D(\ram[199][4] ), 
	.C(\ram[197][4] ), 
	.B(\ram[198][4] ), 
	.A(\ram[196][4] ));
   MUX4EHD U6477 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5027), 
	.D(\ram[195][4] ), 
	.C(\ram[193][4] ), 
	.B(\ram[194][4] ), 
	.A(\ram[192][4] ));
   MUX4EHD U6478 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5028), 
	.D(n5024), 
	.C(n5026), 
	.B(n5025), 
	.A(n5027));
   MUX4EHD U6479 (.S1(n6038), 
	.S0(n7444), 
	.O(n5029), 
	.D(n5013), 
	.C(n5023), 
	.B(n5018), 
	.A(n5028));
   MUX4EHD U6480 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5030), 
	.D(\ram[191][4] ), 
	.C(\ram[189][4] ), 
	.B(\ram[190][4] ), 
	.A(\ram[188][4] ));
   MUX4EHD U6481 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5031), 
	.D(\ram[187][4] ), 
	.C(\ram[185][4] ), 
	.B(\ram[186][4] ), 
	.A(\ram[184][4] ));
   MUX4EHD U6482 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5032), 
	.D(\ram[183][4] ), 
	.C(\ram[181][4] ), 
	.B(\ram[182][4] ), 
	.A(\ram[180][4] ));
   MUX4EHD U6483 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5033), 
	.D(\ram[179][4] ), 
	.C(\ram[177][4] ), 
	.B(\ram[178][4] ), 
	.A(\ram[176][4] ));
   MUX4EHD U6484 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5034), 
	.D(n5030), 
	.C(n5032), 
	.B(n5031), 
	.A(n5033));
   MUX4EHD U6485 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5035), 
	.D(\ram[175][4] ), 
	.C(\ram[173][4] ), 
	.B(\ram[174][4] ), 
	.A(\ram[172][4] ));
   MUX4EHD U6486 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5036), 
	.D(\ram[171][4] ), 
	.C(\ram[169][4] ), 
	.B(\ram[170][4] ), 
	.A(\ram[168][4] ));
   MUX4EHD U6487 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5037), 
	.D(\ram[167][4] ), 
	.C(\ram[165][4] ), 
	.B(\ram[166][4] ), 
	.A(\ram[164][4] ));
   MUX4EHD U6488 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5038), 
	.D(\ram[163][4] ), 
	.C(\ram[161][4] ), 
	.B(\ram[162][4] ), 
	.A(\ram[160][4] ));
   MUX4EHD U6489 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5039), 
	.D(n5035), 
	.C(n5037), 
	.B(n5036), 
	.A(n5038));
   MUX4EHD U6490 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5040), 
	.D(\ram[159][4] ), 
	.C(\ram[157][4] ), 
	.B(\ram[158][4] ), 
	.A(\ram[156][4] ));
   MUX4EHD U6491 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5041), 
	.D(\ram[155][4] ), 
	.C(\ram[153][4] ), 
	.B(\ram[154][4] ), 
	.A(\ram[152][4] ));
   MUX4EHD U6492 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5042), 
	.D(\ram[151][4] ), 
	.C(\ram[149][4] ), 
	.B(\ram[150][4] ), 
	.A(\ram[148][4] ));
   MUX4EHD U6493 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5043), 
	.D(\ram[147][4] ), 
	.C(\ram[145][4] ), 
	.B(\ram[146][4] ), 
	.A(\ram[144][4] ));
   MUX4EHD U6494 (.S1(n6136), 
	.S0(n7442), 
	.O(n5044), 
	.D(n5040), 
	.C(n5042), 
	.B(n5041), 
	.A(n5043));
   MUX4EHD U6495 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5045), 
	.D(\ram[143][4] ), 
	.C(\ram[141][4] ), 
	.B(\ram[142][4] ), 
	.A(\ram[140][4] ));
   MUX4EHD U6496 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5046), 
	.D(\ram[139][4] ), 
	.C(\ram[137][4] ), 
	.B(\ram[138][4] ), 
	.A(\ram[136][4] ));
   MUX4EHD U6497 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5047), 
	.D(\ram[135][4] ), 
	.C(\ram[133][4] ), 
	.B(\ram[134][4] ), 
	.A(\ram[132][4] ));
   MUX4EHD U6498 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5048), 
	.D(\ram[131][4] ), 
	.C(\ram[129][4] ), 
	.B(\ram[130][4] ), 
	.A(\ram[128][4] ));
   MUX4EHD U6499 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5049), 
	.D(n5045), 
	.C(n5047), 
	.B(n5046), 
	.A(n5048));
   MUX4EHD U6500 (.S1(n6038), 
	.S0(n7444), 
	.O(n5050), 
	.D(n5034), 
	.C(n5044), 
	.B(n5039), 
	.A(n5049));
   MUX4EHD U6501 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5051), 
	.D(\ram[127][4] ), 
	.C(\ram[125][4] ), 
	.B(\ram[126][4] ), 
	.A(\ram[124][4] ));
   MUX4EHD U6502 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5052), 
	.D(\ram[123][4] ), 
	.C(\ram[121][4] ), 
	.B(\ram[122][4] ), 
	.A(\ram[120][4] ));
   MUX4EHD U6503 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5053), 
	.D(\ram[119][4] ), 
	.C(\ram[117][4] ), 
	.B(\ram[118][4] ), 
	.A(\ram[116][4] ));
   MUX4EHD U6504 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5054), 
	.D(\ram[115][4] ), 
	.C(\ram[113][4] ), 
	.B(\ram[114][4] ), 
	.A(\ram[112][4] ));
   MUX4EHD U6505 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5055), 
	.D(n5051), 
	.C(n5053), 
	.B(n5052), 
	.A(n5054));
   MUX4EHD U6506 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5056), 
	.D(\ram[111][4] ), 
	.C(\ram[109][4] ), 
	.B(\ram[110][4] ), 
	.A(\ram[108][4] ));
   MUX4EHD U6507 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5057), 
	.D(\ram[107][4] ), 
	.C(\ram[105][4] ), 
	.B(\ram[106][4] ), 
	.A(\ram[104][4] ));
   MUX4EHD U6508 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5058), 
	.D(\ram[103][4] ), 
	.C(\ram[101][4] ), 
	.B(\ram[102][4] ), 
	.A(\ram[100][4] ));
   MUX4EHD U6509 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5059), 
	.D(\ram[99][4] ), 
	.C(\ram[97][4] ), 
	.B(\ram[98][4] ), 
	.A(\ram[96][4] ));
   MUX4EHD U6510 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5060), 
	.D(n5056), 
	.C(n5058), 
	.B(n5057), 
	.A(n5059));
   MUX4EHD U6511 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5061), 
	.D(\ram[95][4] ), 
	.C(\ram[93][4] ), 
	.B(\ram[94][4] ), 
	.A(\ram[92][4] ));
   MUX4EHD U6512 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5062), 
	.D(\ram[91][4] ), 
	.C(\ram[89][4] ), 
	.B(\ram[90][4] ), 
	.A(\ram[88][4] ));
   MUX4EHD U6513 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5063), 
	.D(\ram[87][4] ), 
	.C(\ram[85][4] ), 
	.B(\ram[86][4] ), 
	.A(\ram[84][4] ));
   MUX4EHD U6514 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5064), 
	.D(\ram[83][4] ), 
	.C(\ram[81][4] ), 
	.B(\ram[82][4] ), 
	.A(\ram[80][4] ));
   MUX4EHD U6515 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5065), 
	.D(n5061), 
	.C(n5063), 
	.B(n5062), 
	.A(n5064));
   MUX4EHD U6516 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5066), 
	.D(\ram[79][4] ), 
	.C(\ram[77][4] ), 
	.B(\ram[78][4] ), 
	.A(\ram[76][4] ));
   MUX4EHD U6517 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5067), 
	.D(\ram[75][4] ), 
	.C(\ram[73][4] ), 
	.B(\ram[74][4] ), 
	.A(\ram[72][4] ));
   MUX4EHD U6518 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5068), 
	.D(\ram[71][4] ), 
	.C(\ram[69][4] ), 
	.B(\ram[70][4] ), 
	.A(\ram[68][4] ));
   MUX4EHD U6519 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5069), 
	.D(\ram[67][4] ), 
	.C(\ram[65][4] ), 
	.B(\ram[66][4] ), 
	.A(\ram[64][4] ));
   MUX4EHD U6520 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5070), 
	.D(n5066), 
	.C(n5068), 
	.B(n5067), 
	.A(n5069));
   MUX4EHD U6521 (.S1(n6038), 
	.S0(n7444), 
	.O(n5071), 
	.D(n5055), 
	.C(n5065), 
	.B(n5060), 
	.A(n5070));
   MUX4EHD U6522 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5072), 
	.D(\ram[63][4] ), 
	.C(\ram[61][4] ), 
	.B(\ram[62][4] ), 
	.A(\ram[60][4] ));
   MUX4EHD U6523 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5073), 
	.D(\ram[59][4] ), 
	.C(\ram[57][4] ), 
	.B(\ram[58][4] ), 
	.A(\ram[56][4] ));
   MUX4EHD U6524 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5074), 
	.D(\ram[55][4] ), 
	.C(\ram[53][4] ), 
	.B(\ram[54][4] ), 
	.A(\ram[52][4] ));
   MUX4EHD U6525 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5075), 
	.D(\ram[51][4] ), 
	.C(\ram[49][4] ), 
	.B(\ram[50][4] ), 
	.A(\ram[48][4] ));
   MUX4EHD U6526 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5076), 
	.D(n5072), 
	.C(n5074), 
	.B(n5073), 
	.A(n5075));
   MUX4EHD U6527 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5077), 
	.D(\ram[47][4] ), 
	.C(\ram[45][4] ), 
	.B(\ram[46][4] ), 
	.A(\ram[44][4] ));
   MUX4EHD U6528 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5078), 
	.D(\ram[43][4] ), 
	.C(\ram[41][4] ), 
	.B(\ram[42][4] ), 
	.A(\ram[40][4] ));
   MUX4EHD U6529 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5079), 
	.D(\ram[39][4] ), 
	.C(\ram[37][4] ), 
	.B(\ram[38][4] ), 
	.A(\ram[36][4] ));
   MUX4EHD U6530 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5080), 
	.D(\ram[35][4] ), 
	.C(\ram[33][4] ), 
	.B(\ram[34][4] ), 
	.A(\ram[32][4] ));
   MUX4EHD U6531 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5081), 
	.D(n5077), 
	.C(n5079), 
	.B(n5078), 
	.A(n5080));
   MUX4EHD U6532 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5082), 
	.D(\ram[31][4] ), 
	.C(\ram[29][4] ), 
	.B(\ram[30][4] ), 
	.A(\ram[28][4] ));
   MUX4EHD U6533 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5083), 
	.D(\ram[27][4] ), 
	.C(\ram[25][4] ), 
	.B(\ram[26][4] ), 
	.A(\ram[24][4] ));
   MUX4EHD U6534 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5084), 
	.D(\ram[23][4] ), 
	.C(\ram[21][4] ), 
	.B(\ram[22][4] ), 
	.A(\ram[20][4] ));
   MUX4EHD U6535 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5085), 
	.D(\ram[19][4] ), 
	.C(\ram[17][4] ), 
	.B(\ram[18][4] ), 
	.A(\ram[16][4] ));
   MUX4EHD U6536 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5086), 
	.D(n5082), 
	.C(n5084), 
	.B(n5083), 
	.A(n5085));
   MUX4EHD U6537 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5087), 
	.D(\ram[15][4] ), 
	.C(\ram[13][4] ), 
	.B(\ram[14][4] ), 
	.A(\ram[12][4] ));
   MUX4EHD U6538 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5088), 
	.D(\ram[11][4] ), 
	.C(\ram[9][4] ), 
	.B(\ram[10][4] ), 
	.A(\ram[8][4] ));
   MUX4EHD U6539 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5089), 
	.D(\ram[7][4] ), 
	.C(\ram[5][4] ), 
	.B(\ram[6][4] ), 
	.A(\ram[4][4] ));
   MUX4EHD U6540 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5090), 
	.D(\ram[3][4] ), 
	.C(\ram[1][4] ), 
	.B(\ram[2][4] ), 
	.A(\ram[0][4] ));
   MUX4EHD U6541 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5091), 
	.D(n5087), 
	.C(n5089), 
	.B(n5088), 
	.A(n5090));
   MUX4EHD U6542 (.S1(n6038), 
	.S0(n7444), 
	.O(n5092), 
	.D(n5076), 
	.C(n5086), 
	.B(n5081), 
	.A(n5091));
   MUX4EHD U6543 (.S1(n6469), 
	.S0(n6470), 
	.O(N4137), 
	.D(n5029), 
	.C(n5071), 
	.B(n5050), 
	.A(n5092));
   MUX4EHD U6544 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5093), 
	.D(\ram[255][5] ), 
	.C(\ram[253][5] ), 
	.B(\ram[254][5] ), 
	.A(\ram[252][5] ));
   MUX4EHD U6545 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5094), 
	.D(\ram[251][5] ), 
	.C(\ram[249][5] ), 
	.B(\ram[250][5] ), 
	.A(\ram[248][5] ));
   MUX4EHD U6546 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5095), 
	.D(\ram[247][5] ), 
	.C(\ram[245][5] ), 
	.B(\ram[246][5] ), 
	.A(\ram[244][5] ));
   MUX4EHD U6547 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5096), 
	.D(\ram[243][5] ), 
	.C(\ram[241][5] ), 
	.B(\ram[242][5] ), 
	.A(\ram[240][5] ));
   MUX4EHD U6548 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5097), 
	.D(n5093), 
	.C(n5095), 
	.B(n5094), 
	.A(n5096));
   MUX4EHD U6549 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5098), 
	.D(\ram[239][5] ), 
	.C(\ram[237][5] ), 
	.B(\ram[238][5] ), 
	.A(\ram[236][5] ));
   MUX4EHD U6550 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5099), 
	.D(\ram[235][5] ), 
	.C(\ram[233][5] ), 
	.B(\ram[234][5] ), 
	.A(\ram[232][5] ));
   MUX4EHD U6551 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5100), 
	.D(\ram[231][5] ), 
	.C(\ram[229][5] ), 
	.B(\ram[230][5] ), 
	.A(\ram[228][5] ));
   MUX4EHD U6552 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5101), 
	.D(\ram[227][5] ), 
	.C(\ram[225][5] ), 
	.B(\ram[226][5] ), 
	.A(\ram[224][5] ));
   MUX4EHD U6553 (.S1(n6136), 
	.S0(n7442), 
	.O(n5102), 
	.D(n5098), 
	.C(n5100), 
	.B(n5099), 
	.A(n5101));
   MUX4EHD U6554 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5103), 
	.D(\ram[223][5] ), 
	.C(\ram[221][5] ), 
	.B(\ram[222][5] ), 
	.A(\ram[220][5] ));
   MUX4EHD U6555 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5104), 
	.D(\ram[219][5] ), 
	.C(\ram[217][5] ), 
	.B(\ram[218][5] ), 
	.A(\ram[216][5] ));
   MUX4EHD U6556 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5105), 
	.D(\ram[215][5] ), 
	.C(\ram[213][5] ), 
	.B(\ram[214][5] ), 
	.A(\ram[212][5] ));
   MUX4EHD U6557 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5106), 
	.D(\ram[211][5] ), 
	.C(\ram[209][5] ), 
	.B(\ram[210][5] ), 
	.A(\ram[208][5] ));
   MUX4EHD U6558 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5107), 
	.D(n5103), 
	.C(n5105), 
	.B(n5104), 
	.A(n5106));
   MUX4EHD U6559 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5108), 
	.D(\ram[207][5] ), 
	.C(\ram[205][5] ), 
	.B(\ram[206][5] ), 
	.A(\ram[204][5] ));
   MUX4EHD U6560 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5109), 
	.D(\ram[203][5] ), 
	.C(\ram[201][5] ), 
	.B(\ram[202][5] ), 
	.A(\ram[200][5] ));
   MUX4EHD U6561 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5110), 
	.D(\ram[199][5] ), 
	.C(\ram[197][5] ), 
	.B(\ram[198][5] ), 
	.A(\ram[196][5] ));
   MUX4EHD U6562 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5111), 
	.D(\ram[195][5] ), 
	.C(\ram[193][5] ), 
	.B(\ram[194][5] ), 
	.A(\ram[192][5] ));
   MUX4EHD U6563 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5112), 
	.D(n5108), 
	.C(n5110), 
	.B(n5109), 
	.A(n5111));
   MUX4EHD U6564 (.S1(n6038), 
	.S0(n7444), 
	.O(n5113), 
	.D(n5097), 
	.C(n5107), 
	.B(n5102), 
	.A(n5112));
   MUX4EHD U6565 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5114), 
	.D(\ram[191][5] ), 
	.C(\ram[189][5] ), 
	.B(\ram[190][5] ), 
	.A(\ram[188][5] ));
   MUX4EHD U6566 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5115), 
	.D(\ram[187][5] ), 
	.C(\ram[185][5] ), 
	.B(\ram[186][5] ), 
	.A(\ram[184][5] ));
   MUX4EHD U6567 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5116), 
	.D(\ram[183][5] ), 
	.C(\ram[181][5] ), 
	.B(\ram[182][5] ), 
	.A(\ram[180][5] ));
   MUX4EHD U6568 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5117), 
	.D(\ram[179][5] ), 
	.C(\ram[177][5] ), 
	.B(\ram[178][5] ), 
	.A(\ram[176][5] ));
   MUX4EHD U6569 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5118), 
	.D(n5114), 
	.C(n5116), 
	.B(n5115), 
	.A(n5117));
   MUX4EHD U6570 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5119), 
	.D(\ram[175][5] ), 
	.C(\ram[173][5] ), 
	.B(\ram[174][5] ), 
	.A(\ram[172][5] ));
   MUX4EHD U6571 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5120), 
	.D(\ram[171][5] ), 
	.C(\ram[169][5] ), 
	.B(\ram[170][5] ), 
	.A(\ram[168][5] ));
   MUX4EHD U6572 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5121), 
	.D(\ram[167][5] ), 
	.C(\ram[165][5] ), 
	.B(\ram[166][5] ), 
	.A(\ram[164][5] ));
   MUX4EHD U6573 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5122), 
	.D(\ram[163][5] ), 
	.C(\ram[161][5] ), 
	.B(\ram[162][5] ), 
	.A(\ram[160][5] ));
   MUX4EHD U6574 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5123), 
	.D(n5119), 
	.C(n5121), 
	.B(n5120), 
	.A(n5122));
   MUX4EHD U6575 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5124), 
	.D(\ram[159][5] ), 
	.C(\ram[157][5] ), 
	.B(\ram[158][5] ), 
	.A(\ram[156][5] ));
   MUX4EHD U6576 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5125), 
	.D(\ram[155][5] ), 
	.C(\ram[153][5] ), 
	.B(\ram[154][5] ), 
	.A(\ram[152][5] ));
   MUX4EHD U6577 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5126), 
	.D(\ram[151][5] ), 
	.C(\ram[149][5] ), 
	.B(\ram[150][5] ), 
	.A(\ram[148][5] ));
   MUX4EHD U6578 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5127), 
	.D(\ram[147][5] ), 
	.C(\ram[145][5] ), 
	.B(\ram[146][5] ), 
	.A(\ram[144][5] ));
   MUX4EHD U6579 (.S1(n6136), 
	.S0(n7442), 
	.O(n5128), 
	.D(n5124), 
	.C(n5126), 
	.B(n5125), 
	.A(n5127));
   MUX4EHD U6580 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5129), 
	.D(\ram[143][5] ), 
	.C(\ram[141][5] ), 
	.B(\ram[142][5] ), 
	.A(\ram[140][5] ));
   MUX4EHD U6581 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5130), 
	.D(\ram[139][5] ), 
	.C(\ram[137][5] ), 
	.B(\ram[138][5] ), 
	.A(\ram[136][5] ));
   MUX4EHD U6582 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5131), 
	.D(\ram[135][5] ), 
	.C(\ram[133][5] ), 
	.B(\ram[134][5] ), 
	.A(\ram[132][5] ));
   MUX4EHD U6583 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5132), 
	.D(\ram[131][5] ), 
	.C(\ram[129][5] ), 
	.B(\ram[130][5] ), 
	.A(\ram[128][5] ));
   MUX4EHD U6584 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5133), 
	.D(n5129), 
	.C(n5131), 
	.B(n5130), 
	.A(n5132));
   MUX4EHD U6585 (.S1(n6038), 
	.S0(n7444), 
	.O(n5134), 
	.D(n5118), 
	.C(n5128), 
	.B(n5123), 
	.A(n5133));
   MUX4EHD U6586 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5135), 
	.D(\ram[127][5] ), 
	.C(\ram[125][5] ), 
	.B(\ram[126][5] ), 
	.A(\ram[124][5] ));
   MUX4EHD U6587 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5136), 
	.D(\ram[123][5] ), 
	.C(\ram[121][5] ), 
	.B(\ram[122][5] ), 
	.A(\ram[120][5] ));
   MUX4EHD U6588 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5137), 
	.D(\ram[119][5] ), 
	.C(\ram[117][5] ), 
	.B(\ram[118][5] ), 
	.A(\ram[116][5] ));
   MUX4EHD U6589 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5138), 
	.D(\ram[115][5] ), 
	.C(\ram[113][5] ), 
	.B(\ram[114][5] ), 
	.A(\ram[112][5] ));
   MUX4EHD U6590 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5139), 
	.D(n5135), 
	.C(n5137), 
	.B(n5136), 
	.A(n5138));
   MUX4EHD U6591 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5140), 
	.D(\ram[111][5] ), 
	.C(\ram[109][5] ), 
	.B(\ram[110][5] ), 
	.A(\ram[108][5] ));
   MUX4EHD U6592 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5141), 
	.D(\ram[107][5] ), 
	.C(\ram[105][5] ), 
	.B(\ram[106][5] ), 
	.A(\ram[104][5] ));
   MUX4EHD U6593 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5142), 
	.D(\ram[103][5] ), 
	.C(\ram[101][5] ), 
	.B(\ram[102][5] ), 
	.A(\ram[100][5] ));
   MUX4EHD U6594 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5143), 
	.D(\ram[99][5] ), 
	.C(\ram[97][5] ), 
	.B(\ram[98][5] ), 
	.A(\ram[96][5] ));
   MUX4EHD U6595 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5144), 
	.D(n5140), 
	.C(n5142), 
	.B(n5141), 
	.A(n5143));
   MUX4EHD U6596 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5145), 
	.D(\ram[95][5] ), 
	.C(\ram[93][5] ), 
	.B(\ram[94][5] ), 
	.A(\ram[92][5] ));
   MUX4EHD U6597 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5146), 
	.D(\ram[91][5] ), 
	.C(\ram[89][5] ), 
	.B(\ram[90][5] ), 
	.A(\ram[88][5] ));
   MUX4EHD U6598 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5147), 
	.D(\ram[87][5] ), 
	.C(\ram[85][5] ), 
	.B(\ram[86][5] ), 
	.A(\ram[84][5] ));
   MUX4EHD U6599 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5148), 
	.D(\ram[83][5] ), 
	.C(\ram[81][5] ), 
	.B(\ram[82][5] ), 
	.A(\ram[80][5] ));
   MUX4EHD U6600 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5149), 
	.D(n5145), 
	.C(n5147), 
	.B(n5146), 
	.A(n5148));
   MUX4EHD U6601 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5150), 
	.D(\ram[79][5] ), 
	.C(\ram[77][5] ), 
	.B(\ram[78][5] ), 
	.A(\ram[76][5] ));
   MUX4EHD U6602 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5151), 
	.D(\ram[75][5] ), 
	.C(\ram[73][5] ), 
	.B(\ram[74][5] ), 
	.A(\ram[72][5] ));
   MUX4EHD U6603 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5152), 
	.D(\ram[71][5] ), 
	.C(\ram[69][5] ), 
	.B(\ram[70][5] ), 
	.A(\ram[68][5] ));
   MUX4EHD U6604 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5153), 
	.D(\ram[67][5] ), 
	.C(\ram[65][5] ), 
	.B(\ram[66][5] ), 
	.A(\ram[64][5] ));
   MUX4EHD U6605 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5154), 
	.D(n5150), 
	.C(n5152), 
	.B(n5151), 
	.A(n5153));
   MUX4EHD U6606 (.S1(n6038), 
	.S0(n7444), 
	.O(n5155), 
	.D(n5139), 
	.C(n5149), 
	.B(n5144), 
	.A(n5154));
   MUX4EHD U6607 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5156), 
	.D(\ram[63][5] ), 
	.C(\ram[61][5] ), 
	.B(\ram[62][5] ), 
	.A(\ram[60][5] ));
   MUX4EHD U6608 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5157), 
	.D(\ram[59][5] ), 
	.C(\ram[57][5] ), 
	.B(\ram[58][5] ), 
	.A(\ram[56][5] ));
   MUX4EHD U6609 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5158), 
	.D(\ram[55][5] ), 
	.C(\ram[53][5] ), 
	.B(\ram[54][5] ), 
	.A(\ram[52][5] ));
   MUX4EHD U6610 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5159), 
	.D(\ram[51][5] ), 
	.C(\ram[49][5] ), 
	.B(\ram[50][5] ), 
	.A(\ram[48][5] ));
   MUX4EHD U6611 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5160), 
	.D(n5156), 
	.C(n5158), 
	.B(n5157), 
	.A(n5159));
   MUX4EHD U6612 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5161), 
	.D(\ram[47][5] ), 
	.C(\ram[45][5] ), 
	.B(\ram[46][5] ), 
	.A(\ram[44][5] ));
   MUX4EHD U6613 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5162), 
	.D(\ram[43][5] ), 
	.C(\ram[41][5] ), 
	.B(\ram[42][5] ), 
	.A(\ram[40][5] ));
   MUX4EHD U6614 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5163), 
	.D(\ram[39][5] ), 
	.C(\ram[37][5] ), 
	.B(\ram[38][5] ), 
	.A(\ram[36][5] ));
   MUX4EHD U6615 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5164), 
	.D(\ram[35][5] ), 
	.C(\ram[33][5] ), 
	.B(\ram[34][5] ), 
	.A(\ram[32][5] ));
   MUX4EHD U6616 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5165), 
	.D(n5161), 
	.C(n5163), 
	.B(n5162), 
	.A(n5164));
   MUX4EHD U6617 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5166), 
	.D(\ram[31][5] ), 
	.C(\ram[29][5] ), 
	.B(\ram[30][5] ), 
	.A(\ram[28][5] ));
   MUX4EHD U6618 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5167), 
	.D(\ram[27][5] ), 
	.C(\ram[25][5] ), 
	.B(\ram[26][5] ), 
	.A(\ram[24][5] ));
   MUX4EHD U6619 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5168), 
	.D(\ram[23][5] ), 
	.C(\ram[21][5] ), 
	.B(\ram[22][5] ), 
	.A(\ram[20][5] ));
   MUX4EHD U6620 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5169), 
	.D(\ram[19][5] ), 
	.C(\ram[17][5] ), 
	.B(\ram[18][5] ), 
	.A(\ram[16][5] ));
   MUX4EHD U6621 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5170), 
	.D(n5166), 
	.C(n5168), 
	.B(n5167), 
	.A(n5169));
   MUX4EHD U6622 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5171), 
	.D(\ram[15][5] ), 
	.C(\ram[13][5] ), 
	.B(\ram[14][5] ), 
	.A(\ram[12][5] ));
   MUX4EHD U6623 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5172), 
	.D(\ram[11][5] ), 
	.C(\ram[9][5] ), 
	.B(\ram[10][5] ), 
	.A(\ram[8][5] ));
   MUX4EHD U6624 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5173), 
	.D(\ram[7][5] ), 
	.C(\ram[5][5] ), 
	.B(\ram[6][5] ), 
	.A(\ram[4][5] ));
   MUX4EHD U6625 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5174), 
	.D(\ram[3][5] ), 
	.C(\ram[1][5] ), 
	.B(\ram[2][5] ), 
	.A(\ram[0][5] ));
   MUX4EHD U6626 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5175), 
	.D(n5171), 
	.C(n5173), 
	.B(n5172), 
	.A(n5174));
   MUX4EHD U6627 (.S1(n6038), 
	.S0(n7444), 
	.O(n5176), 
	.D(n5160), 
	.C(n5170), 
	.B(n5165), 
	.A(n5175));
   MUX4EHD U6628 (.S1(n6469), 
	.S0(n6470), 
	.O(N4136), 
	.D(n5113), 
	.C(n5155), 
	.B(n5134), 
	.A(n5176));
   MUX4EHD U6629 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5177), 
	.D(\ram[255][6] ), 
	.C(\ram[253][6] ), 
	.B(\ram[254][6] ), 
	.A(\ram[252][6] ));
   MUX4EHD U6630 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5178), 
	.D(\ram[251][6] ), 
	.C(\ram[249][6] ), 
	.B(\ram[250][6] ), 
	.A(\ram[248][6] ));
   MUX4EHD U6631 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5179), 
	.D(\ram[247][6] ), 
	.C(\ram[245][6] ), 
	.B(\ram[246][6] ), 
	.A(\ram[244][6] ));
   MUX4EHD U6632 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5180), 
	.D(\ram[243][6] ), 
	.C(\ram[241][6] ), 
	.B(\ram[242][6] ), 
	.A(\ram[240][6] ));
   MUX4EHD U6633 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5181), 
	.D(n5177), 
	.C(n5179), 
	.B(n5178), 
	.A(n5180));
   MUX4EHD U6634 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5182), 
	.D(\ram[239][6] ), 
	.C(\ram[237][6] ), 
	.B(\ram[238][6] ), 
	.A(\ram[236][6] ));
   MUX4EHD U6635 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5183), 
	.D(\ram[235][6] ), 
	.C(\ram[233][6] ), 
	.B(\ram[234][6] ), 
	.A(\ram[232][6] ));
   MUX4EHD U6636 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5184), 
	.D(\ram[231][6] ), 
	.C(\ram[229][6] ), 
	.B(\ram[230][6] ), 
	.A(\ram[228][6] ));
   MUX4EHD U6637 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5185), 
	.D(\ram[227][6] ), 
	.C(\ram[225][6] ), 
	.B(\ram[226][6] ), 
	.A(\ram[224][6] ));
   MUX4EHD U6638 (.S1(n6136), 
	.S0(n7442), 
	.O(n5186), 
	.D(n5182), 
	.C(n5184), 
	.B(n5183), 
	.A(n5185));
   MUX4EHD U6639 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5187), 
	.D(\ram[223][6] ), 
	.C(\ram[221][6] ), 
	.B(\ram[222][6] ), 
	.A(\ram[220][6] ));
   MUX4EHD U6640 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5188), 
	.D(\ram[219][6] ), 
	.C(\ram[217][6] ), 
	.B(\ram[218][6] ), 
	.A(\ram[216][6] ));
   MUX4EHD U6641 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5189), 
	.D(\ram[215][6] ), 
	.C(\ram[213][6] ), 
	.B(\ram[214][6] ), 
	.A(\ram[212][6] ));
   MUX4EHD U6642 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5190), 
	.D(\ram[211][6] ), 
	.C(\ram[209][6] ), 
	.B(\ram[210][6] ), 
	.A(\ram[208][6] ));
   MUX4EHD U6643 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5191), 
	.D(n5187), 
	.C(n5189), 
	.B(n5188), 
	.A(n5190));
   MUX4EHD U6644 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5192), 
	.D(\ram[207][6] ), 
	.C(\ram[205][6] ), 
	.B(\ram[206][6] ), 
	.A(\ram[204][6] ));
   MUX4EHD U6645 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5193), 
	.D(\ram[203][6] ), 
	.C(\ram[201][6] ), 
	.B(\ram[202][6] ), 
	.A(\ram[200][6] ));
   MUX4EHD U6646 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5194), 
	.D(\ram[199][6] ), 
	.C(\ram[197][6] ), 
	.B(\ram[198][6] ), 
	.A(\ram[196][6] ));
   MUX4EHD U6647 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5195), 
	.D(\ram[195][6] ), 
	.C(\ram[193][6] ), 
	.B(\ram[194][6] ), 
	.A(\ram[192][6] ));
   MUX4EHD U6648 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5196), 
	.D(n5192), 
	.C(n5194), 
	.B(n5193), 
	.A(n5195));
   MUX4EHD U6649 (.S1(n6038), 
	.S0(n7444), 
	.O(n5197), 
	.D(n5181), 
	.C(n5191), 
	.B(n5186), 
	.A(n5196));
   MUX4EHD U6650 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5198), 
	.D(\ram[191][6] ), 
	.C(\ram[189][6] ), 
	.B(\ram[190][6] ), 
	.A(\ram[188][6] ));
   MUX4EHD U6651 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5199), 
	.D(\ram[187][6] ), 
	.C(\ram[185][6] ), 
	.B(\ram[186][6] ), 
	.A(\ram[184][6] ));
   MUX4EHD U6652 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5200), 
	.D(\ram[183][6] ), 
	.C(\ram[181][6] ), 
	.B(\ram[182][6] ), 
	.A(\ram[180][6] ));
   MUX4EHD U6653 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5201), 
	.D(\ram[179][6] ), 
	.C(\ram[177][6] ), 
	.B(\ram[178][6] ), 
	.A(\ram[176][6] ));
   MUX4EHD U6654 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5202), 
	.D(n5198), 
	.C(n5200), 
	.B(n5199), 
	.A(n5201));
   MUX4EHD U6655 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5203), 
	.D(\ram[175][6] ), 
	.C(\ram[173][6] ), 
	.B(\ram[174][6] ), 
	.A(\ram[172][6] ));
   MUX4EHD U6656 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5204), 
	.D(\ram[171][6] ), 
	.C(\ram[169][6] ), 
	.B(\ram[170][6] ), 
	.A(\ram[168][6] ));
   MUX4EHD U6657 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5205), 
	.D(\ram[167][6] ), 
	.C(\ram[165][6] ), 
	.B(\ram[166][6] ), 
	.A(\ram[164][6] ));
   MUX4EHD U6658 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5206), 
	.D(\ram[163][6] ), 
	.C(\ram[161][6] ), 
	.B(\ram[162][6] ), 
	.A(\ram[160][6] ));
   MUX4EHD U6659 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5207), 
	.D(n5203), 
	.C(n5205), 
	.B(n5204), 
	.A(n5206));
   MUX4EHD U6660 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5208), 
	.D(\ram[159][6] ), 
	.C(\ram[157][6] ), 
	.B(\ram[158][6] ), 
	.A(\ram[156][6] ));
   MUX4EHD U6661 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5209), 
	.D(\ram[155][6] ), 
	.C(\ram[153][6] ), 
	.B(\ram[154][6] ), 
	.A(\ram[152][6] ));
   MUX4EHD U6662 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5210), 
	.D(\ram[151][6] ), 
	.C(\ram[149][6] ), 
	.B(\ram[150][6] ), 
	.A(\ram[148][6] ));
   MUX4EHD U6663 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5211), 
	.D(\ram[147][6] ), 
	.C(\ram[145][6] ), 
	.B(\ram[146][6] ), 
	.A(\ram[144][6] ));
   MUX4EHD U6664 (.S1(n6136), 
	.S0(n7442), 
	.O(n5212), 
	.D(n5208), 
	.C(n5210), 
	.B(n5209), 
	.A(n5211));
   MUX4EHD U6665 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5213), 
	.D(\ram[143][6] ), 
	.C(\ram[141][6] ), 
	.B(\ram[142][6] ), 
	.A(\ram[140][6] ));
   MUX4EHD U6666 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5214), 
	.D(\ram[139][6] ), 
	.C(\ram[137][6] ), 
	.B(\ram[138][6] ), 
	.A(\ram[136][6] ));
   MUX4EHD U6667 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5215), 
	.D(\ram[135][6] ), 
	.C(\ram[133][6] ), 
	.B(\ram[134][6] ), 
	.A(\ram[132][6] ));
   MUX4EHD U6668 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5216), 
	.D(\ram[131][6] ), 
	.C(\ram[129][6] ), 
	.B(\ram[130][6] ), 
	.A(\ram[128][6] ));
   MUX4EHD U6669 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5217), 
	.D(n5213), 
	.C(n5215), 
	.B(n5214), 
	.A(n5216));
   MUX4EHD U6670 (.S1(n6038), 
	.S0(n7444), 
	.O(n5218), 
	.D(n5202), 
	.C(n5212), 
	.B(n5207), 
	.A(n5217));
   MUX4EHD U6671 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5219), 
	.D(\ram[127][6] ), 
	.C(\ram[125][6] ), 
	.B(\ram[126][6] ), 
	.A(\ram[124][6] ));
   MUX4EHD U6672 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5220), 
	.D(\ram[123][6] ), 
	.C(\ram[121][6] ), 
	.B(\ram[122][6] ), 
	.A(\ram[120][6] ));
   MUX4EHD U6673 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5221), 
	.D(\ram[119][6] ), 
	.C(\ram[117][6] ), 
	.B(\ram[118][6] ), 
	.A(\ram[116][6] ));
   MUX4EHD U6674 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5222), 
	.D(\ram[115][6] ), 
	.C(\ram[113][6] ), 
	.B(\ram[114][6] ), 
	.A(\ram[112][6] ));
   MUX4EHD U6675 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5223), 
	.D(n5219), 
	.C(n5221), 
	.B(n5220), 
	.A(n5222));
   MUX4EHD U6676 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5224), 
	.D(\ram[111][6] ), 
	.C(\ram[109][6] ), 
	.B(\ram[110][6] ), 
	.A(\ram[108][6] ));
   MUX4EHD U6677 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5225), 
	.D(\ram[107][6] ), 
	.C(\ram[105][6] ), 
	.B(\ram[106][6] ), 
	.A(\ram[104][6] ));
   MUX4EHD U6678 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5226), 
	.D(\ram[103][6] ), 
	.C(\ram[101][6] ), 
	.B(\ram[102][6] ), 
	.A(\ram[100][6] ));
   MUX4EHD U6679 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5227), 
	.D(\ram[99][6] ), 
	.C(\ram[97][6] ), 
	.B(\ram[98][6] ), 
	.A(\ram[96][6] ));
   MUX4EHD U6680 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5228), 
	.D(n5224), 
	.C(n5226), 
	.B(n5225), 
	.A(n5227));
   MUX4EHD U6681 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5229), 
	.D(\ram[95][6] ), 
	.C(\ram[93][6] ), 
	.B(\ram[94][6] ), 
	.A(\ram[92][6] ));
   MUX4EHD U6682 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5230), 
	.D(\ram[91][6] ), 
	.C(\ram[89][6] ), 
	.B(\ram[90][6] ), 
	.A(\ram[88][6] ));
   MUX4EHD U6683 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5231), 
	.D(\ram[87][6] ), 
	.C(\ram[85][6] ), 
	.B(\ram[86][6] ), 
	.A(\ram[84][6] ));
   MUX4EHD U6684 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5232), 
	.D(\ram[83][6] ), 
	.C(\ram[81][6] ), 
	.B(\ram[82][6] ), 
	.A(\ram[80][6] ));
   MUX4EHD U6685 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5233), 
	.D(n5229), 
	.C(n5231), 
	.B(n5230), 
	.A(n5232));
   MUX4EHD U6686 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5234), 
	.D(\ram[79][6] ), 
	.C(\ram[77][6] ), 
	.B(\ram[78][6] ), 
	.A(\ram[76][6] ));
   MUX4EHD U6687 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5235), 
	.D(\ram[75][6] ), 
	.C(\ram[73][6] ), 
	.B(\ram[74][6] ), 
	.A(\ram[72][6] ));
   MUX4EHD U6688 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5236), 
	.D(\ram[71][6] ), 
	.C(\ram[69][6] ), 
	.B(\ram[70][6] ), 
	.A(\ram[68][6] ));
   MUX4EHD U6689 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5237), 
	.D(\ram[67][6] ), 
	.C(\ram[65][6] ), 
	.B(\ram[66][6] ), 
	.A(\ram[64][6] ));
   MUX4EHD U6690 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5238), 
	.D(n5234), 
	.C(n5236), 
	.B(n5235), 
	.A(n5237));
   MUX4EHD U6691 (.S1(n6038), 
	.S0(n7444), 
	.O(n5239), 
	.D(n5223), 
	.C(n5233), 
	.B(n5228), 
	.A(n5238));
   MUX4EHD U6692 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5240), 
	.D(\ram[63][6] ), 
	.C(\ram[61][6] ), 
	.B(\ram[62][6] ), 
	.A(\ram[60][6] ));
   MUX4EHD U6693 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5241), 
	.D(\ram[59][6] ), 
	.C(\ram[57][6] ), 
	.B(\ram[58][6] ), 
	.A(\ram[56][6] ));
   MUX4EHD U6694 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5242), 
	.D(\ram[55][6] ), 
	.C(\ram[53][6] ), 
	.B(\ram[54][6] ), 
	.A(\ram[52][6] ));
   MUX4EHD U6695 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5243), 
	.D(\ram[51][6] ), 
	.C(\ram[49][6] ), 
	.B(\ram[50][6] ), 
	.A(\ram[48][6] ));
   MUX4EHD U6696 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5244), 
	.D(n5240), 
	.C(n5242), 
	.B(n5241), 
	.A(n5243));
   MUX4EHD U6697 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5245), 
	.D(\ram[47][6] ), 
	.C(\ram[45][6] ), 
	.B(\ram[46][6] ), 
	.A(\ram[44][6] ));
   MUX4EHD U6698 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5246), 
	.D(\ram[43][6] ), 
	.C(\ram[41][6] ), 
	.B(\ram[42][6] ), 
	.A(\ram[40][6] ));
   MUX4EHD U6699 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5247), 
	.D(\ram[39][6] ), 
	.C(\ram[37][6] ), 
	.B(\ram[38][6] ), 
	.A(\ram[36][6] ));
   MUX4EHD U6700 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5248), 
	.D(\ram[35][6] ), 
	.C(\ram[33][6] ), 
	.B(\ram[34][6] ), 
	.A(\ram[32][6] ));
   MUX4EHD U6701 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5249), 
	.D(n5245), 
	.C(n5247), 
	.B(n5246), 
	.A(n5248));
   MUX4EHD U6702 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5250), 
	.D(\ram[31][6] ), 
	.C(\ram[29][6] ), 
	.B(\ram[30][6] ), 
	.A(\ram[28][6] ));
   MUX4EHD U6703 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5251), 
	.D(\ram[27][6] ), 
	.C(\ram[25][6] ), 
	.B(\ram[26][6] ), 
	.A(\ram[24][6] ));
   MUX4EHD U6704 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5252), 
	.D(\ram[23][6] ), 
	.C(\ram[21][6] ), 
	.B(\ram[22][6] ), 
	.A(\ram[20][6] ));
   MUX4EHD U6705 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5253), 
	.D(\ram[19][6] ), 
	.C(\ram[17][6] ), 
	.B(\ram[18][6] ), 
	.A(\ram[16][6] ));
   MUX4EHD U6706 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5254), 
	.D(n5250), 
	.C(n5252), 
	.B(n5251), 
	.A(n5253));
   MUX4EHD U6707 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5255), 
	.D(\ram[15][6] ), 
	.C(\ram[13][6] ), 
	.B(\ram[14][6] ), 
	.A(\ram[12][6] ));
   MUX4EHD U6708 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5256), 
	.D(\ram[11][6] ), 
	.C(\ram[9][6] ), 
	.B(\ram[10][6] ), 
	.A(\ram[8][6] ));
   MUX4EHD U6709 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5257), 
	.D(\ram[7][6] ), 
	.C(\ram[5][6] ), 
	.B(\ram[6][6] ), 
	.A(\ram[4][6] ));
   MUX4EHD U6710 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5258), 
	.D(\ram[3][6] ), 
	.C(\ram[1][6] ), 
	.B(\ram[2][6] ), 
	.A(\ram[0][6] ));
   MUX4EHD U6711 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5259), 
	.D(n5255), 
	.C(n5257), 
	.B(n5256), 
	.A(n5258));
   MUX4EHD U6712 (.S1(n6038), 
	.S0(n7444), 
	.O(n5260), 
	.D(n5244), 
	.C(n5254), 
	.B(n5249), 
	.A(n5259));
   MUX4EHD U6713 (.S1(n6469), 
	.S0(n6470), 
	.O(N4135), 
	.D(n5197), 
	.C(n5239), 
	.B(n5218), 
	.A(n5260));
   MUX4EHD U6714 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5261), 
	.D(\ram[255][7] ), 
	.C(\ram[253][7] ), 
	.B(\ram[254][7] ), 
	.A(\ram[252][7] ));
   MUX4EHD U6715 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5262), 
	.D(\ram[251][7] ), 
	.C(\ram[249][7] ), 
	.B(\ram[250][7] ), 
	.A(\ram[248][7] ));
   MUX4EHD U6716 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5263), 
	.D(\ram[247][7] ), 
	.C(\ram[245][7] ), 
	.B(\ram[246][7] ), 
	.A(\ram[244][7] ));
   MUX4EHD U6717 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5264), 
	.D(\ram[243][7] ), 
	.C(\ram[241][7] ), 
	.B(\ram[242][7] ), 
	.A(\ram[240][7] ));
   MUX4EHD U6718 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5265), 
	.D(n5261), 
	.C(n5263), 
	.B(n5262), 
	.A(n5264));
   MUX4EHD U6719 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5266), 
	.D(\ram[239][7] ), 
	.C(\ram[237][7] ), 
	.B(\ram[238][7] ), 
	.A(\ram[236][7] ));
   MUX4EHD U6720 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5267), 
	.D(\ram[235][7] ), 
	.C(\ram[233][7] ), 
	.B(\ram[234][7] ), 
	.A(\ram[232][7] ));
   MUX4EHD U6721 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5268), 
	.D(\ram[231][7] ), 
	.C(\ram[229][7] ), 
	.B(\ram[230][7] ), 
	.A(\ram[228][7] ));
   MUX4EHD U6722 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5269), 
	.D(\ram[227][7] ), 
	.C(\ram[225][7] ), 
	.B(\ram[226][7] ), 
	.A(\ram[224][7] ));
   MUX4EHD U6723 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5270), 
	.D(n5266), 
	.C(n5268), 
	.B(n5267), 
	.A(n5269));
   MUX4EHD U6724 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5271), 
	.D(\ram[223][7] ), 
	.C(\ram[221][7] ), 
	.B(\ram[222][7] ), 
	.A(\ram[220][7] ));
   MUX4EHD U6725 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5272), 
	.D(\ram[219][7] ), 
	.C(\ram[217][7] ), 
	.B(\ram[218][7] ), 
	.A(\ram[216][7] ));
   MUX4EHD U6726 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5273), 
	.D(\ram[215][7] ), 
	.C(\ram[213][7] ), 
	.B(\ram[214][7] ), 
	.A(\ram[212][7] ));
   MUX4EHD U6727 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5274), 
	.D(\ram[211][7] ), 
	.C(\ram[209][7] ), 
	.B(\ram[210][7] ), 
	.A(\ram[208][7] ));
   MUX4EHD U6728 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5275), 
	.D(n5271), 
	.C(n5273), 
	.B(n5272), 
	.A(n5274));
   MUX4EHD U6729 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5276), 
	.D(\ram[207][7] ), 
	.C(\ram[205][7] ), 
	.B(\ram[206][7] ), 
	.A(\ram[204][7] ));
   MUX4EHD U6730 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5277), 
	.D(\ram[203][7] ), 
	.C(\ram[201][7] ), 
	.B(\ram[202][7] ), 
	.A(\ram[200][7] ));
   MUX4EHD U6731 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5278), 
	.D(\ram[199][7] ), 
	.C(\ram[197][7] ), 
	.B(\ram[198][7] ), 
	.A(\ram[196][7] ));
   MUX4EHD U6732 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5279), 
	.D(\ram[195][7] ), 
	.C(\ram[193][7] ), 
	.B(\ram[194][7] ), 
	.A(\ram[192][7] ));
   MUX4EHD U6733 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5280), 
	.D(n5276), 
	.C(n5278), 
	.B(n5277), 
	.A(n5279));
   MUX4EHD U6734 (.S1(n6038), 
	.S0(n7444), 
	.O(n5281), 
	.D(n5265), 
	.C(n5275), 
	.B(n5270), 
	.A(n5280));
   MUX4EHD U6735 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5282), 
	.D(\ram[191][7] ), 
	.C(\ram[189][7] ), 
	.B(\ram[190][7] ), 
	.A(\ram[188][7] ));
   MUX4EHD U6736 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5283), 
	.D(\ram[187][7] ), 
	.C(\ram[185][7] ), 
	.B(\ram[186][7] ), 
	.A(\ram[184][7] ));
   MUX4EHD U6737 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5284), 
	.D(\ram[183][7] ), 
	.C(\ram[181][7] ), 
	.B(\ram[182][7] ), 
	.A(\ram[180][7] ));
   MUX4EHD U6738 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5285), 
	.D(\ram[179][7] ), 
	.C(\ram[177][7] ), 
	.B(\ram[178][7] ), 
	.A(\ram[176][7] ));
   MUX4EHD U6739 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5286), 
	.D(n5282), 
	.C(n5284), 
	.B(n5283), 
	.A(n5285));
   MUX4EHD U6740 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5287), 
	.D(\ram[175][7] ), 
	.C(\ram[173][7] ), 
	.B(\ram[174][7] ), 
	.A(\ram[172][7] ));
   MUX4EHD U6741 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5288), 
	.D(\ram[171][7] ), 
	.C(\ram[169][7] ), 
	.B(\ram[170][7] ), 
	.A(\ram[168][7] ));
   MUX4EHD U6742 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5289), 
	.D(\ram[167][7] ), 
	.C(\ram[165][7] ), 
	.B(\ram[166][7] ), 
	.A(\ram[164][7] ));
   MUX4EHD U6743 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5290), 
	.D(\ram[163][7] ), 
	.C(\ram[161][7] ), 
	.B(\ram[162][7] ), 
	.A(\ram[160][7] ));
   MUX4EHD U6744 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5291), 
	.D(n5287), 
	.C(n5289), 
	.B(n5288), 
	.A(n5290));
   MUX4EHD U6745 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5292), 
	.D(\ram[159][7] ), 
	.C(\ram[157][7] ), 
	.B(\ram[158][7] ), 
	.A(\ram[156][7] ));
   MUX4EHD U6746 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n5293), 
	.D(\ram[155][7] ), 
	.C(\ram[153][7] ), 
	.B(\ram[154][7] ), 
	.A(\ram[152][7] ));
   MUX4EHD U6747 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5294), 
	.D(\ram[151][7] ), 
	.C(\ram[149][7] ), 
	.B(\ram[150][7] ), 
	.A(\ram[148][7] ));
   MUX4EHD U6748 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5295), 
	.D(\ram[147][7] ), 
	.C(\ram[145][7] ), 
	.B(\ram[146][7] ), 
	.A(\ram[144][7] ));
   MUX4EHD U6749 (.S1(n6136), 
	.S0(n7442), 
	.O(n5296), 
	.D(n5292), 
	.C(n5294), 
	.B(n5293), 
	.A(n5295));
   MUX4EHD U6750 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5297), 
	.D(\ram[143][7] ), 
	.C(\ram[141][7] ), 
	.B(\ram[142][7] ), 
	.A(\ram[140][7] ));
   MUX4EHD U6751 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5298), 
	.D(\ram[139][7] ), 
	.C(\ram[137][7] ), 
	.B(\ram[138][7] ), 
	.A(\ram[136][7] ));
   MUX4EHD U6752 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5299), 
	.D(\ram[135][7] ), 
	.C(\ram[133][7] ), 
	.B(\ram[134][7] ), 
	.A(\ram[132][7] ));
   MUX4EHD U6753 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5300), 
	.D(\ram[131][7] ), 
	.C(\ram[129][7] ), 
	.B(\ram[130][7] ), 
	.A(\ram[128][7] ));
   MUX4EHD U6754 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5301), 
	.D(n5297), 
	.C(n5299), 
	.B(n5298), 
	.A(n5300));
   MUX4EHD U6755 (.S1(n6038), 
	.S0(n7444), 
	.O(n5302), 
	.D(n5286), 
	.C(n5296), 
	.B(n5291), 
	.A(n5301));
   MUX4EHD U6756 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5303), 
	.D(\ram[127][7] ), 
	.C(\ram[125][7] ), 
	.B(\ram[126][7] ), 
	.A(\ram[124][7] ));
   MUX4EHD U6757 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5304), 
	.D(\ram[123][7] ), 
	.C(\ram[121][7] ), 
	.B(\ram[122][7] ), 
	.A(\ram[120][7] ));
   MUX4EHD U6758 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5305), 
	.D(\ram[119][7] ), 
	.C(\ram[117][7] ), 
	.B(\ram[118][7] ), 
	.A(\ram[116][7] ));
   MUX4EHD U6759 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5306), 
	.D(\ram[115][7] ), 
	.C(\ram[113][7] ), 
	.B(\ram[114][7] ), 
	.A(\ram[112][7] ));
   MUX4EHD U6760 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5307), 
	.D(n5303), 
	.C(n5305), 
	.B(n5304), 
	.A(n5306));
   MUX4EHD U6761 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5308), 
	.D(\ram[111][7] ), 
	.C(\ram[109][7] ), 
	.B(\ram[110][7] ), 
	.A(\ram[108][7] ));
   MUX4EHD U6762 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5309), 
	.D(\ram[107][7] ), 
	.C(\ram[105][7] ), 
	.B(\ram[106][7] ), 
	.A(\ram[104][7] ));
   MUX4EHD U6763 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5310), 
	.D(\ram[103][7] ), 
	.C(\ram[101][7] ), 
	.B(\ram[102][7] ), 
	.A(\ram[100][7] ));
   MUX4EHD U6764 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5311), 
	.D(\ram[99][7] ), 
	.C(\ram[97][7] ), 
	.B(\ram[98][7] ), 
	.A(\ram[96][7] ));
   MUX4EHD U6765 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5312), 
	.D(n5308), 
	.C(n5310), 
	.B(n5309), 
	.A(n5311));
   MUX4EHD U6766 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5313), 
	.D(\ram[95][7] ), 
	.C(\ram[93][7] ), 
	.B(\ram[94][7] ), 
	.A(\ram[92][7] ));
   MUX4EHD U6767 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5314), 
	.D(\ram[91][7] ), 
	.C(\ram[89][7] ), 
	.B(\ram[90][7] ), 
	.A(\ram[88][7] ));
   MUX4EHD U6768 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5315), 
	.D(\ram[87][7] ), 
	.C(\ram[85][7] ), 
	.B(\ram[86][7] ), 
	.A(\ram[84][7] ));
   MUX4EHD U6769 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5316), 
	.D(\ram[83][7] ), 
	.C(\ram[81][7] ), 
	.B(\ram[82][7] ), 
	.A(\ram[80][7] ));
   MUX4EHD U6770 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5317), 
	.D(n5313), 
	.C(n5315), 
	.B(n5314), 
	.A(n5316));
   MUX4EHD U6771 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5318), 
	.D(\ram[79][7] ), 
	.C(\ram[77][7] ), 
	.B(\ram[78][7] ), 
	.A(\ram[76][7] ));
   MUX4EHD U6772 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5319), 
	.D(\ram[75][7] ), 
	.C(\ram[73][7] ), 
	.B(\ram[74][7] ), 
	.A(\ram[72][7] ));
   MUX4EHD U6773 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5320), 
	.D(\ram[71][7] ), 
	.C(\ram[69][7] ), 
	.B(\ram[70][7] ), 
	.A(\ram[68][7] ));
   MUX4EHD U6774 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5321), 
	.D(\ram[67][7] ), 
	.C(\ram[65][7] ), 
	.B(\ram[66][7] ), 
	.A(\ram[64][7] ));
   MUX4EHD U6775 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5322), 
	.D(n5318), 
	.C(n5320), 
	.B(n5319), 
	.A(n5321));
   MUX4EHD U6776 (.S1(n6038), 
	.S0(n7444), 
	.O(n5323), 
	.D(n5307), 
	.C(n5317), 
	.B(n5312), 
	.A(n5322));
   MUX4EHD U6777 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5324), 
	.D(\ram[63][7] ), 
	.C(\ram[61][7] ), 
	.B(\ram[62][7] ), 
	.A(\ram[60][7] ));
   MUX4EHD U6778 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5325), 
	.D(\ram[59][7] ), 
	.C(\ram[57][7] ), 
	.B(\ram[58][7] ), 
	.A(\ram[56][7] ));
   MUX4EHD U6779 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5326), 
	.D(\ram[55][7] ), 
	.C(\ram[53][7] ), 
	.B(\ram[54][7] ), 
	.A(\ram[52][7] ));
   MUX4EHD U6780 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5327), 
	.D(\ram[51][7] ), 
	.C(\ram[49][7] ), 
	.B(\ram[50][7] ), 
	.A(\ram[48][7] ));
   MUX4EHD U6781 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5328), 
	.D(n5324), 
	.C(n5326), 
	.B(n5325), 
	.A(n5327));
   MUX4EHD U6782 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5329), 
	.D(\ram[47][7] ), 
	.C(\ram[45][7] ), 
	.B(\ram[46][7] ), 
	.A(\ram[44][7] ));
   MUX4EHD U6783 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5330), 
	.D(\ram[43][7] ), 
	.C(\ram[41][7] ), 
	.B(\ram[42][7] ), 
	.A(\ram[40][7] ));
   MUX4EHD U6784 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5331), 
	.D(\ram[39][7] ), 
	.C(\ram[37][7] ), 
	.B(\ram[38][7] ), 
	.A(\ram[36][7] ));
   MUX4EHD U6785 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5332), 
	.D(\ram[35][7] ), 
	.C(\ram[33][7] ), 
	.B(\ram[34][7] ), 
	.A(\ram[32][7] ));
   MUX4EHD U6786 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5333), 
	.D(n5329), 
	.C(n5331), 
	.B(n5330), 
	.A(n5332));
   MUX4EHD U6787 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5334), 
	.D(\ram[31][7] ), 
	.C(\ram[29][7] ), 
	.B(\ram[30][7] ), 
	.A(\ram[28][7] ));
   MUX4EHD U6788 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5335), 
	.D(\ram[27][7] ), 
	.C(\ram[25][7] ), 
	.B(\ram[26][7] ), 
	.A(\ram[24][7] ));
   MUX4EHD U6789 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5336), 
	.D(\ram[23][7] ), 
	.C(\ram[21][7] ), 
	.B(\ram[22][7] ), 
	.A(\ram[20][7] ));
   MUX4EHD U6790 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5337), 
	.D(\ram[19][7] ), 
	.C(\ram[17][7] ), 
	.B(\ram[18][7] ), 
	.A(\ram[16][7] ));
   MUX4EHD U6791 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5338), 
	.D(n5334), 
	.C(n5336), 
	.B(n5335), 
	.A(n5337));
   MUX4EHD U6792 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5339), 
	.D(\ram[15][7] ), 
	.C(\ram[13][7] ), 
	.B(\ram[14][7] ), 
	.A(\ram[12][7] ));
   MUX4EHD U6793 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5340), 
	.D(\ram[11][7] ), 
	.C(\ram[9][7] ), 
	.B(\ram[10][7] ), 
	.A(\ram[8][7] ));
   MUX4EHD U6794 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5341), 
	.D(\ram[7][7] ), 
	.C(\ram[5][7] ), 
	.B(\ram[6][7] ), 
	.A(\ram[4][7] ));
   MUX4EHD U6795 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5342), 
	.D(\ram[3][7] ), 
	.C(\ram[1][7] ), 
	.B(\ram[2][7] ), 
	.A(\ram[0][7] ));
   MUX4EHD U6796 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5343), 
	.D(n5339), 
	.C(n5341), 
	.B(n5340), 
	.A(n5342));
   MUX4EHD U6797 (.S1(n6038), 
	.S0(n7444), 
	.O(n5344), 
	.D(n5328), 
	.C(n5338), 
	.B(n5333), 
	.A(n5343));
   MUX4EHD U6798 (.S1(n6469), 
	.S0(n6470), 
	.O(N4134), 
	.D(n5281), 
	.C(n5323), 
	.B(n5302), 
	.A(n5344));
   MUX4EHD U6799 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5345), 
	.D(\ram[255][8] ), 
	.C(\ram[253][8] ), 
	.B(\ram[254][8] ), 
	.A(\ram[252][8] ));
   MUX4EHD U6800 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5346), 
	.D(\ram[251][8] ), 
	.C(\ram[249][8] ), 
	.B(\ram[250][8] ), 
	.A(\ram[248][8] ));
   MUX4EHD U6801 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5347), 
	.D(\ram[247][8] ), 
	.C(\ram[245][8] ), 
	.B(\ram[246][8] ), 
	.A(\ram[244][8] ));
   MUX4EHD U6802 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5348), 
	.D(\ram[243][8] ), 
	.C(\ram[241][8] ), 
	.B(\ram[242][8] ), 
	.A(\ram[240][8] ));
   MUX4EHD U6803 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5349), 
	.D(n5345), 
	.C(n5347), 
	.B(n5346), 
	.A(n5348));
   MUX4EHD U6804 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5350), 
	.D(\ram[239][8] ), 
	.C(\ram[237][8] ), 
	.B(\ram[238][8] ), 
	.A(\ram[236][8] ));
   MUX4EHD U6805 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5351), 
	.D(\ram[235][8] ), 
	.C(\ram[233][8] ), 
	.B(\ram[234][8] ), 
	.A(\ram[232][8] ));
   MUX4EHD U6806 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5352), 
	.D(\ram[231][8] ), 
	.C(\ram[229][8] ), 
	.B(\ram[230][8] ), 
	.A(\ram[228][8] ));
   MUX4EHD U6807 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5353), 
	.D(\ram[227][8] ), 
	.C(\ram[225][8] ), 
	.B(\ram[226][8] ), 
	.A(\ram[224][8] ));
   MUX4EHD U6808 (.S1(n6136), 
	.S0(n7442), 
	.O(n5354), 
	.D(n5350), 
	.C(n5352), 
	.B(n5351), 
	.A(n5353));
   MUX4EHD U6809 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5355), 
	.D(\ram[223][8] ), 
	.C(\ram[221][8] ), 
	.B(\ram[222][8] ), 
	.A(\ram[220][8] ));
   MUX4EHD U6810 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5356), 
	.D(\ram[219][8] ), 
	.C(\ram[217][8] ), 
	.B(\ram[218][8] ), 
	.A(\ram[216][8] ));
   MUX4EHD U6811 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5357), 
	.D(\ram[215][8] ), 
	.C(\ram[213][8] ), 
	.B(\ram[214][8] ), 
	.A(\ram[212][8] ));
   MUX4EHD U6812 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5358), 
	.D(\ram[211][8] ), 
	.C(\ram[209][8] ), 
	.B(\ram[210][8] ), 
	.A(\ram[208][8] ));
   MUX4EHD U6813 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5359), 
	.D(n5355), 
	.C(n5357), 
	.B(n5356), 
	.A(n5358));
   MUX4EHD U6814 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5360), 
	.D(\ram[207][8] ), 
	.C(\ram[205][8] ), 
	.B(\ram[206][8] ), 
	.A(\ram[204][8] ));
   MUX4EHD U6815 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5361), 
	.D(\ram[203][8] ), 
	.C(\ram[201][8] ), 
	.B(\ram[202][8] ), 
	.A(\ram[200][8] ));
   MUX4EHD U6816 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5362), 
	.D(\ram[199][8] ), 
	.C(\ram[197][8] ), 
	.B(\ram[198][8] ), 
	.A(\ram[196][8] ));
   MUX4EHD U6817 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5363), 
	.D(\ram[195][8] ), 
	.C(\ram[193][8] ), 
	.B(\ram[194][8] ), 
	.A(\ram[192][8] ));
   MUX4EHD U6818 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5364), 
	.D(n5360), 
	.C(n5362), 
	.B(n5361), 
	.A(n5363));
   MUX4EHD U6819 (.S1(n6038), 
	.S0(n7444), 
	.O(n5365), 
	.D(n5349), 
	.C(n5359), 
	.B(n5354), 
	.A(n5364));
   MUX4EHD U6820 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5366), 
	.D(\ram[191][8] ), 
	.C(\ram[189][8] ), 
	.B(\ram[190][8] ), 
	.A(\ram[188][8] ));
   MUX4EHD U6821 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5367), 
	.D(\ram[187][8] ), 
	.C(\ram[185][8] ), 
	.B(\ram[186][8] ), 
	.A(\ram[184][8] ));
   MUX4EHD U6822 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5368), 
	.D(\ram[183][8] ), 
	.C(\ram[181][8] ), 
	.B(\ram[182][8] ), 
	.A(\ram[180][8] ));
   MUX4EHD U6823 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5369), 
	.D(\ram[179][8] ), 
	.C(\ram[177][8] ), 
	.B(\ram[178][8] ), 
	.A(\ram[176][8] ));
   MUX4EHD U6824 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5370), 
	.D(n5366), 
	.C(n5368), 
	.B(n5367), 
	.A(n5369));
   MUX4EHD U6825 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5371), 
	.D(\ram[175][8] ), 
	.C(\ram[173][8] ), 
	.B(\ram[174][8] ), 
	.A(\ram[172][8] ));
   MUX4EHD U6826 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5372), 
	.D(\ram[171][8] ), 
	.C(\ram[169][8] ), 
	.B(\ram[170][8] ), 
	.A(\ram[168][8] ));
   MUX4EHD U6827 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5373), 
	.D(\ram[167][8] ), 
	.C(\ram[165][8] ), 
	.B(\ram[166][8] ), 
	.A(\ram[164][8] ));
   MUX4EHD U6828 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5374), 
	.D(\ram[163][8] ), 
	.C(\ram[161][8] ), 
	.B(\ram[162][8] ), 
	.A(\ram[160][8] ));
   MUX4EHD U6829 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5375), 
	.D(n5371), 
	.C(n5373), 
	.B(n5372), 
	.A(n5374));
   MUX4EHD U6830 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5376), 
	.D(\ram[159][8] ), 
	.C(\ram[157][8] ), 
	.B(\ram[158][8] ), 
	.A(\ram[156][8] ));
   MUX4EHD U6831 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5377), 
	.D(\ram[155][8] ), 
	.C(\ram[153][8] ), 
	.B(\ram[154][8] ), 
	.A(\ram[152][8] ));
   MUX4EHD U6832 (.S1(FE_OFN28_n6459), 
	.S0(n7440), 
	.O(n5378), 
	.D(\ram[151][8] ), 
	.C(\ram[149][8] ), 
	.B(\ram[150][8] ), 
	.A(\ram[148][8] ));
   MUX4EHD U6833 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5379), 
	.D(\ram[147][8] ), 
	.C(\ram[145][8] ), 
	.B(\ram[146][8] ), 
	.A(\ram[144][8] ));
   MUX4EHD U6834 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5380), 
	.D(n5376), 
	.C(n5378), 
	.B(n5377), 
	.A(n5379));
   MUX4EHD U6835 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5381), 
	.D(\ram[143][8] ), 
	.C(\ram[141][8] ), 
	.B(\ram[142][8] ), 
	.A(\ram[140][8] ));
   MUX4EHD U6836 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5382), 
	.D(\ram[139][8] ), 
	.C(\ram[137][8] ), 
	.B(\ram[138][8] ), 
	.A(\ram[136][8] ));
   MUX4EHD U6837 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5383), 
	.D(\ram[135][8] ), 
	.C(\ram[133][8] ), 
	.B(\ram[134][8] ), 
	.A(\ram[132][8] ));
   MUX4EHD U6838 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5384), 
	.D(\ram[131][8] ), 
	.C(\ram[129][8] ), 
	.B(\ram[130][8] ), 
	.A(\ram[128][8] ));
   MUX4EHD U6839 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5385), 
	.D(n5381), 
	.C(n5383), 
	.B(n5382), 
	.A(n5384));
   MUX4EHD U6840 (.S1(n6038), 
	.S0(n7444), 
	.O(n5386), 
	.D(n5370), 
	.C(n5380), 
	.B(n5375), 
	.A(n5385));
   MUX4EHD U6841 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5387), 
	.D(\ram[127][8] ), 
	.C(\ram[125][8] ), 
	.B(\ram[126][8] ), 
	.A(\ram[124][8] ));
   MUX4EHD U6842 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5388), 
	.D(\ram[123][8] ), 
	.C(\ram[121][8] ), 
	.B(\ram[122][8] ), 
	.A(\ram[120][8] ));
   MUX4EHD U6843 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5389), 
	.D(\ram[119][8] ), 
	.C(\ram[117][8] ), 
	.B(\ram[118][8] ), 
	.A(\ram[116][8] ));
   MUX4EHD U6844 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5390), 
	.D(\ram[115][8] ), 
	.C(\ram[113][8] ), 
	.B(\ram[114][8] ), 
	.A(\ram[112][8] ));
   MUX4EHD U6845 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5391), 
	.D(n5387), 
	.C(n5389), 
	.B(n5388), 
	.A(n5390));
   MUX4EHD U6846 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5392), 
	.D(\ram[111][8] ), 
	.C(\ram[109][8] ), 
	.B(\ram[110][8] ), 
	.A(\ram[108][8] ));
   MUX4EHD U6847 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5393), 
	.D(\ram[107][8] ), 
	.C(\ram[105][8] ), 
	.B(\ram[106][8] ), 
	.A(\ram[104][8] ));
   MUX4EHD U6848 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5394), 
	.D(\ram[103][8] ), 
	.C(\ram[101][8] ), 
	.B(\ram[102][8] ), 
	.A(\ram[100][8] ));
   MUX4EHD U6849 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5395), 
	.D(\ram[99][8] ), 
	.C(\ram[97][8] ), 
	.B(\ram[98][8] ), 
	.A(\ram[96][8] ));
   MUX4EHD U6850 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5396), 
	.D(n5392), 
	.C(n5394), 
	.B(n5393), 
	.A(n5395));
   MUX4EHD U6851 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5397), 
	.D(\ram[95][8] ), 
	.C(\ram[93][8] ), 
	.B(\ram[94][8] ), 
	.A(\ram[92][8] ));
   MUX4EHD U6852 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5398), 
	.D(\ram[91][8] ), 
	.C(\ram[89][8] ), 
	.B(\ram[90][8] ), 
	.A(\ram[88][8] ));
   MUX4EHD U6853 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5399), 
	.D(\ram[87][8] ), 
	.C(\ram[85][8] ), 
	.B(\ram[86][8] ), 
	.A(\ram[84][8] ));
   MUX4EHD U6854 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5400), 
	.D(\ram[83][8] ), 
	.C(\ram[81][8] ), 
	.B(\ram[82][8] ), 
	.A(\ram[80][8] ));
   MUX4EHD U6855 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5401), 
	.D(n5397), 
	.C(n5399), 
	.B(n5398), 
	.A(n5400));
   MUX4EHD U6856 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5402), 
	.D(\ram[79][8] ), 
	.C(\ram[77][8] ), 
	.B(\ram[78][8] ), 
	.A(\ram[76][8] ));
   MUX4EHD U6857 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5403), 
	.D(\ram[75][8] ), 
	.C(\ram[73][8] ), 
	.B(\ram[74][8] ), 
	.A(\ram[72][8] ));
   MUX4EHD U6858 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5404), 
	.D(\ram[71][8] ), 
	.C(\ram[69][8] ), 
	.B(\ram[70][8] ), 
	.A(\ram[68][8] ));
   MUX4EHD U6859 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5405), 
	.D(\ram[67][8] ), 
	.C(\ram[65][8] ), 
	.B(\ram[66][8] ), 
	.A(\ram[64][8] ));
   MUX4EHD U6860 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5406), 
	.D(n5402), 
	.C(n5404), 
	.B(n5403), 
	.A(n5405));
   MUX4EHD U6861 (.S1(n6038), 
	.S0(n7444), 
	.O(n5407), 
	.D(n5391), 
	.C(n5401), 
	.B(n5396), 
	.A(n5406));
   MUX4EHD U6862 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5408), 
	.D(\ram[63][8] ), 
	.C(\ram[61][8] ), 
	.B(\ram[62][8] ), 
	.A(\ram[60][8] ));
   MUX4EHD U6863 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5409), 
	.D(\ram[59][8] ), 
	.C(\ram[57][8] ), 
	.B(\ram[58][8] ), 
	.A(\ram[56][8] ));
   MUX4EHD U6864 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5410), 
	.D(\ram[55][8] ), 
	.C(\ram[53][8] ), 
	.B(\ram[54][8] ), 
	.A(\ram[52][8] ));
   MUX4EHD U6865 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5411), 
	.D(\ram[51][8] ), 
	.C(\ram[49][8] ), 
	.B(\ram[50][8] ), 
	.A(\ram[48][8] ));
   MUX4EHD U6866 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5412), 
	.D(n5408), 
	.C(n5410), 
	.B(n5409), 
	.A(n5411));
   MUX4EHD U6867 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5413), 
	.D(\ram[47][8] ), 
	.C(\ram[45][8] ), 
	.B(\ram[46][8] ), 
	.A(\ram[44][8] ));
   MUX4EHD U6868 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5414), 
	.D(\ram[43][8] ), 
	.C(\ram[41][8] ), 
	.B(\ram[42][8] ), 
	.A(\ram[40][8] ));
   MUX4EHD U6869 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5415), 
	.D(\ram[39][8] ), 
	.C(\ram[37][8] ), 
	.B(\ram[38][8] ), 
	.A(\ram[36][8] ));
   MUX4EHD U6870 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5416), 
	.D(\ram[35][8] ), 
	.C(\ram[33][8] ), 
	.B(\ram[34][8] ), 
	.A(\ram[32][8] ));
   MUX4EHD U6871 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5417), 
	.D(n5413), 
	.C(n5415), 
	.B(n5414), 
	.A(n5416));
   MUX4EHD U6872 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5418), 
	.D(\ram[31][8] ), 
	.C(\ram[29][8] ), 
	.B(\ram[30][8] ), 
	.A(\ram[28][8] ));
   MUX4EHD U6873 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5419), 
	.D(\ram[27][8] ), 
	.C(\ram[25][8] ), 
	.B(\ram[26][8] ), 
	.A(\ram[24][8] ));
   MUX4EHD U6874 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5420), 
	.D(\ram[23][8] ), 
	.C(\ram[21][8] ), 
	.B(\ram[22][8] ), 
	.A(\ram[20][8] ));
   MUX4EHD U6875 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5421), 
	.D(\ram[19][8] ), 
	.C(\ram[17][8] ), 
	.B(\ram[18][8] ), 
	.A(\ram[16][8] ));
   MUX4EHD U6876 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5422), 
	.D(n5418), 
	.C(n5420), 
	.B(n5419), 
	.A(n5421));
   MUX4EHD U6877 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5423), 
	.D(\ram[15][8] ), 
	.C(\ram[13][8] ), 
	.B(\ram[14][8] ), 
	.A(\ram[12][8] ));
   MUX4EHD U6878 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5424), 
	.D(\ram[11][8] ), 
	.C(\ram[9][8] ), 
	.B(\ram[10][8] ), 
	.A(\ram[8][8] ));
   MUX4EHD U6879 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5425), 
	.D(\ram[7][8] ), 
	.C(\ram[5][8] ), 
	.B(\ram[6][8] ), 
	.A(\ram[4][8] ));
   MUX4EHD U6880 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n5426), 
	.D(\ram[3][8] ), 
	.C(\ram[1][8] ), 
	.B(\ram[2][8] ), 
	.A(\ram[0][8] ));
   MUX4EHD U6881 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5427), 
	.D(n5423), 
	.C(n5425), 
	.B(n5424), 
	.A(n5426));
   MUX4EHD U6882 (.S1(n6038), 
	.S0(n7444), 
	.O(n5428), 
	.D(n5412), 
	.C(n5422), 
	.B(n5417), 
	.A(n5427));
   MUX4EHD U6883 (.S1(n6469), 
	.S0(n6470), 
	.O(N4133), 
	.D(n5365), 
	.C(n5407), 
	.B(n5386), 
	.A(n5428));
   MUX4EHD U6884 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5429), 
	.D(\ram[255][9] ), 
	.C(\ram[253][9] ), 
	.B(\ram[254][9] ), 
	.A(\ram[252][9] ));
   MUX4EHD U6885 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5430), 
	.D(\ram[251][9] ), 
	.C(\ram[249][9] ), 
	.B(\ram[250][9] ), 
	.A(\ram[248][9] ));
   MUX4EHD U6886 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5431), 
	.D(\ram[247][9] ), 
	.C(\ram[245][9] ), 
	.B(\ram[246][9] ), 
	.A(\ram[244][9] ));
   MUX4EHD U6887 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5432), 
	.D(\ram[243][9] ), 
	.C(\ram[241][9] ), 
	.B(\ram[242][9] ), 
	.A(\ram[240][9] ));
   MUX4EHD U6888 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5433), 
	.D(n5429), 
	.C(n5431), 
	.B(n5430), 
	.A(n5432));
   MUX4EHD U6889 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5434), 
	.D(\ram[239][9] ), 
	.C(\ram[237][9] ), 
	.B(\ram[238][9] ), 
	.A(\ram[236][9] ));
   MUX4EHD U6890 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5435), 
	.D(\ram[235][9] ), 
	.C(\ram[233][9] ), 
	.B(\ram[234][9] ), 
	.A(\ram[232][9] ));
   MUX4EHD U6891 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5436), 
	.D(\ram[231][9] ), 
	.C(\ram[229][9] ), 
	.B(\ram[230][9] ), 
	.A(\ram[228][9] ));
   MUX4EHD U6892 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5437), 
	.D(\ram[227][9] ), 
	.C(\ram[225][9] ), 
	.B(\ram[226][9] ), 
	.A(\ram[224][9] ));
   MUX4EHD U6893 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5438), 
	.D(n5434), 
	.C(n5436), 
	.B(n5435), 
	.A(n5437));
   MUX4EHD U6894 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5439), 
	.D(\ram[223][9] ), 
	.C(\ram[221][9] ), 
	.B(\ram[222][9] ), 
	.A(\ram[220][9] ));
   MUX4EHD U6895 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5440), 
	.D(\ram[219][9] ), 
	.C(\ram[217][9] ), 
	.B(\ram[218][9] ), 
	.A(\ram[216][9] ));
   MUX4EHD U6896 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5441), 
	.D(\ram[215][9] ), 
	.C(\ram[213][9] ), 
	.B(\ram[214][9] ), 
	.A(\ram[212][9] ));
   MUX4EHD U6897 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5442), 
	.D(\ram[211][9] ), 
	.C(\ram[209][9] ), 
	.B(\ram[210][9] ), 
	.A(\ram[208][9] ));
   MUX4EHD U6898 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5443), 
	.D(n5439), 
	.C(n5441), 
	.B(n5440), 
	.A(n5442));
   MUX4EHD U6899 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5444), 
	.D(\ram[207][9] ), 
	.C(\ram[205][9] ), 
	.B(\ram[206][9] ), 
	.A(\ram[204][9] ));
   MUX4EHD U6900 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5445), 
	.D(\ram[203][9] ), 
	.C(\ram[201][9] ), 
	.B(\ram[202][9] ), 
	.A(\ram[200][9] ));
   MUX4EHD U6901 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5446), 
	.D(\ram[199][9] ), 
	.C(\ram[197][9] ), 
	.B(\ram[198][9] ), 
	.A(\ram[196][9] ));
   MUX4EHD U6902 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5447), 
	.D(\ram[195][9] ), 
	.C(\ram[193][9] ), 
	.B(\ram[194][9] ), 
	.A(\ram[192][9] ));
   MUX4EHD U6903 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5448), 
	.D(n5444), 
	.C(n5446), 
	.B(n5445), 
	.A(n5447));
   MUX4EHD U6904 (.S1(n6038), 
	.S0(n7444), 
	.O(n5449), 
	.D(n5433), 
	.C(n5443), 
	.B(n5438), 
	.A(n5448));
   MUX4EHD U6905 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5450), 
	.D(\ram[191][9] ), 
	.C(\ram[189][9] ), 
	.B(\ram[190][9] ), 
	.A(\ram[188][9] ));
   MUX4EHD U6906 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5451), 
	.D(\ram[187][9] ), 
	.C(\ram[185][9] ), 
	.B(\ram[186][9] ), 
	.A(\ram[184][9] ));
   MUX4EHD U6907 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5452), 
	.D(\ram[183][9] ), 
	.C(\ram[181][9] ), 
	.B(\ram[182][9] ), 
	.A(\ram[180][9] ));
   MUX4EHD U6908 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5453), 
	.D(\ram[179][9] ), 
	.C(\ram[177][9] ), 
	.B(\ram[178][9] ), 
	.A(\ram[176][9] ));
   MUX4EHD U6909 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5454), 
	.D(n5450), 
	.C(n5452), 
	.B(n5451), 
	.A(n5453));
   MUX4EHD U6910 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5455), 
	.D(\ram[175][9] ), 
	.C(\ram[173][9] ), 
	.B(\ram[174][9] ), 
	.A(\ram[172][9] ));
   MUX4EHD U6911 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5456), 
	.D(\ram[171][9] ), 
	.C(\ram[169][9] ), 
	.B(\ram[170][9] ), 
	.A(\ram[168][9] ));
   MUX4EHD U6912 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5457), 
	.D(\ram[167][9] ), 
	.C(\ram[165][9] ), 
	.B(\ram[166][9] ), 
	.A(\ram[164][9] ));
   MUX4EHD U6913 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5458), 
	.D(\ram[163][9] ), 
	.C(\ram[161][9] ), 
	.B(\ram[162][9] ), 
	.A(\ram[160][9] ));
   MUX4EHD U6914 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5459), 
	.D(n5455), 
	.C(n5457), 
	.B(n5456), 
	.A(n5458));
   MUX4EHD U6915 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5460), 
	.D(\ram[159][9] ), 
	.C(\ram[157][9] ), 
	.B(\ram[158][9] ), 
	.A(\ram[156][9] ));
   MUX4EHD U6916 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5461), 
	.D(\ram[155][9] ), 
	.C(\ram[153][9] ), 
	.B(\ram[154][9] ), 
	.A(\ram[152][9] ));
   MUX4EHD U6917 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5462), 
	.D(\ram[151][9] ), 
	.C(\ram[149][9] ), 
	.B(\ram[150][9] ), 
	.A(\ram[148][9] ));
   MUX4EHD U6918 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5463), 
	.D(\ram[147][9] ), 
	.C(\ram[145][9] ), 
	.B(\ram[146][9] ), 
	.A(\ram[144][9] ));
   MUX4EHD U6919 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5464), 
	.D(n5460), 
	.C(n5462), 
	.B(n5461), 
	.A(n5463));
   MUX4EHD U6920 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5465), 
	.D(\ram[143][9] ), 
	.C(\ram[141][9] ), 
	.B(\ram[142][9] ), 
	.A(\ram[140][9] ));
   MUX4EHD U6921 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5466), 
	.D(\ram[139][9] ), 
	.C(\ram[137][9] ), 
	.B(\ram[138][9] ), 
	.A(\ram[136][9] ));
   MUX4EHD U6922 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5467), 
	.D(\ram[135][9] ), 
	.C(\ram[133][9] ), 
	.B(\ram[134][9] ), 
	.A(\ram[132][9] ));
   MUX4EHD U6923 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5468), 
	.D(\ram[131][9] ), 
	.C(\ram[129][9] ), 
	.B(\ram[130][9] ), 
	.A(\ram[128][9] ));
   MUX4EHD U6924 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5469), 
	.D(n5465), 
	.C(n5467), 
	.B(n5466), 
	.A(n5468));
   MUX4EHD U6925 (.S1(n6038), 
	.S0(n7444), 
	.O(n5470), 
	.D(n5454), 
	.C(n5464), 
	.B(n5459), 
	.A(n5469));
   MUX4EHD U6926 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5471), 
	.D(\ram[127][9] ), 
	.C(\ram[125][9] ), 
	.B(\ram[126][9] ), 
	.A(\ram[124][9] ));
   MUX4EHD U6927 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5472), 
	.D(\ram[123][9] ), 
	.C(\ram[121][9] ), 
	.B(\ram[122][9] ), 
	.A(\ram[120][9] ));
   MUX4EHD U6928 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5473), 
	.D(\ram[119][9] ), 
	.C(\ram[117][9] ), 
	.B(\ram[118][9] ), 
	.A(\ram[116][9] ));
   MUX4EHD U6929 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5474), 
	.D(\ram[115][9] ), 
	.C(\ram[113][9] ), 
	.B(\ram[114][9] ), 
	.A(\ram[112][9] ));
   MUX4EHD U6930 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5475), 
	.D(n5471), 
	.C(n5473), 
	.B(n5472), 
	.A(n5474));
   MUX4EHD U6931 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5476), 
	.D(\ram[111][9] ), 
	.C(\ram[109][9] ), 
	.B(\ram[110][9] ), 
	.A(\ram[108][9] ));
   MUX4EHD U6932 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5477), 
	.D(\ram[107][9] ), 
	.C(\ram[105][9] ), 
	.B(\ram[106][9] ), 
	.A(\ram[104][9] ));
   MUX4EHD U6933 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5478), 
	.D(\ram[103][9] ), 
	.C(\ram[101][9] ), 
	.B(\ram[102][9] ), 
	.A(\ram[100][9] ));
   MUX4EHD U6934 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5479), 
	.D(\ram[99][9] ), 
	.C(\ram[97][9] ), 
	.B(\ram[98][9] ), 
	.A(\ram[96][9] ));
   MUX4EHD U6935 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5480), 
	.D(n5476), 
	.C(n5478), 
	.B(n5477), 
	.A(n5479));
   MUX4EHD U6936 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5481), 
	.D(\ram[95][9] ), 
	.C(\ram[93][9] ), 
	.B(\ram[94][9] ), 
	.A(\ram[92][9] ));
   MUX4EHD U6937 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5482), 
	.D(\ram[91][9] ), 
	.C(\ram[89][9] ), 
	.B(\ram[90][9] ), 
	.A(\ram[88][9] ));
   MUX4EHD U6938 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5483), 
	.D(\ram[87][9] ), 
	.C(\ram[85][9] ), 
	.B(\ram[86][9] ), 
	.A(\ram[84][9] ));
   MUX4EHD U6939 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5484), 
	.D(\ram[83][9] ), 
	.C(\ram[81][9] ), 
	.B(\ram[82][9] ), 
	.A(\ram[80][9] ));
   MUX4EHD U6940 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5485), 
	.D(n5481), 
	.C(n5483), 
	.B(n5482), 
	.A(n5484));
   MUX4EHD U6941 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5486), 
	.D(\ram[79][9] ), 
	.C(\ram[77][9] ), 
	.B(\ram[78][9] ), 
	.A(\ram[76][9] ));
   MUX4EHD U6942 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5487), 
	.D(\ram[75][9] ), 
	.C(\ram[73][9] ), 
	.B(\ram[74][9] ), 
	.A(\ram[72][9] ));
   MUX4EHD U6943 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5488), 
	.D(\ram[71][9] ), 
	.C(\ram[69][9] ), 
	.B(\ram[70][9] ), 
	.A(\ram[68][9] ));
   MUX4EHD U6944 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5489), 
	.D(\ram[67][9] ), 
	.C(\ram[65][9] ), 
	.B(\ram[66][9] ), 
	.A(\ram[64][9] ));
   MUX4EHD U6945 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5490), 
	.D(n5486), 
	.C(n5488), 
	.B(n5487), 
	.A(n5489));
   MUX4EHD U6946 (.S1(n6038), 
	.S0(n7444), 
	.O(n5491), 
	.D(n5475), 
	.C(n5485), 
	.B(n5480), 
	.A(n5490));
   MUX4EHD U6947 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5492), 
	.D(\ram[63][9] ), 
	.C(\ram[61][9] ), 
	.B(\ram[62][9] ), 
	.A(\ram[60][9] ));
   MUX4EHD U6948 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5493), 
	.D(\ram[59][9] ), 
	.C(\ram[57][9] ), 
	.B(\ram[58][9] ), 
	.A(\ram[56][9] ));
   MUX4EHD U6949 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5494), 
	.D(\ram[55][9] ), 
	.C(\ram[53][9] ), 
	.B(\ram[54][9] ), 
	.A(\ram[52][9] ));
   MUX4EHD U6950 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5495), 
	.D(\ram[51][9] ), 
	.C(\ram[49][9] ), 
	.B(\ram[50][9] ), 
	.A(\ram[48][9] ));
   MUX4EHD U6951 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5496), 
	.D(n5492), 
	.C(n5494), 
	.B(n5493), 
	.A(n5495));
   MUX4EHD U6952 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5497), 
	.D(\ram[47][9] ), 
	.C(\ram[45][9] ), 
	.B(\ram[46][9] ), 
	.A(\ram[44][9] ));
   MUX4EHD U6953 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5498), 
	.D(\ram[43][9] ), 
	.C(\ram[41][9] ), 
	.B(\ram[42][9] ), 
	.A(\ram[40][9] ));
   MUX4EHD U6954 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5499), 
	.D(\ram[39][9] ), 
	.C(\ram[37][9] ), 
	.B(\ram[38][9] ), 
	.A(\ram[36][9] ));
   MUX4EHD U6955 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5500), 
	.D(\ram[35][9] ), 
	.C(\ram[33][9] ), 
	.B(\ram[34][9] ), 
	.A(\ram[32][9] ));
   MUX4EHD U6956 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5501), 
	.D(n5497), 
	.C(n5499), 
	.B(n5498), 
	.A(n5500));
   MUX4EHD U6957 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5502), 
	.D(\ram[31][9] ), 
	.C(\ram[29][9] ), 
	.B(\ram[30][9] ), 
	.A(\ram[28][9] ));
   MUX4EHD U6958 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5503), 
	.D(\ram[27][9] ), 
	.C(\ram[25][9] ), 
	.B(\ram[26][9] ), 
	.A(\ram[24][9] ));
   MUX4EHD U6959 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5504), 
	.D(\ram[23][9] ), 
	.C(\ram[21][9] ), 
	.B(\ram[22][9] ), 
	.A(\ram[20][9] ));
   MUX4EHD U6960 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5505), 
	.D(\ram[19][9] ), 
	.C(\ram[17][9] ), 
	.B(\ram[18][9] ), 
	.A(\ram[16][9] ));
   MUX4EHD U6961 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5506), 
	.D(n5502), 
	.C(n5504), 
	.B(n5503), 
	.A(n5505));
   MUX4EHD U6962 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5507), 
	.D(\ram[15][9] ), 
	.C(\ram[13][9] ), 
	.B(\ram[14][9] ), 
	.A(\ram[12][9] ));
   MUX4EHD U6963 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5508), 
	.D(\ram[11][9] ), 
	.C(\ram[9][9] ), 
	.B(\ram[10][9] ), 
	.A(\ram[8][9] ));
   MUX4EHD U6964 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5509), 
	.D(\ram[7][9] ), 
	.C(\ram[5][9] ), 
	.B(\ram[6][9] ), 
	.A(\ram[4][9] ));
   MUX4EHD U6965 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5510), 
	.D(\ram[3][9] ), 
	.C(\ram[1][9] ), 
	.B(\ram[2][9] ), 
	.A(\ram[0][9] ));
   MUX4EHD U6966 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5511), 
	.D(n5507), 
	.C(n5509), 
	.B(n5508), 
	.A(n5510));
   MUX4EHD U6967 (.S1(n6038), 
	.S0(n7444), 
	.O(n5512), 
	.D(n5496), 
	.C(n5506), 
	.B(n5501), 
	.A(n5511));
   MUX4EHD U6968 (.S1(n6469), 
	.S0(n6470), 
	.O(N4132), 
	.D(n5449), 
	.C(n5491), 
	.B(n5470), 
	.A(n5512));
   MUX4EHD U6969 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5513), 
	.D(\ram[255][10] ), 
	.C(\ram[253][10] ), 
	.B(\ram[254][10] ), 
	.A(\ram[252][10] ));
   MUX4EHD U6970 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5514), 
	.D(\ram[251][10] ), 
	.C(\ram[249][10] ), 
	.B(\ram[250][10] ), 
	.A(\ram[248][10] ));
   MUX4EHD U6971 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5515), 
	.D(\ram[247][10] ), 
	.C(\ram[245][10] ), 
	.B(\ram[246][10] ), 
	.A(\ram[244][10] ));
   MUX4EHD U6972 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5516), 
	.D(\ram[243][10] ), 
	.C(\ram[241][10] ), 
	.B(\ram[242][10] ), 
	.A(\ram[240][10] ));
   MUX4EHD U6973 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5517), 
	.D(n5513), 
	.C(n5515), 
	.B(n5514), 
	.A(n5516));
   MUX4EHD U6974 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5518), 
	.D(\ram[239][10] ), 
	.C(\ram[237][10] ), 
	.B(\ram[238][10] ), 
	.A(\ram[236][10] ));
   MUX4EHD U6975 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5519), 
	.D(\ram[235][10] ), 
	.C(\ram[233][10] ), 
	.B(\ram[234][10] ), 
	.A(\ram[232][10] ));
   MUX4EHD U6976 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5520), 
	.D(\ram[231][10] ), 
	.C(\ram[229][10] ), 
	.B(\ram[230][10] ), 
	.A(\ram[228][10] ));
   MUX4EHD U6977 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5521), 
	.D(\ram[227][10] ), 
	.C(\ram[225][10] ), 
	.B(\ram[226][10] ), 
	.A(\ram[224][10] ));
   MUX4EHD U6978 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5522), 
	.D(n5518), 
	.C(n5520), 
	.B(n5519), 
	.A(n5521));
   MUX4EHD U6979 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5523), 
	.D(\ram[223][10] ), 
	.C(\ram[221][10] ), 
	.B(\ram[222][10] ), 
	.A(\ram[220][10] ));
   MUX4EHD U6980 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5524), 
	.D(\ram[219][10] ), 
	.C(\ram[217][10] ), 
	.B(\ram[218][10] ), 
	.A(\ram[216][10] ));
   MUX4EHD U6981 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5525), 
	.D(\ram[215][10] ), 
	.C(\ram[213][10] ), 
	.B(\ram[214][10] ), 
	.A(\ram[212][10] ));
   MUX4EHD U6982 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5526), 
	.D(\ram[211][10] ), 
	.C(\ram[209][10] ), 
	.B(\ram[210][10] ), 
	.A(\ram[208][10] ));
   MUX4EHD U6983 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5527), 
	.D(n5523), 
	.C(n5525), 
	.B(n5524), 
	.A(n5526));
   MUX4EHD U6984 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5528), 
	.D(\ram[207][10] ), 
	.C(\ram[205][10] ), 
	.B(\ram[206][10] ), 
	.A(\ram[204][10] ));
   MUX4EHD U6985 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5529), 
	.D(\ram[203][10] ), 
	.C(\ram[201][10] ), 
	.B(\ram[202][10] ), 
	.A(\ram[200][10] ));
   MUX4EHD U6986 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5530), 
	.D(\ram[199][10] ), 
	.C(\ram[197][10] ), 
	.B(\ram[198][10] ), 
	.A(\ram[196][10] ));
   MUX4EHD U6987 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5531), 
	.D(\ram[195][10] ), 
	.C(\ram[193][10] ), 
	.B(\ram[194][10] ), 
	.A(\ram[192][10] ));
   MUX4EHD U6988 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5532), 
	.D(n5528), 
	.C(n5530), 
	.B(n5529), 
	.A(n5531));
   MUX4EHD U6989 (.S1(n6038), 
	.S0(n7444), 
	.O(n5533), 
	.D(n5517), 
	.C(n5527), 
	.B(n5522), 
	.A(n5532));
   MUX4EHD U6990 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5534), 
	.D(\ram[191][10] ), 
	.C(\ram[189][10] ), 
	.B(\ram[190][10] ), 
	.A(\ram[188][10] ));
   MUX4EHD U6991 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5535), 
	.D(\ram[187][10] ), 
	.C(\ram[185][10] ), 
	.B(\ram[186][10] ), 
	.A(\ram[184][10] ));
   MUX4EHD U6992 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5536), 
	.D(\ram[183][10] ), 
	.C(\ram[181][10] ), 
	.B(\ram[182][10] ), 
	.A(\ram[180][10] ));
   MUX4EHD U6993 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5537), 
	.D(\ram[179][10] ), 
	.C(\ram[177][10] ), 
	.B(\ram[178][10] ), 
	.A(\ram[176][10] ));
   MUX4EHD U6994 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5538), 
	.D(n5534), 
	.C(n5536), 
	.B(n5535), 
	.A(n5537));
   MUX4EHD U6995 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5539), 
	.D(\ram[175][10] ), 
	.C(\ram[173][10] ), 
	.B(\ram[174][10] ), 
	.A(\ram[172][10] ));
   MUX4EHD U6996 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5540), 
	.D(\ram[171][10] ), 
	.C(\ram[169][10] ), 
	.B(\ram[170][10] ), 
	.A(\ram[168][10] ));
   MUX4EHD U6997 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5541), 
	.D(\ram[167][10] ), 
	.C(\ram[165][10] ), 
	.B(\ram[166][10] ), 
	.A(\ram[164][10] ));
   MUX4EHD U6998 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5542), 
	.D(\ram[163][10] ), 
	.C(\ram[161][10] ), 
	.B(\ram[162][10] ), 
	.A(\ram[160][10] ));
   MUX4EHD U6999 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5543), 
	.D(n5539), 
	.C(n5541), 
	.B(n5540), 
	.A(n5542));
   MUX4EHD U7000 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5544), 
	.D(\ram[159][10] ), 
	.C(\ram[157][10] ), 
	.B(\ram[158][10] ), 
	.A(\ram[156][10] ));
   MUX4EHD U7001 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5545), 
	.D(\ram[155][10] ), 
	.C(\ram[153][10] ), 
	.B(\ram[154][10] ), 
	.A(\ram[152][10] ));
   MUX4EHD U7002 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5546), 
	.D(\ram[151][10] ), 
	.C(\ram[149][10] ), 
	.B(\ram[150][10] ), 
	.A(\ram[148][10] ));
   MUX4EHD U7003 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5547), 
	.D(\ram[147][10] ), 
	.C(\ram[145][10] ), 
	.B(\ram[146][10] ), 
	.A(\ram[144][10] ));
   MUX4EHD U7004 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5548), 
	.D(n5544), 
	.C(n5546), 
	.B(n5545), 
	.A(n5547));
   MUX4EHD U7005 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5549), 
	.D(\ram[143][10] ), 
	.C(\ram[141][10] ), 
	.B(\ram[142][10] ), 
	.A(\ram[140][10] ));
   MUX4EHD U7006 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5550), 
	.D(\ram[139][10] ), 
	.C(\ram[137][10] ), 
	.B(\ram[138][10] ), 
	.A(\ram[136][10] ));
   MUX4EHD U7007 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5551), 
	.D(\ram[135][10] ), 
	.C(\ram[133][10] ), 
	.B(\ram[134][10] ), 
	.A(\ram[132][10] ));
   MUX4EHD U7008 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5552), 
	.D(\ram[131][10] ), 
	.C(\ram[129][10] ), 
	.B(\ram[130][10] ), 
	.A(\ram[128][10] ));
   MUX4EHD U7009 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5553), 
	.D(n5549), 
	.C(n5551), 
	.B(n5550), 
	.A(n5552));
   MUX4EHD U7010 (.S1(n6038), 
	.S0(n7444), 
	.O(n5554), 
	.D(n5538), 
	.C(n5548), 
	.B(n5543), 
	.A(n5553));
   MUX4EHD U7011 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5555), 
	.D(\ram[127][10] ), 
	.C(\ram[125][10] ), 
	.B(\ram[126][10] ), 
	.A(\ram[124][10] ));
   MUX4EHD U7012 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5556), 
	.D(\ram[123][10] ), 
	.C(\ram[121][10] ), 
	.B(\ram[122][10] ), 
	.A(\ram[120][10] ));
   MUX4EHD U7013 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5557), 
	.D(\ram[119][10] ), 
	.C(\ram[117][10] ), 
	.B(\ram[118][10] ), 
	.A(\ram[116][10] ));
   MUX4EHD U7014 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5558), 
	.D(\ram[115][10] ), 
	.C(\ram[113][10] ), 
	.B(\ram[114][10] ), 
	.A(\ram[112][10] ));
   MUX4EHD U7015 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5559), 
	.D(n5555), 
	.C(n5557), 
	.B(n5556), 
	.A(n5558));
   MUX4EHD U7016 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5560), 
	.D(\ram[111][10] ), 
	.C(\ram[109][10] ), 
	.B(\ram[110][10] ), 
	.A(\ram[108][10] ));
   MUX4EHD U7017 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5561), 
	.D(\ram[107][10] ), 
	.C(\ram[105][10] ), 
	.B(\ram[106][10] ), 
	.A(\ram[104][10] ));
   MUX4EHD U7018 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5562), 
	.D(\ram[103][10] ), 
	.C(\ram[101][10] ), 
	.B(\ram[102][10] ), 
	.A(\ram[100][10] ));
   MUX4EHD U7019 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5563), 
	.D(\ram[99][10] ), 
	.C(\ram[97][10] ), 
	.B(\ram[98][10] ), 
	.A(\ram[96][10] ));
   MUX4EHD U7020 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5564), 
	.D(n5560), 
	.C(n5562), 
	.B(n5561), 
	.A(n5563));
   MUX4EHD U7021 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5565), 
	.D(\ram[95][10] ), 
	.C(\ram[93][10] ), 
	.B(\ram[94][10] ), 
	.A(\ram[92][10] ));
   MUX4EHD U7022 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5566), 
	.D(\ram[91][10] ), 
	.C(\ram[89][10] ), 
	.B(\ram[90][10] ), 
	.A(\ram[88][10] ));
   MUX4EHD U7023 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5567), 
	.D(\ram[87][10] ), 
	.C(\ram[85][10] ), 
	.B(\ram[86][10] ), 
	.A(\ram[84][10] ));
   MUX4EHD U7024 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5568), 
	.D(\ram[83][10] ), 
	.C(\ram[81][10] ), 
	.B(\ram[82][10] ), 
	.A(\ram[80][10] ));
   MUX4EHD U7025 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5569), 
	.D(n5565), 
	.C(n5567), 
	.B(n5566), 
	.A(n5568));
   MUX4EHD U7026 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5570), 
	.D(\ram[79][10] ), 
	.C(\ram[77][10] ), 
	.B(\ram[78][10] ), 
	.A(\ram[76][10] ));
   MUX4EHD U7027 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5571), 
	.D(\ram[75][10] ), 
	.C(\ram[73][10] ), 
	.B(\ram[74][10] ), 
	.A(\ram[72][10] ));
   MUX4EHD U7028 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5572), 
	.D(\ram[71][10] ), 
	.C(\ram[69][10] ), 
	.B(\ram[70][10] ), 
	.A(\ram[68][10] ));
   MUX4EHD U7029 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5573), 
	.D(\ram[67][10] ), 
	.C(\ram[65][10] ), 
	.B(\ram[66][10] ), 
	.A(\ram[64][10] ));
   MUX4EHD U7030 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5574), 
	.D(n5570), 
	.C(n5572), 
	.B(n5571), 
	.A(n5573));
   MUX4EHD U7031 (.S1(n6038), 
	.S0(n7444), 
	.O(n5575), 
	.D(n5559), 
	.C(n5569), 
	.B(n5564), 
	.A(n5574));
   MUX4EHD U7032 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5576), 
	.D(\ram[63][10] ), 
	.C(\ram[61][10] ), 
	.B(\ram[62][10] ), 
	.A(\ram[60][10] ));
   MUX4EHD U7033 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5577), 
	.D(\ram[59][10] ), 
	.C(\ram[57][10] ), 
	.B(\ram[58][10] ), 
	.A(\ram[56][10] ));
   MUX4EHD U7034 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5578), 
	.D(\ram[55][10] ), 
	.C(\ram[53][10] ), 
	.B(\ram[54][10] ), 
	.A(\ram[52][10] ));
   MUX4EHD U7035 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5579), 
	.D(\ram[51][10] ), 
	.C(\ram[49][10] ), 
	.B(\ram[50][10] ), 
	.A(\ram[48][10] ));
   MUX4EHD U7036 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5580), 
	.D(n5576), 
	.C(n5578), 
	.B(n5577), 
	.A(n5579));
   MUX4EHD U7037 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5581), 
	.D(\ram[47][10] ), 
	.C(\ram[45][10] ), 
	.B(\ram[46][10] ), 
	.A(\ram[44][10] ));
   MUX4EHD U7038 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5582), 
	.D(\ram[43][10] ), 
	.C(\ram[41][10] ), 
	.B(\ram[42][10] ), 
	.A(\ram[40][10] ));
   MUX4EHD U7039 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5583), 
	.D(\ram[39][10] ), 
	.C(\ram[37][10] ), 
	.B(\ram[38][10] ), 
	.A(\ram[36][10] ));
   MUX4EHD U7040 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5584), 
	.D(\ram[35][10] ), 
	.C(\ram[33][10] ), 
	.B(\ram[34][10] ), 
	.A(\ram[32][10] ));
   MUX4EHD U7041 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5585), 
	.D(n5581), 
	.C(n5583), 
	.B(n5582), 
	.A(n5584));
   MUX4EHD U7042 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5586), 
	.D(\ram[31][10] ), 
	.C(\ram[29][10] ), 
	.B(\ram[30][10] ), 
	.A(\ram[28][10] ));
   MUX4EHD U7043 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5587), 
	.D(\ram[27][10] ), 
	.C(\ram[25][10] ), 
	.B(\ram[26][10] ), 
	.A(\ram[24][10] ));
   MUX4EHD U7044 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5588), 
	.D(\ram[23][10] ), 
	.C(\ram[21][10] ), 
	.B(\ram[22][10] ), 
	.A(\ram[20][10] ));
   MUX4EHD U7045 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5589), 
	.D(\ram[19][10] ), 
	.C(\ram[17][10] ), 
	.B(\ram[18][10] ), 
	.A(\ram[16][10] ));
   MUX4EHD U7046 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5590), 
	.D(n5586), 
	.C(n5588), 
	.B(n5587), 
	.A(n5589));
   MUX4EHD U7047 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5591), 
	.D(\ram[15][10] ), 
	.C(\ram[13][10] ), 
	.B(\ram[14][10] ), 
	.A(\ram[12][10] ));
   MUX4EHD U7048 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5592), 
	.D(\ram[11][10] ), 
	.C(\ram[9][10] ), 
	.B(\ram[10][10] ), 
	.A(\ram[8][10] ));
   MUX4EHD U7049 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5593), 
	.D(\ram[7][10] ), 
	.C(\ram[5][10] ), 
	.B(\ram[6][10] ), 
	.A(\ram[4][10] ));
   MUX4EHD U7050 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5594), 
	.D(\ram[3][10] ), 
	.C(\ram[1][10] ), 
	.B(\ram[2][10] ), 
	.A(\ram[0][10] ));
   MUX4EHD U7051 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5595), 
	.D(n5591), 
	.C(n5593), 
	.B(n5592), 
	.A(n5594));
   MUX4EHD U7052 (.S1(n6038), 
	.S0(n7444), 
	.O(n5596), 
	.D(n5580), 
	.C(n5590), 
	.B(n5585), 
	.A(n5595));
   MUX4EHD U7053 (.S1(n6469), 
	.S0(n6470), 
	.O(N4131), 
	.D(n5533), 
	.C(n5575), 
	.B(n5554), 
	.A(n5596));
   MUX4EHD U7054 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5597), 
	.D(\ram[255][11] ), 
	.C(\ram[253][11] ), 
	.B(\ram[254][11] ), 
	.A(\ram[252][11] ));
   MUX4EHD U7055 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5598), 
	.D(\ram[251][11] ), 
	.C(\ram[249][11] ), 
	.B(\ram[250][11] ), 
	.A(\ram[248][11] ));
   MUX4EHD U7056 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5599), 
	.D(\ram[247][11] ), 
	.C(\ram[245][11] ), 
	.B(\ram[246][11] ), 
	.A(\ram[244][11] ));
   MUX4EHD U7057 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5600), 
	.D(\ram[243][11] ), 
	.C(\ram[241][11] ), 
	.B(\ram[242][11] ), 
	.A(\ram[240][11] ));
   MUX4EHD U7058 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5601), 
	.D(n5597), 
	.C(n5599), 
	.B(n5598), 
	.A(n5600));
   MUX4EHD U7059 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5602), 
	.D(\ram[239][11] ), 
	.C(\ram[237][11] ), 
	.B(\ram[238][11] ), 
	.A(\ram[236][11] ));
   MUX4EHD U7060 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5603), 
	.D(\ram[235][11] ), 
	.C(\ram[233][11] ), 
	.B(\ram[234][11] ), 
	.A(\ram[232][11] ));
   MUX4EHD U7061 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5604), 
	.D(\ram[231][11] ), 
	.C(\ram[229][11] ), 
	.B(\ram[230][11] ), 
	.A(\ram[228][11] ));
   MUX4EHD U7062 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5605), 
	.D(\ram[227][11] ), 
	.C(\ram[225][11] ), 
	.B(\ram[226][11] ), 
	.A(\ram[224][11] ));
   MUX4EHD U7063 (.S1(n6136), 
	.S0(n7442), 
	.O(n5606), 
	.D(n5602), 
	.C(n5604), 
	.B(n5603), 
	.A(n5605));
   MUX4EHD U7064 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5607), 
	.D(\ram[223][11] ), 
	.C(\ram[221][11] ), 
	.B(\ram[222][11] ), 
	.A(\ram[220][11] ));
   MUX4EHD U7065 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5608), 
	.D(\ram[219][11] ), 
	.C(\ram[217][11] ), 
	.B(\ram[218][11] ), 
	.A(\ram[216][11] ));
   MUX4EHD U7066 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5609), 
	.D(\ram[215][11] ), 
	.C(\ram[213][11] ), 
	.B(\ram[214][11] ), 
	.A(\ram[212][11] ));
   MUX4EHD U7067 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5610), 
	.D(\ram[211][11] ), 
	.C(\ram[209][11] ), 
	.B(\ram[210][11] ), 
	.A(\ram[208][11] ));
   MUX4EHD U7068 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5611), 
	.D(n5607), 
	.C(n5609), 
	.B(n5608), 
	.A(n5610));
   MUX4EHD U7069 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5612), 
	.D(\ram[207][11] ), 
	.C(\ram[205][11] ), 
	.B(\ram[206][11] ), 
	.A(\ram[204][11] ));
   MUX4EHD U7070 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5613), 
	.D(\ram[203][11] ), 
	.C(\ram[201][11] ), 
	.B(\ram[202][11] ), 
	.A(\ram[200][11] ));
   MUX4EHD U7071 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5614), 
	.D(\ram[199][11] ), 
	.C(\ram[197][11] ), 
	.B(\ram[198][11] ), 
	.A(\ram[196][11] ));
   MUX4EHD U7072 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5615), 
	.D(\ram[195][11] ), 
	.C(\ram[193][11] ), 
	.B(\ram[194][11] ), 
	.A(\ram[192][11] ));
   MUX4EHD U7073 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5616), 
	.D(n5612), 
	.C(n5614), 
	.B(n5613), 
	.A(n5615));
   MUX4EHD U7074 (.S1(n6038), 
	.S0(n7444), 
	.O(n5617), 
	.D(n5601), 
	.C(n5611), 
	.B(n5606), 
	.A(n5616));
   MUX4EHD U7075 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5618), 
	.D(\ram[191][11] ), 
	.C(\ram[189][11] ), 
	.B(\ram[190][11] ), 
	.A(\ram[188][11] ));
   MUX4EHD U7076 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5619), 
	.D(\ram[187][11] ), 
	.C(\ram[185][11] ), 
	.B(\ram[186][11] ), 
	.A(\ram[184][11] ));
   MUX4EHD U7077 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5620), 
	.D(\ram[183][11] ), 
	.C(\ram[181][11] ), 
	.B(\ram[182][11] ), 
	.A(\ram[180][11] ));
   MUX4EHD U7078 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5621), 
	.D(\ram[179][11] ), 
	.C(\ram[177][11] ), 
	.B(\ram[178][11] ), 
	.A(\ram[176][11] ));
   MUX4EHD U7079 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5622), 
	.D(n5618), 
	.C(n5620), 
	.B(n5619), 
	.A(n5621));
   MUX4EHD U7080 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5623), 
	.D(\ram[175][11] ), 
	.C(\ram[173][11] ), 
	.B(\ram[174][11] ), 
	.A(\ram[172][11] ));
   MUX4EHD U7081 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5624), 
	.D(\ram[171][11] ), 
	.C(\ram[169][11] ), 
	.B(\ram[170][11] ), 
	.A(\ram[168][11] ));
   MUX4EHD U7082 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5625), 
	.D(\ram[167][11] ), 
	.C(\ram[165][11] ), 
	.B(\ram[166][11] ), 
	.A(\ram[164][11] ));
   MUX4EHD U7083 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5626), 
	.D(\ram[163][11] ), 
	.C(\ram[161][11] ), 
	.B(\ram[162][11] ), 
	.A(\ram[160][11] ));
   MUX4EHD U7084 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5627), 
	.D(n5623), 
	.C(n5625), 
	.B(n5624), 
	.A(n5626));
   MUX4EHD U7085 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5628), 
	.D(\ram[159][11] ), 
	.C(\ram[157][11] ), 
	.B(\ram[158][11] ), 
	.A(\ram[156][11] ));
   MUX4EHD U7086 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5629), 
	.D(\ram[155][11] ), 
	.C(\ram[153][11] ), 
	.B(\ram[154][11] ), 
	.A(\ram[152][11] ));
   MUX4EHD U7087 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5630), 
	.D(\ram[151][11] ), 
	.C(\ram[149][11] ), 
	.B(\ram[150][11] ), 
	.A(\ram[148][11] ));
   MUX4EHD U7088 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5631), 
	.D(\ram[147][11] ), 
	.C(\ram[145][11] ), 
	.B(\ram[146][11] ), 
	.A(\ram[144][11] ));
   MUX4EHD U7089 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5632), 
	.D(n5628), 
	.C(n5630), 
	.B(n5629), 
	.A(n5631));
   MUX4EHD U7090 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5633), 
	.D(\ram[143][11] ), 
	.C(\ram[141][11] ), 
	.B(\ram[142][11] ), 
	.A(\ram[140][11] ));
   MUX4EHD U7091 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5634), 
	.D(\ram[139][11] ), 
	.C(\ram[137][11] ), 
	.B(\ram[138][11] ), 
	.A(\ram[136][11] ));
   MUX4EHD U7092 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5635), 
	.D(\ram[135][11] ), 
	.C(\ram[133][11] ), 
	.B(\ram[134][11] ), 
	.A(\ram[132][11] ));
   MUX4EHD U7093 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5636), 
	.D(\ram[131][11] ), 
	.C(\ram[129][11] ), 
	.B(\ram[130][11] ), 
	.A(\ram[128][11] ));
   MUX4EHD U7094 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5637), 
	.D(n5633), 
	.C(n5635), 
	.B(n5634), 
	.A(n5636));
   MUX4EHD U7095 (.S1(n6038), 
	.S0(n7444), 
	.O(n5638), 
	.D(n5622), 
	.C(n5632), 
	.B(n5627), 
	.A(n5637));
   MUX4EHD U7096 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5639), 
	.D(\ram[127][11] ), 
	.C(\ram[125][11] ), 
	.B(\ram[126][11] ), 
	.A(\ram[124][11] ));
   MUX4EHD U7097 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5640), 
	.D(\ram[123][11] ), 
	.C(\ram[121][11] ), 
	.B(\ram[122][11] ), 
	.A(\ram[120][11] ));
   MUX4EHD U7098 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5641), 
	.D(\ram[119][11] ), 
	.C(\ram[117][11] ), 
	.B(\ram[118][11] ), 
	.A(\ram[116][11] ));
   MUX4EHD U7099 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5642), 
	.D(\ram[115][11] ), 
	.C(\ram[113][11] ), 
	.B(\ram[114][11] ), 
	.A(\ram[112][11] ));
   MUX4EHD U7100 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5643), 
	.D(n5639), 
	.C(n5641), 
	.B(n5640), 
	.A(n5642));
   MUX4EHD U7101 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5644), 
	.D(\ram[111][11] ), 
	.C(\ram[109][11] ), 
	.B(\ram[110][11] ), 
	.A(\ram[108][11] ));
   MUX4EHD U7102 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5645), 
	.D(\ram[107][11] ), 
	.C(\ram[105][11] ), 
	.B(\ram[106][11] ), 
	.A(\ram[104][11] ));
   MUX4EHD U7103 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5646), 
	.D(\ram[103][11] ), 
	.C(\ram[101][11] ), 
	.B(\ram[102][11] ), 
	.A(\ram[100][11] ));
   MUX4EHD U7104 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5647), 
	.D(\ram[99][11] ), 
	.C(\ram[97][11] ), 
	.B(\ram[98][11] ), 
	.A(\ram[96][11] ));
   MUX4EHD U7105 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5648), 
	.D(n5644), 
	.C(n5646), 
	.B(n5645), 
	.A(n5647));
   MUX4EHD U7106 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5649), 
	.D(\ram[95][11] ), 
	.C(\ram[93][11] ), 
	.B(\ram[94][11] ), 
	.A(\ram[92][11] ));
   MUX4EHD U7107 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5650), 
	.D(\ram[91][11] ), 
	.C(\ram[89][11] ), 
	.B(\ram[90][11] ), 
	.A(\ram[88][11] ));
   MUX4EHD U7108 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5651), 
	.D(\ram[87][11] ), 
	.C(\ram[85][11] ), 
	.B(\ram[86][11] ), 
	.A(\ram[84][11] ));
   MUX4EHD U7109 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5652), 
	.D(\ram[83][11] ), 
	.C(\ram[81][11] ), 
	.B(\ram[82][11] ), 
	.A(\ram[80][11] ));
   MUX4EHD U7110 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5653), 
	.D(n5649), 
	.C(n5651), 
	.B(n5650), 
	.A(n5652));
   MUX4EHD U7111 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5654), 
	.D(\ram[79][11] ), 
	.C(\ram[77][11] ), 
	.B(\ram[78][11] ), 
	.A(\ram[76][11] ));
   MUX4EHD U7112 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5655), 
	.D(\ram[75][11] ), 
	.C(\ram[73][11] ), 
	.B(\ram[74][11] ), 
	.A(\ram[72][11] ));
   MUX4EHD U7113 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5656), 
	.D(\ram[71][11] ), 
	.C(\ram[69][11] ), 
	.B(\ram[70][11] ), 
	.A(\ram[68][11] ));
   MUX4EHD U7114 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5657), 
	.D(\ram[67][11] ), 
	.C(\ram[65][11] ), 
	.B(\ram[66][11] ), 
	.A(\ram[64][11] ));
   MUX4EHD U7115 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5658), 
	.D(n5654), 
	.C(n5656), 
	.B(n5655), 
	.A(n5657));
   MUX4EHD U7116 (.S1(n6038), 
	.S0(n7444), 
	.O(n5659), 
	.D(n5643), 
	.C(n5653), 
	.B(n5648), 
	.A(n5658));
   MUX4EHD U7117 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5660), 
	.D(\ram[63][11] ), 
	.C(\ram[61][11] ), 
	.B(\ram[62][11] ), 
	.A(\ram[60][11] ));
   MUX4EHD U7118 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5661), 
	.D(\ram[59][11] ), 
	.C(\ram[57][11] ), 
	.B(\ram[58][11] ), 
	.A(\ram[56][11] ));
   MUX4EHD U7119 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5662), 
	.D(\ram[55][11] ), 
	.C(\ram[53][11] ), 
	.B(\ram[54][11] ), 
	.A(\ram[52][11] ));
   MUX4EHD U7120 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5663), 
	.D(\ram[51][11] ), 
	.C(\ram[49][11] ), 
	.B(\ram[50][11] ), 
	.A(\ram[48][11] ));
   MUX4EHD U7121 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5664), 
	.D(n5660), 
	.C(n5662), 
	.B(n5661), 
	.A(n5663));
   MUX4EHD U7122 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5665), 
	.D(\ram[47][11] ), 
	.C(\ram[45][11] ), 
	.B(\ram[46][11] ), 
	.A(\ram[44][11] ));
   MUX4EHD U7123 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5666), 
	.D(\ram[43][11] ), 
	.C(\ram[41][11] ), 
	.B(\ram[42][11] ), 
	.A(\ram[40][11] ));
   MUX4EHD U7124 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5667), 
	.D(\ram[39][11] ), 
	.C(\ram[37][11] ), 
	.B(\ram[38][11] ), 
	.A(\ram[36][11] ));
   MUX4EHD U7125 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5668), 
	.D(\ram[35][11] ), 
	.C(\ram[33][11] ), 
	.B(\ram[34][11] ), 
	.A(\ram[32][11] ));
   MUX4EHD U7126 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5669), 
	.D(n5665), 
	.C(n5667), 
	.B(n5666), 
	.A(n5668));
   MUX4EHD U7127 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5670), 
	.D(\ram[31][11] ), 
	.C(\ram[29][11] ), 
	.B(\ram[30][11] ), 
	.A(\ram[28][11] ));
   MUX4EHD U7128 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5671), 
	.D(\ram[27][11] ), 
	.C(\ram[25][11] ), 
	.B(\ram[26][11] ), 
	.A(\ram[24][11] ));
   MUX4EHD U7129 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5672), 
	.D(\ram[23][11] ), 
	.C(\ram[21][11] ), 
	.B(\ram[22][11] ), 
	.A(\ram[20][11] ));
   MUX4EHD U7130 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5673), 
	.D(\ram[19][11] ), 
	.C(\ram[17][11] ), 
	.B(\ram[18][11] ), 
	.A(\ram[16][11] ));
   MUX4EHD U7131 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5674), 
	.D(n5670), 
	.C(n5672), 
	.B(n5671), 
	.A(n5673));
   MUX4EHD U7132 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5675), 
	.D(\ram[15][11] ), 
	.C(\ram[13][11] ), 
	.B(\ram[14][11] ), 
	.A(\ram[12][11] ));
   MUX4EHD U7133 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5676), 
	.D(\ram[11][11] ), 
	.C(\ram[9][11] ), 
	.B(\ram[10][11] ), 
	.A(\ram[8][11] ));
   MUX4EHD U7134 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5677), 
	.D(\ram[7][11] ), 
	.C(\ram[5][11] ), 
	.B(\ram[6][11] ), 
	.A(\ram[4][11] ));
   MUX4EHD U7135 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5678), 
	.D(\ram[3][11] ), 
	.C(\ram[1][11] ), 
	.B(\ram[2][11] ), 
	.A(\ram[0][11] ));
   MUX4EHD U7136 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5679), 
	.D(n5675), 
	.C(n5677), 
	.B(n5676), 
	.A(n5678));
   MUX4EHD U7137 (.S1(n6038), 
	.S0(n7444), 
	.O(n5680), 
	.D(n5664), 
	.C(n5674), 
	.B(n5669), 
	.A(n5679));
   MUX4EHD U7138 (.S1(n6469), 
	.S0(n6470), 
	.O(N4130), 
	.D(n5617), 
	.C(n5659), 
	.B(n5638), 
	.A(n5680));
   MUX4EHD U7139 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5681), 
	.D(\ram[255][12] ), 
	.C(\ram[253][12] ), 
	.B(\ram[254][12] ), 
	.A(\ram[252][12] ));
   MUX4EHD U7140 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5682), 
	.D(\ram[251][12] ), 
	.C(\ram[249][12] ), 
	.B(\ram[250][12] ), 
	.A(\ram[248][12] ));
   MUX4EHD U7141 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5683), 
	.D(\ram[247][12] ), 
	.C(\ram[245][12] ), 
	.B(\ram[246][12] ), 
	.A(\ram[244][12] ));
   MUX4EHD U7142 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5684), 
	.D(\ram[243][12] ), 
	.C(\ram[241][12] ), 
	.B(\ram[242][12] ), 
	.A(\ram[240][12] ));
   MUX4EHD U7143 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5685), 
	.D(n5681), 
	.C(n5683), 
	.B(n5682), 
	.A(n5684));
   MUX4EHD U7144 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5686), 
	.D(\ram[239][12] ), 
	.C(\ram[237][12] ), 
	.B(\ram[238][12] ), 
	.A(\ram[236][12] ));
   MUX4EHD U7145 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5687), 
	.D(\ram[235][12] ), 
	.C(\ram[233][12] ), 
	.B(\ram[234][12] ), 
	.A(\ram[232][12] ));
   MUX4EHD U7146 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5688), 
	.D(\ram[231][12] ), 
	.C(\ram[229][12] ), 
	.B(\ram[230][12] ), 
	.A(\ram[228][12] ));
   MUX4EHD U7147 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5689), 
	.D(\ram[227][12] ), 
	.C(\ram[225][12] ), 
	.B(\ram[226][12] ), 
	.A(\ram[224][12] ));
   MUX4EHD U7148 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5690), 
	.D(n5686), 
	.C(n5688), 
	.B(n5687), 
	.A(n5689));
   MUX4EHD U7149 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5691), 
	.D(\ram[223][12] ), 
	.C(\ram[221][12] ), 
	.B(\ram[222][12] ), 
	.A(\ram[220][12] ));
   MUX4EHD U7150 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5692), 
	.D(\ram[219][12] ), 
	.C(\ram[217][12] ), 
	.B(\ram[218][12] ), 
	.A(\ram[216][12] ));
   MUX4EHD U7151 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5693), 
	.D(\ram[215][12] ), 
	.C(\ram[213][12] ), 
	.B(\ram[214][12] ), 
	.A(\ram[212][12] ));
   MUX4EHD U7152 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5694), 
	.D(\ram[211][12] ), 
	.C(\ram[209][12] ), 
	.B(\ram[210][12] ), 
	.A(\ram[208][12] ));
   MUX4EHD U7153 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5695), 
	.D(n5691), 
	.C(n5693), 
	.B(n5692), 
	.A(n5694));
   MUX4EHD U7154 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5696), 
	.D(\ram[207][12] ), 
	.C(\ram[205][12] ), 
	.B(\ram[206][12] ), 
	.A(\ram[204][12] ));
   MUX4EHD U7155 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5697), 
	.D(\ram[203][12] ), 
	.C(\ram[201][12] ), 
	.B(\ram[202][12] ), 
	.A(\ram[200][12] ));
   MUX4EHD U7156 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5698), 
	.D(\ram[199][12] ), 
	.C(\ram[197][12] ), 
	.B(\ram[198][12] ), 
	.A(\ram[196][12] ));
   MUX4EHD U7157 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5699), 
	.D(\ram[195][12] ), 
	.C(\ram[193][12] ), 
	.B(\ram[194][12] ), 
	.A(\ram[192][12] ));
   MUX4EHD U7158 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5700), 
	.D(n5696), 
	.C(n5698), 
	.B(n5697), 
	.A(n5699));
   MUX4EHD U7159 (.S1(n6038), 
	.S0(n7444), 
	.O(n5701), 
	.D(n5685), 
	.C(n5695), 
	.B(n5690), 
	.A(n5700));
   MUX4EHD U7160 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5702), 
	.D(\ram[191][12] ), 
	.C(\ram[189][12] ), 
	.B(\ram[190][12] ), 
	.A(\ram[188][12] ));
   MUX4EHD U7161 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5703), 
	.D(\ram[187][12] ), 
	.C(\ram[185][12] ), 
	.B(\ram[186][12] ), 
	.A(\ram[184][12] ));
   MUX4EHD U7162 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5704), 
	.D(\ram[183][12] ), 
	.C(\ram[181][12] ), 
	.B(\ram[182][12] ), 
	.A(\ram[180][12] ));
   MUX4EHD U7163 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5705), 
	.D(\ram[179][12] ), 
	.C(\ram[177][12] ), 
	.B(\ram[178][12] ), 
	.A(\ram[176][12] ));
   MUX4EHD U7164 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5706), 
	.D(n5702), 
	.C(n5704), 
	.B(n5703), 
	.A(n5705));
   MUX4EHD U7165 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5707), 
	.D(\ram[175][12] ), 
	.C(\ram[173][12] ), 
	.B(\ram[174][12] ), 
	.A(\ram[172][12] ));
   MUX4EHD U7166 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5708), 
	.D(\ram[171][12] ), 
	.C(\ram[169][12] ), 
	.B(\ram[170][12] ), 
	.A(\ram[168][12] ));
   MUX4EHD U7167 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5709), 
	.D(\ram[167][12] ), 
	.C(\ram[165][12] ), 
	.B(\ram[166][12] ), 
	.A(\ram[164][12] ));
   MUX4EHD U7168 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5710), 
	.D(\ram[163][12] ), 
	.C(\ram[161][12] ), 
	.B(\ram[162][12] ), 
	.A(\ram[160][12] ));
   MUX4EHD U7169 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5711), 
	.D(n5707), 
	.C(n5709), 
	.B(n5708), 
	.A(n5710));
   MUX4EHD U7170 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5712), 
	.D(\ram[159][12] ), 
	.C(\ram[157][12] ), 
	.B(\ram[158][12] ), 
	.A(\ram[156][12] ));
   MUX4EHD U7171 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5713), 
	.D(\ram[155][12] ), 
	.C(\ram[153][12] ), 
	.B(\ram[154][12] ), 
	.A(\ram[152][12] ));
   MUX4EHD U7172 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5714), 
	.D(\ram[151][12] ), 
	.C(\ram[149][12] ), 
	.B(\ram[150][12] ), 
	.A(\ram[148][12] ));
   MUX4EHD U7173 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5715), 
	.D(\ram[147][12] ), 
	.C(\ram[145][12] ), 
	.B(\ram[146][12] ), 
	.A(\ram[144][12] ));
   MUX4EHD U7174 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5716), 
	.D(n5712), 
	.C(n5714), 
	.B(n5713), 
	.A(n5715));
   MUX4EHD U7175 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5717), 
	.D(\ram[143][12] ), 
	.C(\ram[141][12] ), 
	.B(\ram[142][12] ), 
	.A(\ram[140][12] ));
   MUX4EHD U7176 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5718), 
	.D(\ram[139][12] ), 
	.C(\ram[137][12] ), 
	.B(\ram[138][12] ), 
	.A(\ram[136][12] ));
   MUX4EHD U7177 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5719), 
	.D(\ram[135][12] ), 
	.C(\ram[133][12] ), 
	.B(\ram[134][12] ), 
	.A(\ram[132][12] ));
   MUX4EHD U7178 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5720), 
	.D(\ram[131][12] ), 
	.C(\ram[129][12] ), 
	.B(\ram[130][12] ), 
	.A(\ram[128][12] ));
   MUX4EHD U7179 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5721), 
	.D(n5717), 
	.C(n5719), 
	.B(n5718), 
	.A(n5720));
   MUX4EHD U7180 (.S1(n6038), 
	.S0(n7444), 
	.O(n5722), 
	.D(n5706), 
	.C(n5716), 
	.B(n5711), 
	.A(n5721));
   MUX4EHD U7181 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5723), 
	.D(\ram[127][12] ), 
	.C(\ram[125][12] ), 
	.B(\ram[126][12] ), 
	.A(\ram[124][12] ));
   MUX4EHD U7182 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5724), 
	.D(\ram[123][12] ), 
	.C(\ram[121][12] ), 
	.B(\ram[122][12] ), 
	.A(\ram[120][12] ));
   MUX4EHD U7183 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5725), 
	.D(\ram[119][12] ), 
	.C(\ram[117][12] ), 
	.B(\ram[118][12] ), 
	.A(\ram[116][12] ));
   MUX4EHD U7184 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5726), 
	.D(\ram[115][12] ), 
	.C(\ram[113][12] ), 
	.B(\ram[114][12] ), 
	.A(\ram[112][12] ));
   MUX4EHD U7185 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5727), 
	.D(n5723), 
	.C(n5725), 
	.B(n5724), 
	.A(n5726));
   MUX4EHD U7186 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5728), 
	.D(\ram[111][12] ), 
	.C(\ram[109][12] ), 
	.B(\ram[110][12] ), 
	.A(\ram[108][12] ));
   MUX4EHD U7187 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5729), 
	.D(\ram[107][12] ), 
	.C(\ram[105][12] ), 
	.B(\ram[106][12] ), 
	.A(\ram[104][12] ));
   MUX4EHD U7188 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5730), 
	.D(\ram[103][12] ), 
	.C(\ram[101][12] ), 
	.B(\ram[102][12] ), 
	.A(\ram[100][12] ));
   MUX4EHD U7189 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5731), 
	.D(\ram[99][12] ), 
	.C(\ram[97][12] ), 
	.B(\ram[98][12] ), 
	.A(\ram[96][12] ));
   MUX4EHD U7190 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5732), 
	.D(n5728), 
	.C(n5730), 
	.B(n5729), 
	.A(n5731));
   MUX4EHD U7191 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5733), 
	.D(\ram[95][12] ), 
	.C(\ram[93][12] ), 
	.B(\ram[94][12] ), 
	.A(\ram[92][12] ));
   MUX4EHD U7192 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5734), 
	.D(\ram[91][12] ), 
	.C(\ram[89][12] ), 
	.B(\ram[90][12] ), 
	.A(\ram[88][12] ));
   MUX4EHD U7193 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5735), 
	.D(\ram[87][12] ), 
	.C(\ram[85][12] ), 
	.B(\ram[86][12] ), 
	.A(\ram[84][12] ));
   MUX4EHD U7194 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5736), 
	.D(\ram[83][12] ), 
	.C(\ram[81][12] ), 
	.B(\ram[82][12] ), 
	.A(\ram[80][12] ));
   MUX4EHD U7195 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5737), 
	.D(n5733), 
	.C(n5735), 
	.B(n5734), 
	.A(n5736));
   MUX4EHD U7196 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5738), 
	.D(\ram[79][12] ), 
	.C(\ram[77][12] ), 
	.B(\ram[78][12] ), 
	.A(\ram[76][12] ));
   MUX4EHD U7197 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5739), 
	.D(\ram[75][12] ), 
	.C(\ram[73][12] ), 
	.B(\ram[74][12] ), 
	.A(\ram[72][12] ));
   MUX4EHD U7198 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5740), 
	.D(\ram[71][12] ), 
	.C(\ram[69][12] ), 
	.B(\ram[70][12] ), 
	.A(\ram[68][12] ));
   MUX4EHD U7199 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5741), 
	.D(\ram[67][12] ), 
	.C(\ram[65][12] ), 
	.B(\ram[66][12] ), 
	.A(\ram[64][12] ));
   MUX4EHD U7200 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5742), 
	.D(n5738), 
	.C(n5740), 
	.B(n5739), 
	.A(n5741));
   MUX4EHD U7201 (.S1(n6038), 
	.S0(n7444), 
	.O(n5743), 
	.D(n5727), 
	.C(n5737), 
	.B(n5732), 
	.A(n5742));
   MUX4EHD U7202 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5744), 
	.D(\ram[63][12] ), 
	.C(\ram[61][12] ), 
	.B(\ram[62][12] ), 
	.A(\ram[60][12] ));
   MUX4EHD U7203 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5745), 
	.D(\ram[59][12] ), 
	.C(\ram[57][12] ), 
	.B(\ram[58][12] ), 
	.A(\ram[56][12] ));
   MUX4EHD U7204 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5746), 
	.D(\ram[55][12] ), 
	.C(\ram[53][12] ), 
	.B(\ram[54][12] ), 
	.A(\ram[52][12] ));
   MUX4EHD U7205 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5747), 
	.D(\ram[51][12] ), 
	.C(\ram[49][12] ), 
	.B(\ram[50][12] ), 
	.A(\ram[48][12] ));
   MUX4EHD U7206 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5748), 
	.D(n5744), 
	.C(n5746), 
	.B(n5745), 
	.A(n5747));
   MUX4EHD U7207 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5749), 
	.D(\ram[47][12] ), 
	.C(\ram[45][12] ), 
	.B(\ram[46][12] ), 
	.A(\ram[44][12] ));
   MUX4EHD U7208 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5750), 
	.D(\ram[43][12] ), 
	.C(\ram[41][12] ), 
	.B(\ram[42][12] ), 
	.A(\ram[40][12] ));
   MUX4EHD U7209 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5751), 
	.D(\ram[39][12] ), 
	.C(\ram[37][12] ), 
	.B(\ram[38][12] ), 
	.A(\ram[36][12] ));
   MUX4EHD U7210 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5752), 
	.D(\ram[35][12] ), 
	.C(\ram[33][12] ), 
	.B(\ram[34][12] ), 
	.A(\ram[32][12] ));
   MUX4EHD U7211 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5753), 
	.D(n5749), 
	.C(n5751), 
	.B(n5750), 
	.A(n5752));
   MUX4EHD U7212 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5754), 
	.D(\ram[31][12] ), 
	.C(\ram[29][12] ), 
	.B(\ram[30][12] ), 
	.A(\ram[28][12] ));
   MUX4EHD U7213 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5755), 
	.D(\ram[27][12] ), 
	.C(\ram[25][12] ), 
	.B(\ram[26][12] ), 
	.A(\ram[24][12] ));
   MUX4EHD U7214 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5756), 
	.D(\ram[23][12] ), 
	.C(\ram[21][12] ), 
	.B(\ram[22][12] ), 
	.A(\ram[20][12] ));
   MUX4EHD U7215 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5757), 
	.D(\ram[19][12] ), 
	.C(\ram[17][12] ), 
	.B(\ram[18][12] ), 
	.A(\ram[16][12] ));
   MUX4EHD U7216 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5758), 
	.D(n5754), 
	.C(n5756), 
	.B(n5755), 
	.A(n5757));
   MUX4EHD U7217 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5759), 
	.D(\ram[15][12] ), 
	.C(\ram[13][12] ), 
	.B(\ram[14][12] ), 
	.A(\ram[12][12] ));
   MUX4EHD U7218 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5760), 
	.D(\ram[11][12] ), 
	.C(\ram[9][12] ), 
	.B(\ram[10][12] ), 
	.A(\ram[8][12] ));
   MUX4EHD U7219 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5761), 
	.D(\ram[7][12] ), 
	.C(\ram[5][12] ), 
	.B(\ram[6][12] ), 
	.A(\ram[4][12] ));
   MUX4EHD U7220 (.S1(FE_OFN30_n6459), 
	.S0(n7440), 
	.O(n5762), 
	.D(\ram[3][12] ), 
	.C(\ram[1][12] ), 
	.B(\ram[2][12] ), 
	.A(\ram[0][12] ));
   MUX4EHD U7221 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5763), 
	.D(n5759), 
	.C(n5761), 
	.B(n5760), 
	.A(n5762));
   MUX4EHD U7222 (.S1(n6038), 
	.S0(n7444), 
	.O(n5764), 
	.D(n5748), 
	.C(n5758), 
	.B(n5753), 
	.A(n5763));
   MUX4EHD U7223 (.S1(n6469), 
	.S0(n6470), 
	.O(N4129), 
	.D(n5701), 
	.C(n5743), 
	.B(n5722), 
	.A(n5764));
   MUX4EHD U7224 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5765), 
	.D(\ram[255][13] ), 
	.C(\ram[253][13] ), 
	.B(\ram[254][13] ), 
	.A(\ram[252][13] ));
   MUX4EHD U7225 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5766), 
	.D(\ram[251][13] ), 
	.C(\ram[249][13] ), 
	.B(\ram[250][13] ), 
	.A(\ram[248][13] ));
   MUX4EHD U7226 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5767), 
	.D(\ram[247][13] ), 
	.C(\ram[245][13] ), 
	.B(\ram[246][13] ), 
	.A(\ram[244][13] ));
   MUX4EHD U7227 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5768), 
	.D(\ram[243][13] ), 
	.C(\ram[241][13] ), 
	.B(\ram[242][13] ), 
	.A(\ram[240][13] ));
   MUX4EHD U7228 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5769), 
	.D(n5765), 
	.C(n5767), 
	.B(n5766), 
	.A(n5768));
   MUX4EHD U7229 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5770), 
	.D(\ram[239][13] ), 
	.C(\ram[237][13] ), 
	.B(\ram[238][13] ), 
	.A(\ram[236][13] ));
   MUX4EHD U7230 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5771), 
	.D(\ram[235][13] ), 
	.C(\ram[233][13] ), 
	.B(\ram[234][13] ), 
	.A(\ram[232][13] ));
   MUX4EHD U7231 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5772), 
	.D(\ram[231][13] ), 
	.C(\ram[229][13] ), 
	.B(\ram[230][13] ), 
	.A(\ram[228][13] ));
   MUX4EHD U7232 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5773), 
	.D(\ram[227][13] ), 
	.C(\ram[225][13] ), 
	.B(\ram[226][13] ), 
	.A(\ram[224][13] ));
   MUX4EHD U7233 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5774), 
	.D(n5770), 
	.C(n5772), 
	.B(n5771), 
	.A(n5773));
   MUX4EHD U7234 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5775), 
	.D(\ram[223][13] ), 
	.C(\ram[221][13] ), 
	.B(\ram[222][13] ), 
	.A(\ram[220][13] ));
   MUX4EHD U7235 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5776), 
	.D(\ram[219][13] ), 
	.C(\ram[217][13] ), 
	.B(\ram[218][13] ), 
	.A(\ram[216][13] ));
   MUX4EHD U7236 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5777), 
	.D(\ram[215][13] ), 
	.C(\ram[213][13] ), 
	.B(\ram[214][13] ), 
	.A(\ram[212][13] ));
   MUX4EHD U7237 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5778), 
	.D(\ram[211][13] ), 
	.C(\ram[209][13] ), 
	.B(\ram[210][13] ), 
	.A(\ram[208][13] ));
   MUX4EHD U7238 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5779), 
	.D(n5775), 
	.C(n5777), 
	.B(n5776), 
	.A(n5778));
   MUX4EHD U7239 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5780), 
	.D(\ram[207][13] ), 
	.C(\ram[205][13] ), 
	.B(\ram[206][13] ), 
	.A(\ram[204][13] ));
   MUX4EHD U7240 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5781), 
	.D(\ram[203][13] ), 
	.C(\ram[201][13] ), 
	.B(\ram[202][13] ), 
	.A(\ram[200][13] ));
   MUX4EHD U7241 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5782), 
	.D(\ram[199][13] ), 
	.C(\ram[197][13] ), 
	.B(\ram[198][13] ), 
	.A(\ram[196][13] ));
   MUX4EHD U7242 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5783), 
	.D(\ram[195][13] ), 
	.C(\ram[193][13] ), 
	.B(\ram[194][13] ), 
	.A(\ram[192][13] ));
   MUX4EHD U7243 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5784), 
	.D(n5780), 
	.C(n5782), 
	.B(n5781), 
	.A(n5783));
   MUX4EHD U7244 (.S1(n6038), 
	.S0(n7444), 
	.O(n5785), 
	.D(n5769), 
	.C(n5779), 
	.B(n5774), 
	.A(n5784));
   MUX4EHD U7245 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5786), 
	.D(\ram[191][13] ), 
	.C(\ram[189][13] ), 
	.B(\ram[190][13] ), 
	.A(\ram[188][13] ));
   MUX4EHD U7246 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5787), 
	.D(\ram[187][13] ), 
	.C(\ram[185][13] ), 
	.B(\ram[186][13] ), 
	.A(\ram[184][13] ));
   MUX4EHD U7247 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5788), 
	.D(\ram[183][13] ), 
	.C(\ram[181][13] ), 
	.B(\ram[182][13] ), 
	.A(\ram[180][13] ));
   MUX4EHD U7248 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5789), 
	.D(\ram[179][13] ), 
	.C(\ram[177][13] ), 
	.B(\ram[178][13] ), 
	.A(\ram[176][13] ));
   MUX4EHD U7249 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5790), 
	.D(n5786), 
	.C(n5788), 
	.B(n5787), 
	.A(n5789));
   MUX4EHD U7250 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5791), 
	.D(\ram[175][13] ), 
	.C(\ram[173][13] ), 
	.B(\ram[174][13] ), 
	.A(\ram[172][13] ));
   MUX4EHD U7251 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5792), 
	.D(\ram[171][13] ), 
	.C(\ram[169][13] ), 
	.B(\ram[170][13] ), 
	.A(\ram[168][13] ));
   MUX4EHD U7252 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5793), 
	.D(\ram[167][13] ), 
	.C(\ram[165][13] ), 
	.B(\ram[166][13] ), 
	.A(\ram[164][13] ));
   MUX4EHD U7253 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5794), 
	.D(\ram[163][13] ), 
	.C(\ram[161][13] ), 
	.B(\ram[162][13] ), 
	.A(\ram[160][13] ));
   MUX4EHD U7254 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5795), 
	.D(n5791), 
	.C(n5793), 
	.B(n5792), 
	.A(n5794));
   MUX4EHD U7255 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5796), 
	.D(\ram[159][13] ), 
	.C(\ram[157][13] ), 
	.B(\ram[158][13] ), 
	.A(\ram[156][13] ));
   MUX4EHD U7256 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5797), 
	.D(\ram[155][13] ), 
	.C(\ram[153][13] ), 
	.B(\ram[154][13] ), 
	.A(\ram[152][13] ));
   MUX4EHD U7257 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5798), 
	.D(\ram[151][13] ), 
	.C(\ram[149][13] ), 
	.B(\ram[150][13] ), 
	.A(\ram[148][13] ));
   MUX4EHD U7258 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5799), 
	.D(\ram[147][13] ), 
	.C(\ram[145][13] ), 
	.B(\ram[146][13] ), 
	.A(\ram[144][13] ));
   MUX4EHD U7259 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5800), 
	.D(n5796), 
	.C(n5798), 
	.B(n5797), 
	.A(n5799));
   MUX4EHD U7260 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5801), 
	.D(\ram[143][13] ), 
	.C(\ram[141][13] ), 
	.B(\ram[142][13] ), 
	.A(\ram[140][13] ));
   MUX4EHD U7261 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5802), 
	.D(\ram[139][13] ), 
	.C(\ram[137][13] ), 
	.B(\ram[138][13] ), 
	.A(\ram[136][13] ));
   MUX4EHD U7262 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5803), 
	.D(\ram[135][13] ), 
	.C(\ram[133][13] ), 
	.B(\ram[134][13] ), 
	.A(\ram[132][13] ));
   MUX4EHD U7263 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5804), 
	.D(\ram[131][13] ), 
	.C(\ram[129][13] ), 
	.B(\ram[130][13] ), 
	.A(\ram[128][13] ));
   MUX4EHD U7264 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5805), 
	.D(n5801), 
	.C(n5803), 
	.B(n5802), 
	.A(n5804));
   MUX4EHD U7265 (.S1(n6038), 
	.S0(n7444), 
	.O(n5806), 
	.D(n5790), 
	.C(n5800), 
	.B(n5795), 
	.A(n5805));
   MUX4EHD U7266 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5807), 
	.D(\ram[127][13] ), 
	.C(\ram[125][13] ), 
	.B(\ram[126][13] ), 
	.A(\ram[124][13] ));
   MUX4EHD U7267 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5808), 
	.D(\ram[123][13] ), 
	.C(\ram[121][13] ), 
	.B(\ram[122][13] ), 
	.A(\ram[120][13] ));
   MUX4EHD U7268 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5809), 
	.D(\ram[119][13] ), 
	.C(\ram[117][13] ), 
	.B(\ram[118][13] ), 
	.A(\ram[116][13] ));
   MUX4EHD U7269 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5810), 
	.D(\ram[115][13] ), 
	.C(\ram[113][13] ), 
	.B(\ram[114][13] ), 
	.A(\ram[112][13] ));
   MUX4EHD U7270 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5811), 
	.D(n5807), 
	.C(n5809), 
	.B(n5808), 
	.A(n5810));
   MUX4EHD U7271 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5812), 
	.D(\ram[111][13] ), 
	.C(\ram[109][13] ), 
	.B(\ram[110][13] ), 
	.A(\ram[108][13] ));
   MUX4EHD U7272 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5813), 
	.D(\ram[107][13] ), 
	.C(\ram[105][13] ), 
	.B(\ram[106][13] ), 
	.A(\ram[104][13] ));
   MUX4EHD U7273 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5814), 
	.D(\ram[103][13] ), 
	.C(\ram[101][13] ), 
	.B(\ram[102][13] ), 
	.A(\ram[100][13] ));
   MUX4EHD U7274 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5815), 
	.D(\ram[99][13] ), 
	.C(\ram[97][13] ), 
	.B(\ram[98][13] ), 
	.A(\ram[96][13] ));
   MUX4EHD U7275 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5816), 
	.D(n5812), 
	.C(n5814), 
	.B(n5813), 
	.A(n5815));
   MUX4EHD U7276 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5817), 
	.D(\ram[95][13] ), 
	.C(\ram[93][13] ), 
	.B(\ram[94][13] ), 
	.A(\ram[92][13] ));
   MUX4EHD U7277 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5818), 
	.D(\ram[91][13] ), 
	.C(\ram[89][13] ), 
	.B(\ram[90][13] ), 
	.A(\ram[88][13] ));
   MUX4EHD U7278 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5819), 
	.D(\ram[87][13] ), 
	.C(\ram[85][13] ), 
	.B(\ram[86][13] ), 
	.A(\ram[84][13] ));
   MUX4EHD U7279 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5820), 
	.D(\ram[83][13] ), 
	.C(\ram[81][13] ), 
	.B(\ram[82][13] ), 
	.A(\ram[80][13] ));
   MUX4EHD U7280 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5821), 
	.D(n5817), 
	.C(n5819), 
	.B(n5818), 
	.A(n5820));
   MUX4EHD U7281 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5822), 
	.D(\ram[79][13] ), 
	.C(\ram[77][13] ), 
	.B(\ram[78][13] ), 
	.A(\ram[76][13] ));
   MUX4EHD U7282 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5823), 
	.D(\ram[75][13] ), 
	.C(\ram[73][13] ), 
	.B(\ram[74][13] ), 
	.A(\ram[72][13] ));
   MUX4EHD U7283 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5824), 
	.D(\ram[71][13] ), 
	.C(\ram[69][13] ), 
	.B(\ram[70][13] ), 
	.A(\ram[68][13] ));
   MUX4EHD U7284 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5825), 
	.D(\ram[67][13] ), 
	.C(\ram[65][13] ), 
	.B(\ram[66][13] ), 
	.A(\ram[64][13] ));
   MUX4EHD U7285 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5826), 
	.D(n5822), 
	.C(n5824), 
	.B(n5823), 
	.A(n5825));
   MUX4EHD U7286 (.S1(n6038), 
	.S0(n7444), 
	.O(n5827), 
	.D(n5811), 
	.C(n5821), 
	.B(n5816), 
	.A(n5826));
   MUX4EHD U7287 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5828), 
	.D(\ram[63][13] ), 
	.C(\ram[61][13] ), 
	.B(\ram[62][13] ), 
	.A(\ram[60][13] ));
   MUX4EHD U7288 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5829), 
	.D(\ram[59][13] ), 
	.C(\ram[57][13] ), 
	.B(\ram[58][13] ), 
	.A(\ram[56][13] ));
   MUX4EHD U7289 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5830), 
	.D(\ram[55][13] ), 
	.C(\ram[53][13] ), 
	.B(\ram[54][13] ), 
	.A(\ram[52][13] ));
   MUX4EHD U7290 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5831), 
	.D(\ram[51][13] ), 
	.C(\ram[49][13] ), 
	.B(\ram[50][13] ), 
	.A(\ram[48][13] ));
   MUX4EHD U7291 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5832), 
	.D(n5828), 
	.C(n5830), 
	.B(n5829), 
	.A(n5831));
   MUX4EHD U7292 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5833), 
	.D(\ram[47][13] ), 
	.C(\ram[45][13] ), 
	.B(\ram[46][13] ), 
	.A(\ram[44][13] ));
   MUX4EHD U7293 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5834), 
	.D(\ram[43][13] ), 
	.C(\ram[41][13] ), 
	.B(\ram[42][13] ), 
	.A(\ram[40][13] ));
   MUX4EHD U7294 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5835), 
	.D(\ram[39][13] ), 
	.C(\ram[37][13] ), 
	.B(\ram[38][13] ), 
	.A(\ram[36][13] ));
   MUX4EHD U7295 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5836), 
	.D(\ram[35][13] ), 
	.C(\ram[33][13] ), 
	.B(\ram[34][13] ), 
	.A(\ram[32][13] ));
   MUX4EHD U7296 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5837), 
	.D(n5833), 
	.C(n5835), 
	.B(n5834), 
	.A(n5836));
   MUX4EHD U7297 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5838), 
	.D(\ram[31][13] ), 
	.C(\ram[29][13] ), 
	.B(\ram[30][13] ), 
	.A(\ram[28][13] ));
   MUX4EHD U7298 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5839), 
	.D(\ram[27][13] ), 
	.C(\ram[25][13] ), 
	.B(\ram[26][13] ), 
	.A(\ram[24][13] ));
   MUX4EHD U7299 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5840), 
	.D(\ram[23][13] ), 
	.C(\ram[21][13] ), 
	.B(\ram[22][13] ), 
	.A(\ram[20][13] ));
   MUX4EHD U7300 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5841), 
	.D(\ram[19][13] ), 
	.C(\ram[17][13] ), 
	.B(\ram[18][13] ), 
	.A(\ram[16][13] ));
   MUX4EHD U7301 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5842), 
	.D(n5838), 
	.C(n5840), 
	.B(n5839), 
	.A(n5841));
   MUX4EHD U7302 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5843), 
	.D(\ram[15][13] ), 
	.C(\ram[13][13] ), 
	.B(\ram[14][13] ), 
	.A(\ram[12][13] ));
   MUX4EHD U7303 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5844), 
	.D(\ram[11][13] ), 
	.C(\ram[9][13] ), 
	.B(\ram[10][13] ), 
	.A(\ram[8][13] ));
   MUX4EHD U7304 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5845), 
	.D(\ram[7][13] ), 
	.C(\ram[5][13] ), 
	.B(\ram[6][13] ), 
	.A(\ram[4][13] ));
   MUX4EHD U7305 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5846), 
	.D(\ram[3][13] ), 
	.C(\ram[1][13] ), 
	.B(\ram[2][13] ), 
	.A(\ram[0][13] ));
   MUX4EHD U7306 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5847), 
	.D(n5843), 
	.C(n5845), 
	.B(n5844), 
	.A(n5846));
   MUX4EHD U7307 (.S1(n6038), 
	.S0(n7444), 
	.O(n5848), 
	.D(n5832), 
	.C(n5842), 
	.B(n5837), 
	.A(n5847));
   MUX4EHD U7308 (.S1(n6469), 
	.S0(n6470), 
	.O(N4128), 
	.D(n5785), 
	.C(n5827), 
	.B(n5806), 
	.A(n5848));
   MUX4EHD U7309 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5849), 
	.D(\ram[255][14] ), 
	.C(\ram[253][14] ), 
	.B(\ram[254][14] ), 
	.A(\ram[252][14] ));
   MUX4EHD U7310 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5850), 
	.D(\ram[251][14] ), 
	.C(\ram[249][14] ), 
	.B(\ram[250][14] ), 
	.A(\ram[248][14] ));
   MUX4EHD U7311 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5851), 
	.D(\ram[247][14] ), 
	.C(\ram[245][14] ), 
	.B(\ram[246][14] ), 
	.A(\ram[244][14] ));
   MUX4EHD U7312 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5852), 
	.D(\ram[243][14] ), 
	.C(\ram[241][14] ), 
	.B(\ram[242][14] ), 
	.A(\ram[240][14] ));
   MUX4EHD U7313 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5853), 
	.D(n5849), 
	.C(n5851), 
	.B(n5850), 
	.A(n5852));
   MUX4EHD U7314 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5854), 
	.D(\ram[239][14] ), 
	.C(\ram[237][14] ), 
	.B(\ram[238][14] ), 
	.A(\ram[236][14] ));
   MUX4EHD U7315 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5855), 
	.D(\ram[235][14] ), 
	.C(\ram[233][14] ), 
	.B(\ram[234][14] ), 
	.A(\ram[232][14] ));
   MUX4EHD U7316 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5856), 
	.D(\ram[231][14] ), 
	.C(\ram[229][14] ), 
	.B(\ram[230][14] ), 
	.A(\ram[228][14] ));
   MUX4EHD U7317 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5857), 
	.D(\ram[227][14] ), 
	.C(\ram[225][14] ), 
	.B(\ram[226][14] ), 
	.A(\ram[224][14] ));
   MUX4EHD U7318 (.S1(n6136), 
	.S0(n7442), 
	.O(n5858), 
	.D(n5854), 
	.C(n5856), 
	.B(n5855), 
	.A(n5857));
   MUX4EHD U7319 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5859), 
	.D(\ram[223][14] ), 
	.C(\ram[221][14] ), 
	.B(\ram[222][14] ), 
	.A(\ram[220][14] ));
   MUX4EHD U7320 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5860), 
	.D(\ram[219][14] ), 
	.C(\ram[217][14] ), 
	.B(\ram[218][14] ), 
	.A(\ram[216][14] ));
   MUX4EHD U7321 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5861), 
	.D(\ram[215][14] ), 
	.C(\ram[213][14] ), 
	.B(\ram[214][14] ), 
	.A(\ram[212][14] ));
   MUX4EHD U7322 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5862), 
	.D(\ram[211][14] ), 
	.C(\ram[209][14] ), 
	.B(\ram[210][14] ), 
	.A(\ram[208][14] ));
   MUX4EHD U7323 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5863), 
	.D(n5859), 
	.C(n5861), 
	.B(n5860), 
	.A(n5862));
   MUX4EHD U7324 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5864), 
	.D(\ram[207][14] ), 
	.C(\ram[205][14] ), 
	.B(\ram[206][14] ), 
	.A(\ram[204][14] ));
   MUX4EHD U7325 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5865), 
	.D(\ram[203][14] ), 
	.C(\ram[201][14] ), 
	.B(\ram[202][14] ), 
	.A(\ram[200][14] ));
   MUX4EHD U7326 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5866), 
	.D(\ram[199][14] ), 
	.C(\ram[197][14] ), 
	.B(\ram[198][14] ), 
	.A(\ram[196][14] ));
   MUX4EHD U7327 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5867), 
	.D(\ram[195][14] ), 
	.C(\ram[193][14] ), 
	.B(\ram[194][14] ), 
	.A(\ram[192][14] ));
   MUX4EHD U7328 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5868), 
	.D(n5864), 
	.C(n5866), 
	.B(n5865), 
	.A(n5867));
   MUX4EHD U7329 (.S1(n6038), 
	.S0(n7444), 
	.O(n5869), 
	.D(n5853), 
	.C(n5863), 
	.B(n5858), 
	.A(n5868));
   MUX4EHD U7330 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5870), 
	.D(\ram[191][14] ), 
	.C(\ram[189][14] ), 
	.B(\ram[190][14] ), 
	.A(\ram[188][14] ));
   MUX4EHD U7331 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5871), 
	.D(\ram[187][14] ), 
	.C(\ram[185][14] ), 
	.B(\ram[186][14] ), 
	.A(\ram[184][14] ));
   MUX4EHD U7332 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5872), 
	.D(\ram[183][14] ), 
	.C(\ram[181][14] ), 
	.B(\ram[182][14] ), 
	.A(\ram[180][14] ));
   MUX4EHD U7333 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5873), 
	.D(\ram[179][14] ), 
	.C(\ram[177][14] ), 
	.B(\ram[178][14] ), 
	.A(\ram[176][14] ));
   MUX4EHD U7334 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5874), 
	.D(n5870), 
	.C(n5872), 
	.B(n5871), 
	.A(n5873));
   MUX4EHD U7335 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5875), 
	.D(\ram[175][14] ), 
	.C(\ram[173][14] ), 
	.B(\ram[174][14] ), 
	.A(\ram[172][14] ));
   MUX4EHD U7336 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5876), 
	.D(\ram[171][14] ), 
	.C(\ram[169][14] ), 
	.B(\ram[170][14] ), 
	.A(\ram[168][14] ));
   MUX4EHD U7337 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5877), 
	.D(\ram[167][14] ), 
	.C(\ram[165][14] ), 
	.B(\ram[166][14] ), 
	.A(\ram[164][14] ));
   MUX4EHD U7338 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5878), 
	.D(\ram[163][14] ), 
	.C(\ram[161][14] ), 
	.B(\ram[162][14] ), 
	.A(\ram[160][14] ));
   MUX4EHD U7339 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5879), 
	.D(n5875), 
	.C(n5877), 
	.B(n5876), 
	.A(n5878));
   MUX4EHD U7340 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5880), 
	.D(\ram[159][14] ), 
	.C(\ram[157][14] ), 
	.B(\ram[158][14] ), 
	.A(\ram[156][14] ));
   MUX4EHD U7341 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5881), 
	.D(\ram[155][14] ), 
	.C(\ram[153][14] ), 
	.B(\ram[154][14] ), 
	.A(\ram[152][14] ));
   MUX4EHD U7342 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5882), 
	.D(\ram[151][14] ), 
	.C(\ram[149][14] ), 
	.B(\ram[150][14] ), 
	.A(\ram[148][14] ));
   MUX4EHD U7343 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5883), 
	.D(\ram[147][14] ), 
	.C(\ram[145][14] ), 
	.B(\ram[146][14] ), 
	.A(\ram[144][14] ));
   MUX4EHD U7344 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5884), 
	.D(n5880), 
	.C(n5882), 
	.B(n5881), 
	.A(n5883));
   MUX4EHD U7345 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5885), 
	.D(\ram[143][14] ), 
	.C(\ram[141][14] ), 
	.B(\ram[142][14] ), 
	.A(\ram[140][14] ));
   MUX4EHD U7346 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5886), 
	.D(\ram[139][14] ), 
	.C(\ram[137][14] ), 
	.B(\ram[138][14] ), 
	.A(\ram[136][14] ));
   MUX4EHD U7347 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5887), 
	.D(\ram[135][14] ), 
	.C(\ram[133][14] ), 
	.B(\ram[134][14] ), 
	.A(\ram[132][14] ));
   MUX4EHD U7348 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5888), 
	.D(\ram[131][14] ), 
	.C(\ram[129][14] ), 
	.B(\ram[130][14] ), 
	.A(\ram[128][14] ));
   MUX4EHD U7349 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5889), 
	.D(n5885), 
	.C(n5887), 
	.B(n5886), 
	.A(n5888));
   MUX4EHD U7350 (.S1(n6038), 
	.S0(n7444), 
	.O(n5890), 
	.D(n5874), 
	.C(n5884), 
	.B(n5879), 
	.A(n5889));
   MUX4EHD U7351 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5891), 
	.D(\ram[127][14] ), 
	.C(\ram[125][14] ), 
	.B(\ram[126][14] ), 
	.A(\ram[124][14] ));
   MUX4EHD U7352 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5892), 
	.D(\ram[123][14] ), 
	.C(\ram[121][14] ), 
	.B(\ram[122][14] ), 
	.A(\ram[120][14] ));
   MUX4EHD U7353 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5893), 
	.D(\ram[119][14] ), 
	.C(\ram[117][14] ), 
	.B(\ram[118][14] ), 
	.A(\ram[116][14] ));
   MUX4EHD U7354 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5894), 
	.D(\ram[115][14] ), 
	.C(\ram[113][14] ), 
	.B(\ram[114][14] ), 
	.A(\ram[112][14] ));
   MUX4EHD U7355 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5895), 
	.D(n5891), 
	.C(n5893), 
	.B(n5892), 
	.A(n5894));
   MUX4EHD U7356 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5896), 
	.D(\ram[111][14] ), 
	.C(\ram[109][14] ), 
	.B(\ram[110][14] ), 
	.A(\ram[108][14] ));
   MUX4EHD U7357 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5897), 
	.D(\ram[107][14] ), 
	.C(\ram[105][14] ), 
	.B(\ram[106][14] ), 
	.A(\ram[104][14] ));
   MUX4EHD U7358 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5898), 
	.D(\ram[103][14] ), 
	.C(\ram[101][14] ), 
	.B(\ram[102][14] ), 
	.A(\ram[100][14] ));
   MUX4EHD U7359 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5899), 
	.D(\ram[99][14] ), 
	.C(\ram[97][14] ), 
	.B(\ram[98][14] ), 
	.A(\ram[96][14] ));
   MUX4EHD U7360 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5900), 
	.D(n5896), 
	.C(n5898), 
	.B(n5897), 
	.A(n5899));
   MUX4EHD U7361 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5901), 
	.D(\ram[95][14] ), 
	.C(\ram[93][14] ), 
	.B(\ram[94][14] ), 
	.A(\ram[92][14] ));
   MUX4EHD U7362 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5902), 
	.D(\ram[91][14] ), 
	.C(\ram[89][14] ), 
	.B(\ram[90][14] ), 
	.A(\ram[88][14] ));
   MUX4EHD U7363 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5903), 
	.D(\ram[87][14] ), 
	.C(\ram[85][14] ), 
	.B(\ram[86][14] ), 
	.A(\ram[84][14] ));
   MUX4EHD U7364 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5904), 
	.D(\ram[83][14] ), 
	.C(\ram[81][14] ), 
	.B(\ram[82][14] ), 
	.A(\ram[80][14] ));
   MUX4EHD U7365 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5905), 
	.D(n5901), 
	.C(n5903), 
	.B(n5902), 
	.A(n5904));
   MUX4EHD U7366 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5906), 
	.D(\ram[79][14] ), 
	.C(\ram[77][14] ), 
	.B(\ram[78][14] ), 
	.A(\ram[76][14] ));
   MUX4EHD U7367 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5907), 
	.D(\ram[75][14] ), 
	.C(\ram[73][14] ), 
	.B(\ram[74][14] ), 
	.A(\ram[72][14] ));
   MUX4EHD U7368 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5908), 
	.D(\ram[71][14] ), 
	.C(\ram[69][14] ), 
	.B(\ram[70][14] ), 
	.A(\ram[68][14] ));
   MUX4EHD U7369 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5909), 
	.D(\ram[67][14] ), 
	.C(\ram[65][14] ), 
	.B(\ram[66][14] ), 
	.A(\ram[64][14] ));
   MUX4EHD U7370 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5910), 
	.D(n5906), 
	.C(n5908), 
	.B(n5907), 
	.A(n5909));
   MUX4EHD U7371 (.S1(n6038), 
	.S0(n7444), 
	.O(n5911), 
	.D(n5895), 
	.C(n5905), 
	.B(n5900), 
	.A(n5910));
   MUX4EHD U7372 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5912), 
	.D(\ram[63][14] ), 
	.C(\ram[61][14] ), 
	.B(\ram[62][14] ), 
	.A(\ram[60][14] ));
   MUX4EHD U7373 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5913), 
	.D(\ram[59][14] ), 
	.C(\ram[57][14] ), 
	.B(\ram[58][14] ), 
	.A(\ram[56][14] ));
   MUX4EHD U7374 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5914), 
	.D(\ram[55][14] ), 
	.C(\ram[53][14] ), 
	.B(\ram[54][14] ), 
	.A(\ram[52][14] ));
   MUX4EHD U7375 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5915), 
	.D(\ram[51][14] ), 
	.C(\ram[49][14] ), 
	.B(\ram[50][14] ), 
	.A(\ram[48][14] ));
   MUX4EHD U7376 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5916), 
	.D(n5912), 
	.C(n5914), 
	.B(n5913), 
	.A(n5915));
   MUX4EHD U7377 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5917), 
	.D(\ram[47][14] ), 
	.C(\ram[45][14] ), 
	.B(\ram[46][14] ), 
	.A(\ram[44][14] ));
   MUX4EHD U7378 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5918), 
	.D(\ram[43][14] ), 
	.C(\ram[41][14] ), 
	.B(\ram[42][14] ), 
	.A(\ram[40][14] ));
   MUX4EHD U7379 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5919), 
	.D(\ram[39][14] ), 
	.C(\ram[37][14] ), 
	.B(\ram[38][14] ), 
	.A(\ram[36][14] ));
   MUX4EHD U7380 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n5920), 
	.D(\ram[35][14] ), 
	.C(\ram[33][14] ), 
	.B(\ram[34][14] ), 
	.A(\ram[32][14] ));
   MUX4EHD U7381 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5921), 
	.D(n5917), 
	.C(n5919), 
	.B(n5918), 
	.A(n5920));
   MUX4EHD U7382 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5922), 
	.D(\ram[31][14] ), 
	.C(\ram[29][14] ), 
	.B(\ram[30][14] ), 
	.A(\ram[28][14] ));
   MUX4EHD U7383 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5923), 
	.D(\ram[27][14] ), 
	.C(\ram[25][14] ), 
	.B(\ram[26][14] ), 
	.A(\ram[24][14] ));
   MUX4EHD U7384 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5924), 
	.D(\ram[23][14] ), 
	.C(\ram[21][14] ), 
	.B(\ram[22][14] ), 
	.A(\ram[20][14] ));
   MUX4EHD U7385 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN12_n7440), 
	.O(n5925), 
	.D(\ram[19][14] ), 
	.C(\ram[17][14] ), 
	.B(\ram[18][14] ), 
	.A(\ram[16][14] ));
   MUX4EHD U7386 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5926), 
	.D(n5922), 
	.C(n5924), 
	.B(n5923), 
	.A(n5925));
   MUX4EHD U7387 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5927), 
	.D(\ram[15][14] ), 
	.C(\ram[13][14] ), 
	.B(\ram[14][14] ), 
	.A(\ram[12][14] ));
   MUX4EHD U7388 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5928), 
	.D(\ram[11][14] ), 
	.C(\ram[9][14] ), 
	.B(\ram[10][14] ), 
	.A(\ram[8][14] ));
   MUX4EHD U7389 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n5929), 
	.D(\ram[7][14] ), 
	.C(\ram[5][14] ), 
	.B(\ram[6][14] ), 
	.A(\ram[4][14] ));
   MUX4EHD U7390 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n5930), 
	.D(\ram[3][14] ), 
	.C(\ram[1][14] ), 
	.B(\ram[2][14] ), 
	.A(\ram[0][14] ));
   MUX4EHD U7391 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n5931), 
	.D(n5927), 
	.C(n5929), 
	.B(n5928), 
	.A(n5930));
   MUX4EHD U7392 (.S1(n6038), 
	.S0(n7444), 
	.O(n5932), 
	.D(n5916), 
	.C(n5926), 
	.B(n5921), 
	.A(n5931));
   MUX4EHD U7393 (.S1(n6469), 
	.S0(n6470), 
	.O(N4127), 
	.D(n5869), 
	.C(n5911), 
	.B(n5890), 
	.A(n5932));
   MUX4EHD U7394 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5933), 
	.D(\ram[255][15] ), 
	.C(\ram[253][15] ), 
	.B(\ram[254][15] ), 
	.A(\ram[252][15] ));
   MUX4EHD U7395 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5934), 
	.D(\ram[251][15] ), 
	.C(\ram[249][15] ), 
	.B(\ram[250][15] ), 
	.A(\ram[248][15] ));
   MUX4EHD U7396 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5935), 
	.D(\ram[247][15] ), 
	.C(\ram[245][15] ), 
	.B(\ram[246][15] ), 
	.A(\ram[244][15] ));
   MUX4EHD U7397 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5936), 
	.D(\ram[243][15] ), 
	.C(\ram[241][15] ), 
	.B(\ram[242][15] ), 
	.A(\ram[240][15] ));
   MUX4EHD U7398 (.S1(n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5937), 
	.D(n5933), 
	.C(n5935), 
	.B(n5934), 
	.A(n5936));
   MUX4EHD U7399 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5938), 
	.D(\ram[239][15] ), 
	.C(\ram[237][15] ), 
	.B(\ram[238][15] ), 
	.A(\ram[236][15] ));
   MUX4EHD U7400 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN7_n7440), 
	.O(n5939), 
	.D(\ram[235][15] ), 
	.C(\ram[233][15] ), 
	.B(\ram[234][15] ), 
	.A(\ram[232][15] ));
   MUX4EHD U7401 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5940), 
	.D(\ram[231][15] ), 
	.C(\ram[229][15] ), 
	.B(\ram[230][15] ), 
	.A(\ram[228][15] ));
   MUX4EHD U7402 (.S1(FE_OFN32_n6459), 
	.S0(FE_OFN11_n7440), 
	.O(n5941), 
	.D(\ram[227][15] ), 
	.C(\ram[225][15] ), 
	.B(\ram[226][15] ), 
	.A(\ram[224][15] ));
   MUX4EHD U7403 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5942), 
	.D(n5938), 
	.C(n5940), 
	.B(n5939), 
	.A(n5941));
   MUX4EHD U7404 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5943), 
	.D(\ram[223][15] ), 
	.C(\ram[221][15] ), 
	.B(\ram[222][15] ), 
	.A(\ram[220][15] ));
   MUX4EHD U7405 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5944), 
	.D(\ram[219][15] ), 
	.C(\ram[217][15] ), 
	.B(\ram[218][15] ), 
	.A(\ram[216][15] ));
   MUX4EHD U7406 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5945), 
	.D(\ram[215][15] ), 
	.C(\ram[213][15] ), 
	.B(\ram[214][15] ), 
	.A(\ram[212][15] ));
   MUX4EHD U7407 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5946), 
	.D(\ram[211][15] ), 
	.C(\ram[209][15] ), 
	.B(\ram[210][15] ), 
	.A(\ram[208][15] ));
   MUX4EHD U7408 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN1_n7442), 
	.O(n5947), 
	.D(n5943), 
	.C(n5945), 
	.B(n5944), 
	.A(n5946));
   MUX4EHD U7409 (.S1(FE_OFN31_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5948), 
	.D(\ram[207][15] ), 
	.C(\ram[205][15] ), 
	.B(\ram[206][15] ), 
	.A(\ram[204][15] ));
   MUX4EHD U7410 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5949), 
	.D(\ram[203][15] ), 
	.C(\ram[201][15] ), 
	.B(\ram[202][15] ), 
	.A(\ram[200][15] ));
   MUX4EHD U7411 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5950), 
	.D(\ram[199][15] ), 
	.C(\ram[197][15] ), 
	.B(\ram[198][15] ), 
	.A(\ram[196][15] ));
   MUX4EHD U7412 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5951), 
	.D(\ram[195][15] ), 
	.C(\ram[193][15] ), 
	.B(\ram[194][15] ), 
	.A(\ram[192][15] ));
   MUX4EHD U7413 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5952), 
	.D(n5948), 
	.C(n5950), 
	.B(n5949), 
	.A(n5951));
   MUX4EHD U7414 (.S1(n6038), 
	.S0(n7444), 
	.O(n5953), 
	.D(n5937), 
	.C(n5947), 
	.B(n5942), 
	.A(n5952));
   MUX4EHD U7415 (.S1(FE_OFN26_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5954), 
	.D(\ram[191][15] ), 
	.C(\ram[189][15] ), 
	.B(\ram[190][15] ), 
	.A(\ram[188][15] ));
   MUX4EHD U7416 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5955), 
	.D(\ram[187][15] ), 
	.C(\ram[185][15] ), 
	.B(\ram[186][15] ), 
	.A(\ram[184][15] ));
   MUX4EHD U7417 (.S1(FE_OFN26_n6459), 
	.S0(n7440), 
	.O(n5956), 
	.D(\ram[183][15] ), 
	.C(\ram[181][15] ), 
	.B(\ram[182][15] ), 
	.A(\ram[180][15] ));
   MUX4EHD U7418 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n5957), 
	.D(\ram[179][15] ), 
	.C(\ram[177][15] ), 
	.B(\ram[178][15] ), 
	.A(\ram[176][15] ));
   MUX4EHD U7419 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5958), 
	.D(n5954), 
	.C(n5956), 
	.B(n5955), 
	.A(n5957));
   MUX4EHD U7420 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5959), 
	.D(\ram[175][15] ), 
	.C(\ram[173][15] ), 
	.B(\ram[174][15] ), 
	.A(\ram[172][15] ));
   MUX4EHD U7421 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5960), 
	.D(\ram[171][15] ), 
	.C(\ram[169][15] ), 
	.B(\ram[170][15] ), 
	.A(\ram[168][15] ));
   MUX4EHD U7422 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN10_n7440), 
	.O(n5961), 
	.D(\ram[167][15] ), 
	.C(\ram[165][15] ), 
	.B(\ram[166][15] ), 
	.A(\ram[164][15] ));
   MUX4EHD U7423 (.S1(FE_OFN27_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5962), 
	.D(\ram[163][15] ), 
	.C(\ram[161][15] ), 
	.B(\ram[162][15] ), 
	.A(\ram[160][15] ));
   MUX4EHD U7424 (.S1(FE_OFN22_n6136), 
	.S0(n7442), 
	.O(n5963), 
	.D(n5959), 
	.C(n5961), 
	.B(n5960), 
	.A(n5962));
   MUX4EHD U7425 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5964), 
	.D(\ram[159][15] ), 
	.C(\ram[157][15] ), 
	.B(\ram[158][15] ), 
	.A(\ram[156][15] ));
   MUX4EHD U7426 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5965), 
	.D(\ram[155][15] ), 
	.C(\ram[153][15] ), 
	.B(\ram[154][15] ), 
	.A(\ram[152][15] ));
   MUX4EHD U7427 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n5966), 
	.D(\ram[151][15] ), 
	.C(\ram[149][15] ), 
	.B(\ram[150][15] ), 
	.A(\ram[148][15] ));
   MUX4EHD U7428 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN6_n7440), 
	.O(n5967), 
	.D(\ram[147][15] ), 
	.C(\ram[145][15] ), 
	.B(\ram[146][15] ), 
	.A(\ram[144][15] ));
   MUX4EHD U7429 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5968), 
	.D(n5964), 
	.C(n5966), 
	.B(n5965), 
	.A(n5967));
   MUX4EHD U7430 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5969), 
	.D(\ram[143][15] ), 
	.C(\ram[141][15] ), 
	.B(\ram[142][15] ), 
	.A(\ram[140][15] ));
   MUX4EHD U7431 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5970), 
	.D(\ram[139][15] ), 
	.C(\ram[137][15] ), 
	.B(\ram[138][15] ), 
	.A(\ram[136][15] ));
   MUX4EHD U7432 (.S1(FE_OFN25_n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5971), 
	.D(\ram[135][15] ), 
	.C(\ram[133][15] ), 
	.B(\ram[134][15] ), 
	.A(\ram[132][15] ));
   MUX4EHD U7433 (.S1(n6459), 
	.S0(FE_OFN8_n7440), 
	.O(n5972), 
	.D(\ram[131][15] ), 
	.C(\ram[129][15] ), 
	.B(\ram[130][15] ), 
	.A(\ram[128][15] ));
   MUX4EHD U7434 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN0_n7442), 
	.O(n5973), 
	.D(n5969), 
	.C(n5971), 
	.B(n5970), 
	.A(n5972));
   MUX4EHD U7435 (.S1(n6038), 
	.S0(n7444), 
	.O(n5974), 
	.D(n5958), 
	.C(n5968), 
	.B(n5963), 
	.A(n5973));
   MUX4EHD U7436 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5975), 
	.D(\ram[127][15] ), 
	.C(\ram[125][15] ), 
	.B(\ram[126][15] ), 
	.A(\ram[124][15] ));
   MUX4EHD U7437 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5976), 
	.D(\ram[123][15] ), 
	.C(\ram[121][15] ), 
	.B(\ram[122][15] ), 
	.A(\ram[120][15] ));
   MUX4EHD U7438 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5977), 
	.D(\ram[119][15] ), 
	.C(\ram[117][15] ), 
	.B(\ram[118][15] ), 
	.A(\ram[116][15] ));
   MUX4EHD U7439 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5978), 
	.D(\ram[115][15] ), 
	.C(\ram[113][15] ), 
	.B(\ram[114][15] ), 
	.A(\ram[112][15] ));
   MUX4EHD U7440 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5979), 
	.D(n5975), 
	.C(n5977), 
	.B(n5976), 
	.A(n5978));
   MUX4EHD U7441 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5980), 
	.D(\ram[111][15] ), 
	.C(\ram[109][15] ), 
	.B(\ram[110][15] ), 
	.A(\ram[108][15] ));
   MUX4EHD U7442 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN14_n7440), 
	.O(n5981), 
	.D(\ram[107][15] ), 
	.C(\ram[105][15] ), 
	.B(\ram[106][15] ), 
	.A(\ram[104][15] ));
   MUX4EHD U7443 (.S1(FE_OFN40_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5982), 
	.D(\ram[103][15] ), 
	.C(\ram[101][15] ), 
	.B(\ram[102][15] ), 
	.A(\ram[100][15] ));
   MUX4EHD U7444 (.S1(FE_OFN36_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n5983), 
	.D(\ram[99][15] ), 
	.C(\ram[97][15] ), 
	.B(\ram[98][15] ), 
	.A(\ram[96][15] ));
   MUX4EHD U7445 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5984), 
	.D(n5980), 
	.C(n5982), 
	.B(n5981), 
	.A(n5983));
   MUX4EHD U7446 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN9_n7440), 
	.O(n5985), 
	.D(\ram[95][15] ), 
	.C(\ram[93][15] ), 
	.B(\ram[94][15] ), 
	.A(\ram[92][15] ));
   MUX4EHD U7447 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5986), 
	.D(\ram[91][15] ), 
	.C(\ram[89][15] ), 
	.B(\ram[90][15] ), 
	.A(\ram[88][15] ));
   MUX4EHD U7448 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN21_n7440), 
	.O(n5987), 
	.D(\ram[87][15] ), 
	.C(\ram[85][15] ), 
	.B(\ram[86][15] ), 
	.A(\ram[84][15] ));
   MUX4EHD U7449 (.S1(FE_OFN37_n6459), 
	.S0(FE_OFN20_n7440), 
	.O(n5988), 
	.D(\ram[83][15] ), 
	.C(\ram[81][15] ), 
	.B(\ram[82][15] ), 
	.A(\ram[80][15] ));
   MUX4EHD U7450 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n5989), 
	.D(n5985), 
	.C(n5987), 
	.B(n5986), 
	.A(n5988));
   MUX4EHD U7451 (.S1(FE_OFN33_n6459), 
	.S0(FE_OFN13_n7440), 
	.O(n5990), 
	.D(\ram[79][15] ), 
	.C(\ram[77][15] ), 
	.B(\ram[78][15] ), 
	.A(\ram[76][15] ));
   MUX4EHD U7452 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5991), 
	.D(\ram[75][15] ), 
	.C(\ram[73][15] ), 
	.B(\ram[74][15] ), 
	.A(\ram[72][15] ));
   MUX4EHD U7453 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5992), 
	.D(\ram[71][15] ), 
	.C(\ram[69][15] ), 
	.B(\ram[70][15] ), 
	.A(\ram[68][15] ));
   MUX4EHD U7454 (.S1(FE_OFN38_n6459), 
	.S0(FE_OFN19_n7440), 
	.O(n5993), 
	.D(\ram[67][15] ), 
	.C(\ram[65][15] ), 
	.B(\ram[66][15] ), 
	.A(\ram[64][15] ));
   MUX4EHD U7455 (.S1(FE_OFN23_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n5994), 
	.D(n5990), 
	.C(n5992), 
	.B(n5991), 
	.A(n5993));
   MUX4EHD U7456 (.S1(n6038), 
	.S0(n7444), 
	.O(n5995), 
	.D(n5979), 
	.C(n5989), 
	.B(n5984), 
	.A(n5994));
   MUX4EHD U7457 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5996), 
	.D(\ram[63][15] ), 
	.C(\ram[61][15] ), 
	.B(\ram[62][15] ), 
	.A(\ram[60][15] ));
   MUX4EHD U7458 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5997), 
	.D(\ram[59][15] ), 
	.C(\ram[57][15] ), 
	.B(\ram[58][15] ), 
	.A(\ram[56][15] ));
   MUX4EHD U7459 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5998), 
	.D(\ram[55][15] ), 
	.C(\ram[53][15] ), 
	.B(\ram[54][15] ), 
	.A(\ram[52][15] ));
   MUX4EHD U7460 (.S1(FE_OFN39_n6459), 
	.S0(FE_OFN15_n7440), 
	.O(n5999), 
	.D(\ram[51][15] ), 
	.C(\ram[49][15] ), 
	.B(\ram[50][15] ), 
	.A(\ram[48][15] ));
   MUX4EHD U7461 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN4_n7442), 
	.O(n6000), 
	.D(n5996), 
	.C(n5998), 
	.B(n5997), 
	.A(n5999));
   MUX4EHD U7462 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6001), 
	.D(\ram[47][15] ), 
	.C(\ram[45][15] ), 
	.B(\ram[46][15] ), 
	.A(\ram[44][15] ));
   MUX4EHD U7463 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6002), 
	.D(\ram[43][15] ), 
	.C(\ram[41][15] ), 
	.B(\ram[42][15] ), 
	.A(\ram[40][15] ));
   MUX4EHD U7464 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6003), 
	.D(\ram[39][15] ), 
	.C(\ram[37][15] ), 
	.B(\ram[38][15] ), 
	.A(\ram[36][15] ));
   MUX4EHD U7465 (.S1(FE_OFN35_n6459), 
	.S0(FE_OFN16_n7440), 
	.O(n6004), 
	.D(\ram[35][15] ), 
	.C(\ram[33][15] ), 
	.B(\ram[34][15] ), 
	.A(\ram[32][15] ));
   MUX4EHD U7466 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n6005), 
	.D(n6001), 
	.C(n6003), 
	.B(n6002), 
	.A(n6004));
   MUX4EHD U7467 (.S1(FE_OFN30_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n6006), 
	.D(\ram[31][15] ), 
	.C(\ram[29][15] ), 
	.B(\ram[30][15] ), 
	.A(\ram[28][15] ));
   MUX4EHD U7468 (.S1(FE_OFN28_n6459), 
	.S0(FE_OFN5_n7440), 
	.O(n6007), 
	.D(\ram[27][15] ), 
	.C(\ram[25][15] ), 
	.B(\ram[26][15] ), 
	.A(\ram[24][15] ));
   MUX4EHD U7469 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n6008), 
	.D(\ram[23][15] ), 
	.C(\ram[21][15] ), 
	.B(\ram[22][15] ), 
	.A(\ram[20][15] ));
   MUX4EHD U7470 (.S1(FE_OFN34_n6459), 
	.S0(FE_OFN18_n7440), 
	.O(n6009), 
	.D(\ram[19][15] ), 
	.C(\ram[17][15] ), 
	.B(\ram[18][15] ), 
	.A(\ram[16][15] ));
   MUX4EHD U7471 (.S1(FE_OFN24_n6136), 
	.S0(FE_OFN2_n7442), 
	.O(n6010), 
	.D(n6006), 
	.C(n6008), 
	.B(n6007), 
	.A(n6009));
   MUX4EHD U7472 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n6011), 
	.D(\ram[15][15] ), 
	.C(\ram[13][15] ), 
	.B(\ram[14][15] ), 
	.A(\ram[12][15] ));
   MUX4EHD U7473 (.S1(FE_OFN29_n6459), 
	.S0(FE_OFN17_n7440), 
	.O(n6012), 
	.D(\ram[11][15] ), 
	.C(\ram[9][15] ), 
	.B(\ram[10][15] ), 
	.A(\ram[8][15] ));
   MUX4EHD U7474 (.S1(FE_OFN35_n6459), 
	.S0(n7440), 
	.O(n6013), 
	.D(\ram[7][15] ), 
	.C(\ram[5][15] ), 
	.B(\ram[6][15] ), 
	.A(\ram[4][15] ));
   MUX4EHD U7475 (.S1(FE_OFN29_n6459), 
	.S0(n7440), 
	.O(n6014), 
	.D(\ram[3][15] ), 
	.C(\ram[1][15] ), 
	.B(\ram[2][15] ), 
	.A(\ram[0][15] ));
   MUX4EHD U7476 (.S1(FE_OFN22_n6136), 
	.S0(FE_OFN3_n7442), 
	.O(n6015), 
	.D(n6011), 
	.C(n6013), 
	.B(n6012), 
	.A(n6014));
   MUX4EHD U7477 (.S1(n6038), 
	.S0(n7444), 
	.O(n6016), 
	.D(n6000), 
	.C(n6010), 
	.B(n6005), 
	.A(n6015));
   MUX4EHD U7478 (.S1(n6469), 
	.S0(n6470), 
	.O(N4126), 
	.D(n5953), 
	.C(n5995), 
	.B(n5974), 
	.A(n6016));
endmodule

module alu (
	a, 
	b, 
	alu_control, 
	result, 
	zero);
   input [15:0] a;
   input [15:0] b;
   input [2:0] alu_control;
   output [15:0] result;
   output zero;

   // Internal wires
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N46;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N90;
   wire n10;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;

   OR3B1EHD U19 (.O(n31), 
	.I2(result[14]), 
	.I1(result[13]), 
	.B1(n44));
   NR6EHD U69 (.O(zero), 
	.I6(result[0]), 
	.I5(result[10]), 
	.I4(result[11]), 
	.I3(result[12]), 
	.I2(n31), 
	.I1(n74));
   NR8EHD U70 (.O(n49), 
	.I8(result[9]), 
	.I7(result[8]), 
	.I6(result[7]), 
	.I5(result[6]), 
	.I4(result[5]), 
	.I3(result[4]), 
	.I2(result[3]), 
	.I1(result[2]));
   alu_DW01_sub_0 sub_14 (.A({ a[15],
		a[14],
		a[13],
		a[12],
		a[11],
		a[10],
		a[9],
		a[8],
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }), 
	.B({ b[15],
		b[14],
		b[13],
		b[12],
		b[11],
		b[10],
		b[9],
		b[8],
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }), 
	.CI(n10), 
	.DIFF({ N57,
		N56,
		N55,
		N54,
		N53,
		N52,
		N51,
		N50,
		N49,
		N48,
		N47,
		N46,
		N45,
		N44,
		N43,
		N42 }));
   alu_DW01_add_0 r53 (.A({ a[15],
		a[14],
		a[13],
		a[12],
		a[11],
		a[10],
		a[9],
		a[8],
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }), 
	.B({ b[15],
		b[14],
		b[13],
		b[12],
		b[11],
		b[10],
		b[9],
		b[8],
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }), 
	.CI(n10), 
	.SUM({ N41,
		N40,
		N39,
		N38,
		N37,
		N36,
		N35,
		N34,
		N33,
		N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26 }));
   XNR2EHD U2 (.O(n35), 
	.I2(n37), 
	.I1(n80));
   INVDHD U3 (.O(n79), 
	.I(n32));
   NR2CHD U4 (.O(n44), 
	.I2(result[15]), 
	.I1(result[1]));
   AO2222EHD U5 (.O(result[9]), 
	.D2(n50), 
	.D1(b[9]), 
	.C2(n35), 
	.C1(N35), 
	.B2(a[9]), 
	.B1(n79), 
	.A2(n40), 
	.A1(N51));
   OAI12CHD U6 (.O(n50), 
	.B2(n64), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U7 (.O(result[15]), 
	.D2(n45), 
	.D1(b[15]), 
	.C2(n35), 
	.C1(N41), 
	.B2(n79), 
	.B1(a[15]), 
	.A2(n40), 
	.A1(N57));
   OAI12CHD U8 (.O(n45), 
	.B2(n73), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U9 (.O(result[13]), 
	.D2(n48), 
	.D1(b[13]), 
	.C2(n35), 
	.C1(N39), 
	.B2(n79), 
	.B1(a[13]), 
	.A2(n40), 
	.A1(N55));
   OAI12CHD U10 (.O(n48), 
	.B2(n70), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U11 (.O(result[11]), 
	.D2(n42), 
	.D1(b[11]), 
	.C2(n35), 
	.C1(N37), 
	.B2(n79), 
	.B1(a[11]), 
	.A2(n40), 
	.A1(N53));
   OAI12CHD U12 (.O(n42), 
	.B2(n67), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U13 (.O(result[14]), 
	.D2(n47), 
	.D1(b[14]), 
	.C2(n35), 
	.C1(N40), 
	.B2(n79), 
	.B1(a[14]), 
	.A2(n40), 
	.A1(N56));
   OAI12CHD U14 (.O(n47), 
	.B2(n75), 
	.B1(n39), 
	.A1(n32));
   INVDHD U15 (.O(n75), 
	.I(a[14]));
   AO2222CHD U16 (.O(result[12]), 
	.D2(n43), 
	.D1(b[12]), 
	.C2(n35), 
	.C1(N38), 
	.B2(n79), 
	.B1(a[12]), 
	.A2(n40), 
	.A1(N54));
   OAI12CHD U17 (.O(n43), 
	.B2(n69), 
	.B1(n39), 
	.A1(n32));
   INVDHD U18 (.O(n29), 
	.I(b[4]));
   INVDHD U20 (.O(n30), 
	.I(a[4]));
   INVDHD U21 (.O(n59), 
	.I(b[6]));
   INVDHD U22 (.O(n60), 
	.I(a[6]));
   INVDHD U23 (.O(n62), 
	.I(b[8]));
   INVDHD U24 (.O(n63), 
	.I(a[8]));
   INVDHD U25 (.O(n65), 
	.I(b[10]));
   INVDHD U26 (.O(n66), 
	.I(a[10]));
   INVDHD U27 (.O(n68), 
	.I(b[12]));
   INVDHD U28 (.O(n69), 
	.I(a[12]));
   INVDHD U29 (.O(n27), 
	.I(b[2]));
   INVDHD U30 (.O(n26), 
	.I(b[1]));
   INVDHD U31 (.O(n71), 
	.I(b[14]));
   AN2EHD U32 (.O(n36), 
	.I2(alu_control[2]), 
	.I1(N90));
   INVDHD U33 (.O(n72), 
	.I(b[15]));
   OAI112BHD U34 (.O(result[0]), 
	.C2(n78), 
	.C1(n32), 
	.B1(n34), 
	.A1(n33));
   ND2DHD U35 (.O(n33), 
	.I2(n40), 
	.I1(N42));
   AOI222BHD U36 (.O(n34), 
	.C2(n38), 
	.C1(b[0]), 
	.B2(n37), 
	.B1(n36), 
	.A2(n35), 
	.A1(N26));
   OAI12CHD U37 (.O(n38), 
	.B2(n78), 
	.B1(n39), 
	.A1(n32));
   AO2222EHD U38 (.O(result[8]), 
	.D2(n51), 
	.D1(b[8]), 
	.C2(n35), 
	.C1(N34), 
	.B2(n79), 
	.B1(a[8]), 
	.A2(n40), 
	.A1(N50));
   OAI12CHD U39 (.O(n51), 
	.B2(n63), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U40 (.O(result[10]), 
	.D2(n41), 
	.D1(b[10]), 
	.C2(n35), 
	.C1(N36), 
	.B2(n79), 
	.B1(a[10]), 
	.A2(n40), 
	.A1(N52));
   OAI12CHD U41 (.O(n41), 
	.B2(n66), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U42 (.O(result[7]), 
	.D2(n52), 
	.D1(b[7]), 
	.C2(n35), 
	.C1(N33), 
	.B2(n79), 
	.B1(a[7]), 
	.A2(n40), 
	.A1(N49));
   OAI12CHD U43 (.O(n52), 
	.B2(n61), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U44 (.O(result[6]), 
	.D2(n53), 
	.D1(b[6]), 
	.C2(n35), 
	.C1(N32), 
	.B2(n79), 
	.B1(a[6]), 
	.A2(n40), 
	.A1(N48));
   OAI12CHD U45 (.O(n53), 
	.B2(n60), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U46 (.O(result[1]), 
	.D2(n46), 
	.D1(b[1]), 
	.C2(n35), 
	.C1(N27), 
	.B2(n79), 
	.B1(a[1]), 
	.A2(n40), 
	.A1(N43));
   OAI12CHD U47 (.O(n46), 
	.B2(n77), 
	.B1(n39), 
	.A1(n32));
   INVDHD U48 (.O(n77), 
	.I(a[1]));
   ND3CHD U49 (.O(n32), 
	.I3(alu_control[0]), 
	.I2(n80), 
	.I1(alu_control[1]));
   AO2222CHD U50 (.O(result[5]), 
	.D2(n54), 
	.D1(b[5]), 
	.C2(n35), 
	.C1(N31), 
	.B2(n79), 
	.B1(a[5]), 
	.A2(n40), 
	.A1(N47));
   OAI12CHD U51 (.O(n54), 
	.B2(n58), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U52 (.O(result[3]), 
	.D2(n56), 
	.D1(b[3]), 
	.C2(n35), 
	.C1(N29), 
	.B2(n79), 
	.B1(a[3]), 
	.A2(n40), 
	.A1(N45));
   OAI12CHD U53 (.O(n56), 
	.B2(n28), 
	.B1(n39), 
	.A1(n32));
   AO2222CHD U54 (.O(result[4]), 
	.D2(n55), 
	.D1(b[4]), 
	.C2(n35), 
	.C1(N30), 
	.B2(n79), 
	.B1(a[4]), 
	.A2(n40), 
	.A1(N46));
   OAI12CHD U55 (.O(n55), 
	.B2(n30), 
	.B1(n39), 
	.A1(n32));
   ND2DHD U56 (.O(n39), 
	.I2(n80), 
	.I1(alu_control[1]));
   NR2CHD U57 (.O(n37), 
	.I2(alu_control[0]), 
	.I1(alu_control[1]));
   INVDHD U58 (.O(n80), 
	.I(alu_control[2]));
   AN3B2BHD U60 (.O(n40), 
	.I1(alu_control[0]), 
	.B2(alu_control[2]), 
	.B1(alu_control[1]));
   AO2222CHD U61 (.O(result[2]), 
	.D2(n57), 
	.D1(b[2]), 
	.C2(n35), 
	.C1(N28), 
	.B2(n79), 
	.B1(a[2]), 
	.A2(n40), 
	.A1(N44));
   OAI12CHD U62 (.O(n57), 
	.B2(n76), 
	.B1(n39), 
	.A1(n32));
   INVDHD U63 (.O(n76), 
	.I(a[2]));
   INVDHD U64 (.O(n74), 
	.I(n49));
   INVDHD U65 (.O(n28), 
	.I(a[3]));
   INVDHD U66 (.O(n58), 
	.I(a[5]));
   INVDHD U67 (.O(n64), 
	.I(a[9]));
   INVDHD U68 (.O(n61), 
	.I(a[7]));
   INVDHD U71 (.O(n67), 
	.I(a[11]));
   INVDHD U72 (.O(n70), 
	.I(a[13]));
   INVDHD U73 (.O(n78), 
	.I(a[0]));
   INVDHD U74 (.O(n73), 
	.I(a[15]));
   TIE0DHD U75 (.O(n10));
   AN2CHD U76 (.O(n22), 
	.I2(b[13]), 
	.I1(n70));
   AN2CHD U77 (.O(n19), 
	.I2(b[11]), 
	.I1(n67));
   AN2CHD U78 (.O(n16), 
	.I2(b[9]), 
	.I1(n64));
   AN2CHD U79 (.O(n13), 
	.I2(b[7]), 
	.I1(n61));
   AN2CHD U80 (.O(n9), 
	.I2(b[5]), 
	.I1(n58));
   AN2CHD U81 (.O(n6), 
	.I2(b[3]), 
	.I1(n28));
   OR2B1CHD U82 (.O(n3), 
	.I1(a[0]), 
	.B1(b[0]));
   OR2CHD U83 (.O(n2), 
	.I2(n3), 
	.I1(a[1]));
   AO222CHD U84 (.O(n4), 
	.C2(a[2]), 
	.C1(n27), 
	.B2(n2), 
	.B1(n26), 
	.A2(a[1]), 
	.A1(n3));
   OAI12CHD U85 (.O(n5), 
	.B2(n27), 
	.B1(a[2]), 
	.A1(n4));
   OAI222BHD U86 (.O(n7), 
	.C2(n30), 
	.C1(b[4]), 
	.B2(n5), 
	.B1(n6), 
	.A2(n28), 
	.A1(b[3]));
   OAI12CHD U87 (.O(n8), 
	.B2(n29), 
	.B1(a[4]), 
	.A1(n7));
   OAI222BHD U88 (.O(n11), 
	.C2(n60), 
	.C1(b[6]), 
	.B2(n8), 
	.B1(n9), 
	.A2(n58), 
	.A1(b[5]));
   OAI12CHD U89 (.O(n12), 
	.B2(n59), 
	.B1(a[6]), 
	.A1(n11));
   OAI222BHD U90 (.O(n14), 
	.C2(n63), 
	.C1(b[8]), 
	.B2(n12), 
	.B1(n13), 
	.A2(n61), 
	.A1(b[7]));
   OAI12CHD U91 (.O(n15), 
	.B2(n62), 
	.B1(a[8]), 
	.A1(n14));
   OAI222BHD U92 (.O(n17), 
	.C2(n64), 
	.C1(b[9]), 
	.B2(n15), 
	.B1(n16), 
	.A2(n66), 
	.A1(b[10]));
   OAI12CHD U93 (.O(n18), 
	.B2(n65), 
	.B1(a[10]), 
	.A1(n17));
   OAI222BHD U94 (.O(n20), 
	.C2(n69), 
	.C1(b[12]), 
	.B2(n18), 
	.B1(n19), 
	.A2(n67), 
	.A1(b[11]));
   OAI12CHD U95 (.O(n21), 
	.B2(n68), 
	.B1(a[12]), 
	.A1(n20));
   OAI222BHD U96 (.O(n23), 
	.C2(n75), 
	.C1(b[14]), 
	.B2(n21), 
	.B1(n22), 
	.A2(n70), 
	.A1(b[13]));
   OAI12CHD U97 (.O(n24), 
	.B2(n71), 
	.B1(a[14]), 
	.A1(n23));
   OAI12CHD U98 (.O(n25), 
	.B2(n73), 
	.B1(b[15]), 
	.A1(n24));
   OAI12CHD U99 (.O(N90), 
	.B2(n72), 
	.B1(a[15]), 
	.A1(n25));
endmodule

module ALUControl (
	ALU_Control, 
	ALUOp, 
	Function);
   output [2:0] ALU_Control;
   input [1:0] ALUOp;
   input [3:0] Function;

   // Internal wires
   wire N9;
   wire N15;
   wire N20;
   wire n3;
   wire n4;
   wire n5;
   wire n1;
   wire n2;

   assign ALU_Control[2] = N9 ;
   assign ALU_Control[1] = N15 ;
   assign ALU_Control[0] = N20 ;

   OAI22CHD U8 (.O(N20), 
	.B2(n2), 
	.B1(n5), 
	.A2(n1), 
	.A1(ALUOp[1]));
   INVDHD U1 (.O(n1), 
	.I(ALUOp[0]));
   AN3B2BHD U2 (.O(N15), 
	.I1(Function[1]), 
	.B2(n5), 
	.B1(ALUOp[0]));
   NR2CHD U3 (.O(N9), 
	.I2(n3), 
	.I1(ALUOp[0]));
   AOI13BHD U4 (.O(n3), 
	.B3(n4), 
	.B2(n2), 
	.B1(Function[2]), 
	.A1(ALUOp[1]));
   NR2CHD U5 (.O(n4), 
	.I2(Function[1]), 
	.I1(Function[3]));
   OR3EHD U6 (.O(n5), 
	.I3(ALUOp[1]), 
	.I2(Function[3]), 
	.I1(Function[2]));
   INVDHD U7 (.O(n2), 
	.I(Function[0]));
endmodule

module JR_Control (
	alu_op, 
	funct, 
	JRControl);
   input [1:0] alu_op;
   input [3:0] funct;
   output JRControl;

   // Internal wires
   wire n1;

   NR6EHD U2 (.O(JRControl), 
	.I6(alu_op[0]), 
	.I5(alu_op[1]), 
	.I4(n1), 
	.I3(funct[1]), 
	.I2(funct[2]), 
	.I1(funct[0]));
   INVDHD U1 (.O(n1), 
	.I(funct[3]));
endmodule

module register_file (
	clk, 
	rst, 
	reg_write_en, 
	reg_write_dest, 
	reg_write_data, 
	reg_read_addr_1, 
	reg_read_data_1, 
	reg_read_addr_2, 
	reg_read_data_2, 
	clk_m__L3_N123, 
	clk_m__L3_N124, 
	clk_m__L3_N126, 
	clk_m__L3_N154, 
	clk_m__L3_N49, 
	clk_m__L3_N50, 
	clk_m__L3_N51, 
	clk_m__L3_N53, 
	clk_m__L3_N54, 
	clk_m__L3_N80);
   input clk;
   input rst;
   input reg_write_en;
   input [2:0] reg_write_dest;
   input [15:0] reg_write_data;
   input [2:0] reg_read_addr_1;
   output [15:0] reg_read_data_1;
   input [2:0] reg_read_addr_2;
   output [15:0] reg_read_data_2;
   input clk_m__L3_N123;
   input clk_m__L3_N124;
   input clk_m__L3_N126;
   input clk_m__L3_N154;
   input clk_m__L3_N49;
   input clk_m__L3_N50;
   input clk_m__L3_N51;
   input clk_m__L3_N53;
   input clk_m__L3_N54;
   input clk_m__L3_N80;

   // Internal wires
   wire FE_OFN95_n240;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire \reg_array[7][15] ;
   wire \reg_array[7][14] ;
   wire \reg_array[7][13] ;
   wire \reg_array[7][12] ;
   wire \reg_array[7][11] ;
   wire \reg_array[7][10] ;
   wire \reg_array[7][9] ;
   wire \reg_array[7][8] ;
   wire \reg_array[7][7] ;
   wire \reg_array[7][6] ;
   wire \reg_array[7][5] ;
   wire \reg_array[7][4] ;
   wire \reg_array[7][3] ;
   wire \reg_array[7][2] ;
   wire \reg_array[7][1] ;
   wire \reg_array[7][0] ;
   wire \reg_array[6][15] ;
   wire \reg_array[6][14] ;
   wire \reg_array[6][13] ;
   wire \reg_array[6][12] ;
   wire \reg_array[6][11] ;
   wire \reg_array[6][10] ;
   wire \reg_array[6][9] ;
   wire \reg_array[6][8] ;
   wire \reg_array[6][7] ;
   wire \reg_array[6][6] ;
   wire \reg_array[6][5] ;
   wire \reg_array[6][4] ;
   wire \reg_array[6][3] ;
   wire \reg_array[6][2] ;
   wire \reg_array[6][1] ;
   wire \reg_array[6][0] ;
   wire \reg_array[5][15] ;
   wire \reg_array[5][14] ;
   wire \reg_array[5][13] ;
   wire \reg_array[5][12] ;
   wire \reg_array[5][11] ;
   wire \reg_array[5][10] ;
   wire \reg_array[5][9] ;
   wire \reg_array[5][8] ;
   wire \reg_array[5][7] ;
   wire \reg_array[5][6] ;
   wire \reg_array[5][5] ;
   wire \reg_array[5][4] ;
   wire \reg_array[5][3] ;
   wire \reg_array[5][2] ;
   wire \reg_array[5][1] ;
   wire \reg_array[5][0] ;
   wire \reg_array[4][15] ;
   wire \reg_array[4][14] ;
   wire \reg_array[4][13] ;
   wire \reg_array[4][12] ;
   wire \reg_array[4][11] ;
   wire \reg_array[4][10] ;
   wire \reg_array[4][9] ;
   wire \reg_array[4][8] ;
   wire \reg_array[4][7] ;
   wire \reg_array[4][6] ;
   wire \reg_array[4][5] ;
   wire \reg_array[4][4] ;
   wire \reg_array[4][3] ;
   wire \reg_array[4][2] ;
   wire \reg_array[4][1] ;
   wire \reg_array[4][0] ;
   wire \reg_array[3][15] ;
   wire \reg_array[3][14] ;
   wire \reg_array[3][13] ;
   wire \reg_array[3][12] ;
   wire \reg_array[3][11] ;
   wire \reg_array[3][10] ;
   wire \reg_array[3][9] ;
   wire \reg_array[3][8] ;
   wire \reg_array[3][7] ;
   wire \reg_array[3][6] ;
   wire \reg_array[3][5] ;
   wire \reg_array[3][4] ;
   wire \reg_array[3][3] ;
   wire \reg_array[3][2] ;
   wire \reg_array[3][1] ;
   wire \reg_array[3][0] ;
   wire \reg_array[2][15] ;
   wire \reg_array[2][14] ;
   wire \reg_array[2][13] ;
   wire \reg_array[2][12] ;
   wire \reg_array[2][11] ;
   wire \reg_array[2][10] ;
   wire \reg_array[2][9] ;
   wire \reg_array[2][8] ;
   wire \reg_array[2][7] ;
   wire \reg_array[2][6] ;
   wire \reg_array[2][5] ;
   wire \reg_array[2][4] ;
   wire \reg_array[2][3] ;
   wire \reg_array[2][2] ;
   wire \reg_array[2][1] ;
   wire \reg_array[2][0] ;
   wire \reg_array[1][15] ;
   wire \reg_array[1][14] ;
   wire \reg_array[1][13] ;
   wire \reg_array[1][12] ;
   wire \reg_array[1][11] ;
   wire \reg_array[1][10] ;
   wire \reg_array[1][9] ;
   wire \reg_array[1][8] ;
   wire \reg_array[1][7] ;
   wire \reg_array[1][6] ;
   wire \reg_array[1][5] ;
   wire \reg_array[1][4] ;
   wire \reg_array[1][3] ;
   wire \reg_array[1][2] ;
   wire \reg_array[1][1] ;
   wire \reg_array[1][0] ;
   wire \reg_array[0][15] ;
   wire \reg_array[0][14] ;
   wire \reg_array[0][13] ;
   wire \reg_array[0][12] ;
   wire \reg_array[0][11] ;
   wire \reg_array[0][10] ;
   wire \reg_array[0][9] ;
   wire \reg_array[0][8] ;
   wire \reg_array[0][7] ;
   wire \reg_array[0][6] ;
   wire \reg_array[0][5] ;
   wire \reg_array[0][4] ;
   wire \reg_array[0][3] ;
   wire \reg_array[0][2] ;
   wire \reg_array[0][1] ;
   wire \reg_array[0][0] ;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n238;
   wire n239;
   wire n240;

   assign N18 = reg_read_addr_1[0] ;
   assign N19 = reg_read_addr_1[1] ;
   assign N20 = reg_read_addr_1[2] ;
   assign N21 = reg_read_addr_2[0] ;
   assign N22 = reg_read_addr_2[1] ;
   assign N23 = reg_read_addr_2[2] ;

   BUFGHD FE_OFC95_n240 (.O(FE_OFN95_n240), 
	.I(n240));
   DFERBCHD \reg_array_reg[5][15]  (.RB(n240), 
	.Q(\reg_array[5][15] ), 
	.EB(n144), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[1][15]  (.RB(n240), 
	.Q(\reg_array[1][15] ), 
	.EB(n137), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[1][14]  (.RB(n240), 
	.Q(\reg_array[1][14] ), 
	.EB(n137), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[6][15]  (.RB(n240), 
	.Q(\reg_array[6][15] ), 
	.EB(n146), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[6][14]  (.RB(n240), 
	.Q(\reg_array[6][14] ), 
	.EB(n146), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[2][15]  (.RB(n240), 
	.Q(\reg_array[2][15] ), 
	.EB(n138), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[2][14]  (.RB(n240), 
	.Q(\reg_array[2][14] ), 
	.EB(n138), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[4][15]  (.RB(n240), 
	.Q(\reg_array[4][15] ), 
	.EB(n142), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[4][14]  (.RB(n240), 
	.Q(\reg_array[4][14] ), 
	.EB(n142), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[0][15]  (.RB(n240), 
	.Q(\reg_array[0][15] ), 
	.EB(n135), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[0][14]  (.RB(n240), 
	.Q(\reg_array[0][14] ), 
	.EB(n135), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[7][15]  (.RB(n240), 
	.Q(\reg_array[7][15] ), 
	.EB(n148), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[7][14]  (.RB(n240), 
	.Q(\reg_array[7][14] ), 
	.EB(n148), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[3][15]  (.RB(n240), 
	.Q(\reg_array[3][15] ), 
	.EB(n140), 
	.D(reg_write_data[15]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[3][14]  (.RB(n240), 
	.Q(\reg_array[3][14] ), 
	.EB(n140), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[5][14]  (.RB(n240), 
	.Q(\reg_array[5][14] ), 
	.EB(n144), 
	.D(reg_write_data[14]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[5][13]  (.RB(n240), 
	.Q(\reg_array[5][13] ), 
	.EB(n144), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[5][12]  (.RB(n240), 
	.Q(\reg_array[5][12] ), 
	.EB(n144), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[5][11]  (.RB(n240), 
	.Q(\reg_array[5][11] ), 
	.EB(n144), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[5][10]  (.RB(n240), 
	.Q(\reg_array[5][10] ), 
	.EB(n144), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[5][9]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][9] ), 
	.EB(n144), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[1][13]  (.RB(n240), 
	.Q(\reg_array[1][13] ), 
	.EB(n137), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[1][12]  (.RB(n240), 
	.Q(\reg_array[1][12] ), 
	.EB(n137), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[1][11]  (.RB(n240), 
	.Q(\reg_array[1][11] ), 
	.EB(n137), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[1][10]  (.RB(n240), 
	.Q(\reg_array[1][10] ), 
	.EB(n137), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[1][9]  (.RB(n240), 
	.Q(\reg_array[1][9] ), 
	.EB(n137), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[6][13]  (.RB(n240), 
	.Q(\reg_array[6][13] ), 
	.EB(n146), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[6][12]  (.RB(n240), 
	.Q(\reg_array[6][12] ), 
	.EB(n146), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[6][11]  (.RB(n240), 
	.Q(\reg_array[6][11] ), 
	.EB(n146), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[6][10]  (.RB(n240), 
	.Q(\reg_array[6][10] ), 
	.EB(n146), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[6][9]  (.RB(n240), 
	.Q(\reg_array[6][9] ), 
	.EB(n146), 
	.D(reg_write_data[9]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[2][13]  (.RB(n240), 
	.Q(\reg_array[2][13] ), 
	.EB(n138), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[2][12]  (.RB(n240), 
	.Q(\reg_array[2][12] ), 
	.EB(n138), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[2][11]  (.RB(n240), 
	.Q(\reg_array[2][11] ), 
	.EB(n138), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[2][10]  (.RB(n240), 
	.Q(\reg_array[2][10] ), 
	.EB(n138), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[2][9]  (.RB(n240), 
	.Q(\reg_array[2][9] ), 
	.EB(n138), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[4][13]  (.RB(n240), 
	.Q(\reg_array[4][13] ), 
	.EB(n142), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[4][12]  (.RB(n240), 
	.Q(\reg_array[4][12] ), 
	.EB(n142), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[4][11]  (.RB(n240), 
	.Q(\reg_array[4][11] ), 
	.EB(n142), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[4][10]  (.RB(n240), 
	.Q(\reg_array[4][10] ), 
	.EB(n142), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[4][9]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][9] ), 
	.EB(n142), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[0][13]  (.RB(n240), 
	.Q(\reg_array[0][13] ), 
	.EB(n135), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[0][12]  (.RB(n240), 
	.Q(\reg_array[0][12] ), 
	.EB(n135), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[0][11]  (.RB(n240), 
	.Q(\reg_array[0][11] ), 
	.EB(n135), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[0][10]  (.RB(n240), 
	.Q(\reg_array[0][10] ), 
	.EB(n135), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[0][9]  (.RB(n240), 
	.Q(\reg_array[0][9] ), 
	.EB(n135), 
	.D(reg_write_data[9]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[7][13]  (.RB(n240), 
	.Q(\reg_array[7][13] ), 
	.EB(n148), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[7][12]  (.RB(n240), 
	.Q(\reg_array[7][12] ), 
	.EB(n148), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[7][11]  (.RB(n240), 
	.Q(\reg_array[7][11] ), 
	.EB(n148), 
	.D(reg_write_data[11]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[7][10]  (.RB(n240), 
	.Q(\reg_array[7][10] ), 
	.EB(n148), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[7][9]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][9] ), 
	.EB(n148), 
	.D(reg_write_data[9]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[7][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][8] ), 
	.EB(n148), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[3][13]  (.RB(n240), 
	.Q(\reg_array[3][13] ), 
	.EB(n140), 
	.D(reg_write_data[13]), 
	.CK(clk_m__L3_N124));
   DFERBCHD \reg_array_reg[3][12]  (.RB(n240), 
	.Q(\reg_array[3][12] ), 
	.EB(n140), 
	.D(reg_write_data[12]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[3][11]  (.RB(n240), 
	.Q(\reg_array[3][11] ), 
	.EB(n140), 
	.D(reg_write_data[11]), 
	.CK(clk_m__L3_N123));
   DFERBCHD \reg_array_reg[3][10]  (.RB(n240), 
	.Q(\reg_array[3][10] ), 
	.EB(n140), 
	.D(reg_write_data[10]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[3][9]  (.RB(n240), 
	.Q(\reg_array[3][9] ), 
	.EB(n140), 
	.D(reg_write_data[9]), 
	.CK(clk));
   DFERBCHD \reg_array_reg[3][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][8] ), 
	.EB(n140), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[5][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][8] ), 
	.EB(n144), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[5][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][7] ), 
	.EB(n144), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[5][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][6] ), 
	.EB(n144), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[5][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][5] ), 
	.EB(n144), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[5][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][4] ), 
	.EB(n144), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[5][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][3] ), 
	.EB(n144), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[1][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][8] ), 
	.EB(n137), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[1][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][7] ), 
	.EB(n137), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[1][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][6] ), 
	.EB(n137), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[1][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][5] ), 
	.EB(n137), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[1][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][4] ), 
	.EB(n137), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[1][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][3] ), 
	.EB(n137), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[6][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][8] ), 
	.EB(n146), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[6][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][7] ), 
	.EB(n146), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[6][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][6] ), 
	.EB(n146), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[6][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][5] ), 
	.EB(n146), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[6][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][4] ), 
	.EB(n146), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[6][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][3] ), 
	.EB(n146), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[2][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][8] ), 
	.EB(n138), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[2][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][7] ), 
	.EB(n138), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[2][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][6] ), 
	.EB(n138), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[2][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][5] ), 
	.EB(n138), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[2][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][4] ), 
	.EB(n138), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[2][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][3] ), 
	.EB(n138), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[4][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][8] ), 
	.EB(n142), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[4][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][7] ), 
	.EB(n142), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[4][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][6] ), 
	.EB(n142), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[4][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][5] ), 
	.EB(n142), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[4][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][4] ), 
	.EB(n142), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[4][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][3] ), 
	.EB(n142), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][8]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][8] ), 
	.EB(n135), 
	.D(reg_write_data[8]), 
	.CK(clk_m__L3_N126));
   DFERBCHD \reg_array_reg[0][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][7] ), 
	.EB(n135), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[0][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][6] ), 
	.EB(n135), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N53));
   DFERBCHD \reg_array_reg[0][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][5] ), 
	.EB(n135), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[0][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][4] ), 
	.EB(n135), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][3] ), 
	.EB(n135), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[7][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][7] ), 
	.EB(n148), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[7][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][6] ), 
	.EB(n148), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N49));
   DFERBCHD \reg_array_reg[7][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][5] ), 
	.EB(n148), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[7][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][4] ), 
	.EB(n148), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[7][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][3] ), 
	.EB(n148), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[3][7]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][7] ), 
	.EB(n140), 
	.D(reg_write_data[7]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][6]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][6] ), 
	.EB(n140), 
	.D(reg_write_data[6]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][5]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][5] ), 
	.EB(n140), 
	.D(reg_write_data[5]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][4]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][4] ), 
	.EB(n140), 
	.D(reg_write_data[4]), 
	.CK(clk_m__L3_N50));
   DFERBCHD \reg_array_reg[3][3]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][3] ), 
	.EB(n140), 
	.D(reg_write_data[3]), 
	.CK(clk_m__L3_N54));
   DFERBCHD \reg_array_reg[5][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][2] ), 
	.EB(n144), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[5][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][1] ), 
	.EB(n144), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[5][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[5][0] ), 
	.EB(n144), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[1][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][2] ), 
	.EB(n137), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[1][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][1] ), 
	.EB(n137), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[1][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[1][0] ), 
	.EB(n137), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[6][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][2] ), 
	.EB(n146), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[6][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][1] ), 
	.EB(n146), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[6][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[6][0] ), 
	.EB(n146), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[2][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][2] ), 
	.EB(n138), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[2][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][1] ), 
	.EB(n138), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[2][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[2][0] ), 
	.EB(n138), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[4][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][2] ), 
	.EB(n142), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N80));
   DFERBCHD \reg_array_reg[4][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][1] ), 
	.EB(n142), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[4][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[4][0] ), 
	.EB(n142), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[0][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][2] ), 
	.EB(n135), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][1] ), 
	.EB(n135), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[0][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[0][0] ), 
	.EB(n135), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[7][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][2] ), 
	.EB(n148), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[7][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][1] ), 
	.EB(n148), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N80));
   DFERBCHD \reg_array_reg[7][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[7][0] ), 
	.EB(n148), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   DFERBCHD \reg_array_reg[3][2]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][2] ), 
	.EB(n140), 
	.D(reg_write_data[2]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[3][1]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][1] ), 
	.EB(n140), 
	.D(reg_write_data[1]), 
	.CK(clk_m__L3_N51));
   DFERBCHD \reg_array_reg[3][0]  (.RB(FE_OFN95_n240), 
	.Q(\reg_array[3][0] ), 
	.EB(n140), 
	.D(reg_write_data[0]), 
	.CK(clk_m__L3_N154));
   NR2CHD U2 (.O(n136), 
	.I2(reg_write_dest[1]), 
	.I1(reg_write_dest[2]));
   INVDHD U3 (.O(n239), 
	.I(reg_write_dest[0]));
   ND3CHD U17 (.O(n140), 
	.I3(n141), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[1]));
   NR2CHD U18 (.O(n141), 
	.I2(n238), 
	.I1(reg_write_dest[2]));
   ND3CHD U20 (.O(n144), 
	.I3(n145), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[2]));
   NR2CHD U21 (.O(n145), 
	.I2(n238), 
	.I1(reg_write_dest[1]));
   ND3CHD U23 (.O(n146), 
	.I3(n147), 
	.I2(reg_write_dest[1]), 
	.I1(reg_write_dest[2]));
   NR2CHD U24 (.O(n147), 
	.I2(n238), 
	.I1(reg_write_dest[0]));
   ND3CHD U26 (.O(n148), 
	.I3(n149), 
	.I2(reg_write_dest[1]), 
	.I1(reg_write_dest[2]));
   NR2CHD U27 (.O(n149), 
	.I2(n239), 
	.I1(n238));
   INVDHD U34 (.O(n238), 
	.I(reg_write_en));
   ND3CHD U36 (.O(n137), 
	.I3(n136), 
	.I2(reg_write_en), 
	.I1(reg_write_dest[0]));
   ND3CHD U38 (.O(n138), 
	.I3(n139), 
	.I2(reg_write_en), 
	.I1(reg_write_dest[1]));
   NR2CHD U39 (.O(n139), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[2]));
   ND3CHD U41 (.O(n142), 
	.I3(n143), 
	.I2(reg_write_en), 
	.I1(reg_write_dest[2]));
   NR2CHD U42 (.O(n143), 
	.I2(reg_write_dest[0]), 
	.I1(reg_write_dest[1]));
   ND3CHD U44 (.O(n135), 
	.I3(n136), 
	.I2(n239), 
	.I1(reg_write_en));
   AN2EHD U47 (.O(reg_read_data_1[1]), 
	.I2(n134), 
	.I1(N167));
   MUX2EHD U48 (.S(N20), 
	.O(N167), 
	.B(n131), 
	.A(n132));
   AN2EHD U49 (.O(reg_read_data_2[1]), 
	.I2(n133), 
	.I1(N183));
   MUX2EHD U50 (.S(N23), 
	.O(N183), 
	.B(n180), 
	.A(n181));
   AN2EHD U51 (.O(reg_read_data_2[2]), 
	.I2(n133), 
	.I1(N182));
   MUX2EHD U52 (.S(N23), 
	.O(N182), 
	.B(n182), 
	.A(n183));
   AN2EHD U53 (.O(reg_read_data_2[0]), 
	.I2(n133), 
	.I1(N184));
   MUX2EHD U54 (.S(N23), 
	.O(N184), 
	.B(n178), 
	.A(n179));
   AN2EHD U55 (.O(reg_read_data_1[0]), 
	.I2(n134), 
	.I1(N168));
   MUX2EHD U56 (.S(N20), 
	.O(N168), 
	.B(n129), 
	.A(n130));
   AN2EHD U57 (.O(reg_read_data_2[7]), 
	.I2(n133), 
	.I1(N177));
   MUX2EHD U58 (.S(N23), 
	.O(N177), 
	.B(n192), 
	.A(n193));
   AN2EHD U59 (.O(reg_read_data_2[8]), 
	.I2(n133), 
	.I1(N176));
   MUX2EHD U60 (.S(N23), 
	.O(N176), 
	.B(n194), 
	.A(n195));
   AN2EHD U61 (.O(reg_read_data_2[3]), 
	.I2(n133), 
	.I1(N181));
   MUX2EHD U62 (.S(N23), 
	.O(N181), 
	.B(n184), 
	.A(n185));
   AN2EHD U63 (.O(reg_read_data_2[4]), 
	.I2(n133), 
	.I1(N180));
   MUX2EHD U64 (.S(N23), 
	.O(N180), 
	.B(n186), 
	.A(n187));
   AN2EHD U65 (.O(reg_read_data_2[5]), 
	.I2(n133), 
	.I1(N179));
   MUX2EHD U66 (.S(N23), 
	.O(N179), 
	.B(n188), 
	.A(n189));
   AN2EHD U67 (.O(reg_read_data_2[6]), 
	.I2(n133), 
	.I1(N178));
   MUX2EHD U68 (.S(N23), 
	.O(N178), 
	.B(n190), 
	.A(n191));
   AN2EHD U69 (.O(reg_read_data_1[2]), 
	.I2(n134), 
	.I1(N166));
   MUX2EHD U70 (.S(N20), 
	.O(N166), 
	.B(n150), 
	.A(n151));
   AN2EHD U71 (.O(reg_read_data_1[3]), 
	.I2(n134), 
	.I1(N165));
   MUX2EHD U72 (.S(N20), 
	.O(N165), 
	.B(n152), 
	.A(n153));
   AN2EHD U73 (.O(reg_read_data_1[4]), 
	.I2(n134), 
	.I1(N164));
   MUX2EHD U74 (.S(N20), 
	.O(N164), 
	.B(n154), 
	.A(n155));
   AN2EHD U75 (.O(reg_read_data_1[5]), 
	.I2(n134), 
	.I1(N163));
   MUX2EHD U76 (.S(N20), 
	.O(N163), 
	.B(n156), 
	.A(n157));
   AN2EHD U77 (.O(reg_read_data_1[6]), 
	.I2(n134), 
	.I1(N162));
   MUX2EHD U78 (.S(N20), 
	.O(N162), 
	.B(n158), 
	.A(n159));
   AN2EHD U79 (.O(reg_read_data_1[7]), 
	.I2(n134), 
	.I1(N161));
   MUX2EHD U80 (.S(N20), 
	.O(N161), 
	.B(n160), 
	.A(n161));
   AN2EHD U81 (.O(reg_read_data_1[9]), 
	.I2(n134), 
	.I1(N159));
   MUX2EHD U82 (.S(N20), 
	.O(N159), 
	.B(n164), 
	.A(n165));
   AN2EHD U83 (.O(reg_read_data_1[13]), 
	.I2(n134), 
	.I1(N155));
   MUX2EHD U84 (.S(N20), 
	.O(N155), 
	.B(n172), 
	.A(n173));
   AN2EHD U85 (.O(reg_read_data_2[9]), 
	.I2(n133), 
	.I1(N175));
   MUX2EHD U86 (.S(N23), 
	.O(N175), 
	.B(n196), 
	.A(n197));
   AN2EHD U87 (.O(reg_read_data_2[10]), 
	.I2(n133), 
	.I1(N174));
   MUX2EHD U88 (.S(N23), 
	.O(N174), 
	.B(n198), 
	.A(n199));
   AN2EHD U89 (.O(reg_read_data_2[11]), 
	.I2(n133), 
	.I1(N173));
   MUX2EHD U90 (.S(N23), 
	.O(N173), 
	.B(n200), 
	.A(n201));
   AN2EHD U91 (.O(reg_read_data_2[12]), 
	.I2(n133), 
	.I1(N172));
   MUX2EHD U92 (.S(N23), 
	.O(N172), 
	.B(n202), 
	.A(n203));
   AN2EHD U93 (.O(reg_read_data_2[13]), 
	.I2(n133), 
	.I1(N171));
   MUX2EHD U94 (.S(N23), 
	.O(N171), 
	.B(n204), 
	.A(n205));
   AN2EHD U95 (.O(reg_read_data_2[14]), 
	.I2(n133), 
	.I1(N170));
   MUX2EHD U96 (.S(N23), 
	.O(N170), 
	.B(n206), 
	.A(n207));
   AN2EHD U97 (.O(reg_read_data_1[12]), 
	.I2(n134), 
	.I1(N156));
   MUX2EHD U98 (.S(N20), 
	.O(N156), 
	.B(n170), 
	.A(n171));
   AN2EHD U99 (.O(reg_read_data_1[8]), 
	.I2(n134), 
	.I1(N160));
   MUX2EHD U100 (.S(N20), 
	.O(N160), 
	.B(n162), 
	.A(n163));
   AN2EHD U101 (.O(reg_read_data_1[10]), 
	.I2(n134), 
	.I1(N158));
   MUX2EHD U102 (.S(N20), 
	.O(N158), 
	.B(n166), 
	.A(n167));
   AN2EHD U103 (.O(reg_read_data_1[11]), 
	.I2(n134), 
	.I1(N157));
   MUX2EHD U104 (.S(N20), 
	.O(N157), 
	.B(n168), 
	.A(n169));
   AN2EHD U105 (.O(reg_read_data_1[15]), 
	.I2(n134), 
	.I1(N153));
   MUX2EHD U106 (.S(N20), 
	.O(N153), 
	.B(n176), 
	.A(n177));
   AN2EHD U107 (.O(reg_read_data_2[15]), 
	.I2(n133), 
	.I1(N169));
   MUX2EHD U108 (.S(N23), 
	.O(N169), 
	.B(n208), 
	.A(n209));
   AN2EHD U109 (.O(reg_read_data_1[14]), 
	.I2(n134), 
	.I1(N154));
   MUX2EHD U110 (.S(N20), 
	.O(N154), 
	.B(n174), 
	.A(n175));
   INVDHD U111 (.O(n240), 
	.I(rst));
   OR3EHD U112 (.O(n133), 
	.I3(N21), 
	.I2(N23), 
	.I1(N22));
   OR3EHD U113 (.O(n134), 
	.I3(N18), 
	.I2(N20), 
	.I1(N19));
   MUX4EHD U114 (.S1(N18), 
	.S0(N19), 
	.O(n129), 
	.D(\reg_array[7][0] ), 
	.C(\reg_array[5][0] ), 
	.B(\reg_array[6][0] ), 
	.A(\reg_array[4][0] ));
   MUX4EHD U115 (.S1(N18), 
	.S0(N19), 
	.O(n130), 
	.D(\reg_array[3][0] ), 
	.C(\reg_array[1][0] ), 
	.B(\reg_array[2][0] ), 
	.A(\reg_array[0][0] ));
   MUX4EHD U116 (.S1(N18), 
	.S0(N19), 
	.O(n131), 
	.D(\reg_array[7][1] ), 
	.C(\reg_array[5][1] ), 
	.B(\reg_array[6][1] ), 
	.A(\reg_array[4][1] ));
   MUX4EHD U117 (.S1(N18), 
	.S0(N19), 
	.O(n132), 
	.D(\reg_array[3][1] ), 
	.C(\reg_array[1][1] ), 
	.B(\reg_array[2][1] ), 
	.A(\reg_array[0][1] ));
   MUX4EHD U118 (.S1(N18), 
	.S0(N19), 
	.O(n150), 
	.D(\reg_array[7][2] ), 
	.C(\reg_array[5][2] ), 
	.B(\reg_array[6][2] ), 
	.A(\reg_array[4][2] ));
   MUX4EHD U119 (.S1(N18), 
	.S0(N19), 
	.O(n151), 
	.D(\reg_array[3][2] ), 
	.C(\reg_array[1][2] ), 
	.B(\reg_array[2][2] ), 
	.A(\reg_array[0][2] ));
   MUX4EHD U120 (.S1(N18), 
	.S0(N19), 
	.O(n152), 
	.D(\reg_array[7][3] ), 
	.C(\reg_array[5][3] ), 
	.B(\reg_array[6][3] ), 
	.A(\reg_array[4][3] ));
   MUX4EHD U121 (.S1(N18), 
	.S0(N19), 
	.O(n153), 
	.D(\reg_array[3][3] ), 
	.C(\reg_array[1][3] ), 
	.B(\reg_array[2][3] ), 
	.A(\reg_array[0][3] ));
   MUX4EHD U122 (.S1(N18), 
	.S0(N19), 
	.O(n154), 
	.D(\reg_array[7][4] ), 
	.C(\reg_array[5][4] ), 
	.B(\reg_array[6][4] ), 
	.A(\reg_array[4][4] ));
   MUX4EHD U123 (.S1(N18), 
	.S0(N19), 
	.O(n155), 
	.D(\reg_array[3][4] ), 
	.C(\reg_array[1][4] ), 
	.B(\reg_array[2][4] ), 
	.A(\reg_array[0][4] ));
   MUX4EHD U124 (.S1(N18), 
	.S0(N19), 
	.O(n156), 
	.D(\reg_array[7][5] ), 
	.C(\reg_array[5][5] ), 
	.B(\reg_array[6][5] ), 
	.A(\reg_array[4][5] ));
   MUX4EHD U125 (.S1(N18), 
	.S0(N19), 
	.O(n157), 
	.D(\reg_array[3][5] ), 
	.C(\reg_array[1][5] ), 
	.B(\reg_array[2][5] ), 
	.A(\reg_array[0][5] ));
   MUX4EHD U126 (.S1(N18), 
	.S0(N19), 
	.O(n158), 
	.D(\reg_array[7][6] ), 
	.C(\reg_array[5][6] ), 
	.B(\reg_array[6][6] ), 
	.A(\reg_array[4][6] ));
   MUX4EHD U127 (.S1(N18), 
	.S0(N19), 
	.O(n159), 
	.D(\reg_array[3][6] ), 
	.C(\reg_array[1][6] ), 
	.B(\reg_array[2][6] ), 
	.A(\reg_array[0][6] ));
   MUX4EHD U128 (.S1(N18), 
	.S0(N19), 
	.O(n160), 
	.D(\reg_array[7][7] ), 
	.C(\reg_array[5][7] ), 
	.B(\reg_array[6][7] ), 
	.A(\reg_array[4][7] ));
   MUX4EHD U129 (.S1(N18), 
	.S0(N19), 
	.O(n161), 
	.D(\reg_array[3][7] ), 
	.C(\reg_array[1][7] ), 
	.B(\reg_array[2][7] ), 
	.A(\reg_array[0][7] ));
   MUX4EHD U130 (.S1(N18), 
	.S0(N19), 
	.O(n162), 
	.D(\reg_array[7][8] ), 
	.C(\reg_array[5][8] ), 
	.B(\reg_array[6][8] ), 
	.A(\reg_array[4][8] ));
   MUX4EHD U131 (.S1(N18), 
	.S0(N19), 
	.O(n163), 
	.D(\reg_array[3][8] ), 
	.C(\reg_array[1][8] ), 
	.B(\reg_array[2][8] ), 
	.A(\reg_array[0][8] ));
   MUX4EHD U132 (.S1(N18), 
	.S0(N19), 
	.O(n164), 
	.D(\reg_array[7][9] ), 
	.C(\reg_array[5][9] ), 
	.B(\reg_array[6][9] ), 
	.A(\reg_array[4][9] ));
   MUX4EHD U133 (.S1(N18), 
	.S0(N19), 
	.O(n165), 
	.D(\reg_array[3][9] ), 
	.C(\reg_array[1][9] ), 
	.B(\reg_array[2][9] ), 
	.A(\reg_array[0][9] ));
   MUX4EHD U134 (.S1(N18), 
	.S0(N19), 
	.O(n166), 
	.D(\reg_array[7][10] ), 
	.C(\reg_array[5][10] ), 
	.B(\reg_array[6][10] ), 
	.A(\reg_array[4][10] ));
   MUX4EHD U135 (.S1(N18), 
	.S0(N19), 
	.O(n167), 
	.D(\reg_array[3][10] ), 
	.C(\reg_array[1][10] ), 
	.B(\reg_array[2][10] ), 
	.A(\reg_array[0][10] ));
   MUX4EHD U136 (.S1(N18), 
	.S0(N19), 
	.O(n168), 
	.D(\reg_array[7][11] ), 
	.C(\reg_array[5][11] ), 
	.B(\reg_array[6][11] ), 
	.A(\reg_array[4][11] ));
   MUX4EHD U137 (.S1(N18), 
	.S0(N19), 
	.O(n169), 
	.D(\reg_array[3][11] ), 
	.C(\reg_array[1][11] ), 
	.B(\reg_array[2][11] ), 
	.A(\reg_array[0][11] ));
   MUX4EHD U138 (.S1(N18), 
	.S0(N19), 
	.O(n170), 
	.D(\reg_array[7][12] ), 
	.C(\reg_array[5][12] ), 
	.B(\reg_array[6][12] ), 
	.A(\reg_array[4][12] ));
   MUX4EHD U139 (.S1(N18), 
	.S0(N19), 
	.O(n171), 
	.D(\reg_array[3][12] ), 
	.C(\reg_array[1][12] ), 
	.B(\reg_array[2][12] ), 
	.A(\reg_array[0][12] ));
   MUX4EHD U140 (.S1(N18), 
	.S0(N19), 
	.O(n172), 
	.D(\reg_array[7][13] ), 
	.C(\reg_array[5][13] ), 
	.B(\reg_array[6][13] ), 
	.A(\reg_array[4][13] ));
   MUX4EHD U141 (.S1(N18), 
	.S0(N19), 
	.O(n173), 
	.D(\reg_array[3][13] ), 
	.C(\reg_array[1][13] ), 
	.B(\reg_array[2][13] ), 
	.A(\reg_array[0][13] ));
   MUX4EHD U142 (.S1(N18), 
	.S0(N19), 
	.O(n174), 
	.D(\reg_array[7][14] ), 
	.C(\reg_array[5][14] ), 
	.B(\reg_array[6][14] ), 
	.A(\reg_array[4][14] ));
   MUX4EHD U143 (.S1(N18), 
	.S0(N19), 
	.O(n175), 
	.D(\reg_array[3][14] ), 
	.C(\reg_array[1][14] ), 
	.B(\reg_array[2][14] ), 
	.A(\reg_array[0][14] ));
   MUX4EHD U144 (.S1(N18), 
	.S0(N19), 
	.O(n176), 
	.D(\reg_array[7][15] ), 
	.C(\reg_array[5][15] ), 
	.B(\reg_array[6][15] ), 
	.A(\reg_array[4][15] ));
   MUX4EHD U145 (.S1(N18), 
	.S0(N19), 
	.O(n177), 
	.D(\reg_array[3][15] ), 
	.C(\reg_array[1][15] ), 
	.B(\reg_array[2][15] ), 
	.A(\reg_array[0][15] ));
   MUX4EHD U146 (.S1(N21), 
	.S0(N22), 
	.O(n178), 
	.D(\reg_array[7][0] ), 
	.C(\reg_array[5][0] ), 
	.B(\reg_array[6][0] ), 
	.A(\reg_array[4][0] ));
   MUX4EHD U147 (.S1(N21), 
	.S0(N22), 
	.O(n179), 
	.D(\reg_array[3][0] ), 
	.C(\reg_array[1][0] ), 
	.B(\reg_array[2][0] ), 
	.A(\reg_array[0][0] ));
   MUX4EHD U148 (.S1(N21), 
	.S0(N22), 
	.O(n180), 
	.D(\reg_array[7][1] ), 
	.C(\reg_array[5][1] ), 
	.B(\reg_array[6][1] ), 
	.A(\reg_array[4][1] ));
   MUX4EHD U149 (.S1(N21), 
	.S0(N22), 
	.O(n181), 
	.D(\reg_array[3][1] ), 
	.C(\reg_array[1][1] ), 
	.B(\reg_array[2][1] ), 
	.A(\reg_array[0][1] ));
   MUX4EHD U150 (.S1(N21), 
	.S0(N22), 
	.O(n182), 
	.D(\reg_array[7][2] ), 
	.C(\reg_array[5][2] ), 
	.B(\reg_array[6][2] ), 
	.A(\reg_array[4][2] ));
   MUX4EHD U151 (.S1(N21), 
	.S0(N22), 
	.O(n183), 
	.D(\reg_array[3][2] ), 
	.C(\reg_array[1][2] ), 
	.B(\reg_array[2][2] ), 
	.A(\reg_array[0][2] ));
   MUX4EHD U152 (.S1(N21), 
	.S0(N22), 
	.O(n184), 
	.D(\reg_array[7][3] ), 
	.C(\reg_array[5][3] ), 
	.B(\reg_array[6][3] ), 
	.A(\reg_array[4][3] ));
   MUX4EHD U153 (.S1(N21), 
	.S0(N22), 
	.O(n185), 
	.D(\reg_array[3][3] ), 
	.C(\reg_array[1][3] ), 
	.B(\reg_array[2][3] ), 
	.A(\reg_array[0][3] ));
   MUX4EHD U154 (.S1(N21), 
	.S0(N22), 
	.O(n186), 
	.D(\reg_array[7][4] ), 
	.C(\reg_array[5][4] ), 
	.B(\reg_array[6][4] ), 
	.A(\reg_array[4][4] ));
   MUX4EHD U155 (.S1(N21), 
	.S0(N22), 
	.O(n187), 
	.D(\reg_array[3][4] ), 
	.C(\reg_array[1][4] ), 
	.B(\reg_array[2][4] ), 
	.A(\reg_array[0][4] ));
   MUX4EHD U156 (.S1(N21), 
	.S0(N22), 
	.O(n188), 
	.D(\reg_array[7][5] ), 
	.C(\reg_array[5][5] ), 
	.B(\reg_array[6][5] ), 
	.A(\reg_array[4][5] ));
   MUX4EHD U157 (.S1(N21), 
	.S0(N22), 
	.O(n189), 
	.D(\reg_array[3][5] ), 
	.C(\reg_array[1][5] ), 
	.B(\reg_array[2][5] ), 
	.A(\reg_array[0][5] ));
   MUX4EHD U158 (.S1(N21), 
	.S0(N22), 
	.O(n190), 
	.D(\reg_array[7][6] ), 
	.C(\reg_array[5][6] ), 
	.B(\reg_array[6][6] ), 
	.A(\reg_array[4][6] ));
   MUX4EHD U159 (.S1(N21), 
	.S0(N22), 
	.O(n191), 
	.D(\reg_array[3][6] ), 
	.C(\reg_array[1][6] ), 
	.B(\reg_array[2][6] ), 
	.A(\reg_array[0][6] ));
   MUX4EHD U160 (.S1(N21), 
	.S0(N22), 
	.O(n192), 
	.D(\reg_array[7][7] ), 
	.C(\reg_array[5][7] ), 
	.B(\reg_array[6][7] ), 
	.A(\reg_array[4][7] ));
   MUX4EHD U161 (.S1(N21), 
	.S0(N22), 
	.O(n193), 
	.D(\reg_array[3][7] ), 
	.C(\reg_array[1][7] ), 
	.B(\reg_array[2][7] ), 
	.A(\reg_array[0][7] ));
   MUX4EHD U162 (.S1(N21), 
	.S0(N22), 
	.O(n194), 
	.D(\reg_array[7][8] ), 
	.C(\reg_array[5][8] ), 
	.B(\reg_array[6][8] ), 
	.A(\reg_array[4][8] ));
   MUX4EHD U163 (.S1(N21), 
	.S0(N22), 
	.O(n195), 
	.D(\reg_array[3][8] ), 
	.C(\reg_array[1][8] ), 
	.B(\reg_array[2][8] ), 
	.A(\reg_array[0][8] ));
   MUX4EHD U164 (.S1(N21), 
	.S0(N22), 
	.O(n196), 
	.D(\reg_array[7][9] ), 
	.C(\reg_array[5][9] ), 
	.B(\reg_array[6][9] ), 
	.A(\reg_array[4][9] ));
   MUX4EHD U165 (.S1(N21), 
	.S0(N22), 
	.O(n197), 
	.D(\reg_array[3][9] ), 
	.C(\reg_array[1][9] ), 
	.B(\reg_array[2][9] ), 
	.A(\reg_array[0][9] ));
   MUX4EHD U166 (.S1(N21), 
	.S0(N22), 
	.O(n198), 
	.D(\reg_array[7][10] ), 
	.C(\reg_array[5][10] ), 
	.B(\reg_array[6][10] ), 
	.A(\reg_array[4][10] ));
   MUX4EHD U167 (.S1(N21), 
	.S0(N22), 
	.O(n199), 
	.D(\reg_array[3][10] ), 
	.C(\reg_array[1][10] ), 
	.B(\reg_array[2][10] ), 
	.A(\reg_array[0][10] ));
   MUX4EHD U168 (.S1(N21), 
	.S0(N22), 
	.O(n200), 
	.D(\reg_array[7][11] ), 
	.C(\reg_array[5][11] ), 
	.B(\reg_array[6][11] ), 
	.A(\reg_array[4][11] ));
   MUX4EHD U169 (.S1(N21), 
	.S0(N22), 
	.O(n201), 
	.D(\reg_array[3][11] ), 
	.C(\reg_array[1][11] ), 
	.B(\reg_array[2][11] ), 
	.A(\reg_array[0][11] ));
   MUX4EHD U170 (.S1(N21), 
	.S0(N22), 
	.O(n202), 
	.D(\reg_array[7][12] ), 
	.C(\reg_array[5][12] ), 
	.B(\reg_array[6][12] ), 
	.A(\reg_array[4][12] ));
   MUX4EHD U171 (.S1(N21), 
	.S0(N22), 
	.O(n203), 
	.D(\reg_array[3][12] ), 
	.C(\reg_array[1][12] ), 
	.B(\reg_array[2][12] ), 
	.A(\reg_array[0][12] ));
   MUX4EHD U172 (.S1(N21), 
	.S0(N22), 
	.O(n204), 
	.D(\reg_array[7][13] ), 
	.C(\reg_array[5][13] ), 
	.B(\reg_array[6][13] ), 
	.A(\reg_array[4][13] ));
   MUX4EHD U173 (.S1(N21), 
	.S0(N22), 
	.O(n205), 
	.D(\reg_array[3][13] ), 
	.C(\reg_array[1][13] ), 
	.B(\reg_array[2][13] ), 
	.A(\reg_array[0][13] ));
   MUX4EHD U174 (.S1(N21), 
	.S0(N22), 
	.O(n206), 
	.D(\reg_array[7][14] ), 
	.C(\reg_array[5][14] ), 
	.B(\reg_array[6][14] ), 
	.A(\reg_array[4][14] ));
   MUX4EHD U175 (.S1(N21), 
	.S0(N22), 
	.O(n207), 
	.D(\reg_array[3][14] ), 
	.C(\reg_array[1][14] ), 
	.B(\reg_array[2][14] ), 
	.A(\reg_array[0][14] ));
   MUX4EHD U176 (.S1(N21), 
	.S0(N22), 
	.O(n208), 
	.D(\reg_array[7][15] ), 
	.C(\reg_array[5][15] ), 
	.B(\reg_array[6][15] ), 
	.A(\reg_array[4][15] ));
   MUX4EHD U177 (.S1(N21), 
	.S0(N22), 
	.O(n209), 
	.D(\reg_array[3][15] ), 
	.C(\reg_array[1][15] ), 
	.B(\reg_array[2][15] ), 
	.A(\reg_array[0][15] ));
endmodule

module control (
	opcode, 
	reset, 
	reg_dst, 
	mem_to_reg, 
	alu_op, 
	jump, 
	branch, 
	mem_read, 
	mem_write, 
	alu_src, 
	reg_write, 
	sign_or_zero, 
	n75);
   input [2:0] opcode;
   input reset;
   output [1:0] reg_dst;
   output [1:0] mem_to_reg;
   output [1:0] alu_op;
   output jump;
   output branch;
   output mem_read;
   output mem_write;
   output alu_src;
   output reg_write;
   output sign_or_zero;
   input n75;

   // Internal wires
   wire \mem_to_reg[1] ;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n1;
   wire n2;
   wire n3;

   assign reg_dst[1] = \mem_to_reg[1]  ;
   assign mem_to_reg[1] = \mem_to_reg[1]  ;
   assign mem_to_reg[0] = mem_read ;
   assign alu_op[1] = alu_src ;

   AO12EHD U4 (.O(reg_write), 
	.B2(n75), 
	.B1(n7), 
	.A1(\mem_to_reg[1] ));
   OA13EHD U11 (.O(alu_src), 
	.B3(n13), 
	.B2(n9), 
	.B1(n12), 
	.A1(n75));
   ND2DHD U3 (.O(n12), 
	.I2(n8), 
	.I1(n14));
   OR3EHD U5 (.O(alu_op[0]), 
	.I3(branch), 
	.I2(mem_write), 
	.I1(mem_read));
   AN2HHD U6 (.O(mem_write), 
	.I2(n75), 
	.I1(n13));
   AN2EHD U7 (.O(reg_dst[0]), 
	.I2(n6), 
	.I1(n3));
   ND2DHD U8 (.O(sign_or_zero), 
	.I2(n6), 
	.I1(opcode[0]));
   NR2CHD U10 (.O(mem_read), 
	.I2(reset), 
	.I1(n14));
   AN2EHD U12 (.O(branch), 
	.I2(opcode[2]), 
	.I1(n11));
   NR2CHD U13 (.O(n11), 
	.I2(reset), 
	.I1(n2));
   OAI112BHD U14 (.O(n7), 
	.C2(opcode[0]), 
	.C1(opcode[1]), 
	.B1(n8), 
	.A1(n1));
   INVDHD U15 (.O(n1), 
	.I(n9));
   AN3EHD U16 (.O(\mem_to_reg[1] ), 
	.I3(n10), 
	.I2(opcode[1]), 
	.I1(opcode[0]));
   NR2CHD U17 (.O(n10), 
	.I2(opcode[2]), 
	.I1(reset));
   NR3BHD U18 (.O(n6), 
	.I3(opcode[1]), 
	.I2(reset), 
	.I1(opcode[2]));
   AN2B1CHD U19 (.O(jump), 
	.I1(n11), 
	.B1(opcode[2]));
   INVDHD U20 (.O(n2), 
	.I(opcode[1]));
   ND3CHD U21 (.O(n14), 
	.I3(opcode[2]), 
	.I2(n2), 
	.I1(n3));
   ND3CHD U22 (.O(n8), 
	.I3(opcode[0]), 
	.I2(opcode[2]), 
	.I1(opcode[1]));
   NR3BHD U23 (.O(n9), 
	.I3(n3), 
	.I2(opcode[2]), 
	.I1(opcode[1]));
   INVDHD U24 (.O(n3), 
	.I(opcode[0]));
   AN3EHD U25 (.O(n13), 
	.I3(opcode[0]), 
	.I2(n2), 
	.I1(opcode[2]));
endmodule

module instr_mem (
	pc, 
	instruction);
   input [15:0] pc;
   output [15:0] instruction;

   // Internal wires
   wire \instruction[0] ;

   assign instruction[15] = \instruction[0]  ;
   assign instruction[14] = \instruction[0]  ;
   assign instruction[13] = \instruction[0]  ;
   assign instruction[12] = \instruction[0]  ;
   assign instruction[11] = \instruction[0]  ;
   assign instruction[10] = \instruction[0]  ;
   assign instruction[9] = \instruction[0]  ;
   assign instruction[8] = \instruction[0]  ;
   assign instruction[7] = \instruction[0]  ;
   assign instruction[6] = \instruction[0]  ;
   assign instruction[5] = \instruction[0]  ;
   assign instruction[4] = \instruction[0]  ;
   assign instruction[3] = \instruction[0]  ;
   assign instruction[2] = \instruction[0]  ;
   assign instruction[1] = \instruction[0]  ;
   assign instruction[0] = \instruction[0]  ;

   TIE0DHD U2 (.O(\instruction[0] ));
endmodule

module mips_16 (
	clk, 
	reset, 
	pc_out, 
	alu_result, 
	clk_m__L3_N1, 
	clk_m__L3_N10, 
	clk_m__L3_N100, 
	clk_m__L3_N101, 
	clk_m__L3_N102, 
	clk_m__L3_N103, 
	clk_m__L3_N104, 
	clk_m__L3_N105, 
	clk_m__L3_N106, 
	clk_m__L3_N107, 
	clk_m__L3_N108, 
	clk_m__L3_N109, 
	clk_m__L3_N11, 
	clk_m__L3_N110, 
	clk_m__L3_N111, 
	clk_m__L3_N112, 
	clk_m__L3_N113, 
	clk_m__L3_N114, 
	clk_m__L3_N115, 
	clk_m__L3_N116, 
	clk_m__L3_N117, 
	clk_m__L3_N118, 
	clk_m__L3_N119, 
	clk_m__L3_N12, 
	clk_m__L3_N120, 
	clk_m__L3_N121, 
	clk_m__L3_N122, 
	clk_m__L3_N123, 
	clk_m__L3_N124, 
	clk_m__L3_N125, 
	clk_m__L3_N126, 
	clk_m__L3_N127, 
	clk_m__L3_N128, 
	clk_m__L3_N129, 
	clk_m__L3_N13, 
	clk_m__L3_N130, 
	clk_m__L3_N131, 
	clk_m__L3_N132, 
	clk_m__L3_N133, 
	clk_m__L3_N134, 
	clk_m__L3_N135, 
	clk_m__L3_N136, 
	clk_m__L3_N137, 
	clk_m__L3_N138, 
	clk_m__L3_N139, 
	clk_m__L3_N14, 
	clk_m__L3_N140, 
	clk_m__L3_N141, 
	clk_m__L3_N142, 
	clk_m__L3_N143, 
	clk_m__L3_N144, 
	clk_m__L3_N145, 
	clk_m__L3_N146, 
	clk_m__L3_N147, 
	clk_m__L3_N148, 
	clk_m__L3_N149, 
	clk_m__L3_N15, 
	clk_m__L3_N150, 
	clk_m__L3_N151, 
	clk_m__L3_N152, 
	clk_m__L3_N153, 
	clk_m__L3_N154, 
	clk_m__L3_N155, 
	clk_m__L3_N156, 
	clk_m__L3_N157, 
	clk_m__L3_N158, 
	clk_m__L3_N159, 
	clk_m__L3_N16, 
	clk_m__L3_N160, 
	clk_m__L3_N161, 
	clk_m__L3_N162, 
	clk_m__L3_N163, 
	clk_m__L3_N164, 
	clk_m__L3_N165, 
	clk_m__L3_N166, 
	clk_m__L3_N167, 
	clk_m__L3_N168, 
	clk_m__L3_N169, 
	clk_m__L3_N17, 
	clk_m__L3_N170, 
	clk_m__L3_N171, 
	clk_m__L3_N172, 
	clk_m__L3_N173, 
	clk_m__L3_N174, 
	clk_m__L3_N175, 
	clk_m__L3_N176, 
	clk_m__L3_N177, 
	clk_m__L3_N18, 
	clk_m__L3_N19, 
	clk_m__L3_N2, 
	clk_m__L3_N20, 
	clk_m__L3_N21, 
	clk_m__L3_N22, 
	clk_m__L3_N23, 
	clk_m__L3_N24, 
	clk_m__L3_N25, 
	clk_m__L3_N26, 
	clk_m__L3_N27, 
	clk_m__L3_N28, 
	clk_m__L3_N29, 
	clk_m__L3_N3, 
	clk_m__L3_N30, 
	clk_m__L3_N31, 
	clk_m__L3_N32, 
	clk_m__L3_N33, 
	clk_m__L3_N34, 
	clk_m__L3_N35, 
	clk_m__L3_N36, 
	clk_m__L3_N37, 
	clk_m__L3_N38, 
	clk_m__L3_N39, 
	clk_m__L3_N4, 
	clk_m__L3_N40, 
	clk_m__L3_N41, 
	clk_m__L3_N42, 
	clk_m__L3_N43, 
	clk_m__L3_N44, 
	clk_m__L3_N45, 
	clk_m__L3_N46, 
	clk_m__L3_N47, 
	clk_m__L3_N48, 
	clk_m__L3_N49, 
	clk_m__L3_N5, 
	clk_m__L3_N50, 
	clk_m__L3_N51, 
	clk_m__L3_N52, 
	clk_m__L3_N53, 
	clk_m__L3_N54, 
	clk_m__L3_N55, 
	clk_m__L3_N56, 
	clk_m__L3_N57, 
	clk_m__L3_N58, 
	clk_m__L3_N59, 
	clk_m__L3_N6, 
	clk_m__L3_N60, 
	clk_m__L3_N61, 
	clk_m__L3_N62, 
	clk_m__L3_N63, 
	clk_m__L3_N64, 
	clk_m__L3_N65, 
	clk_m__L3_N66, 
	clk_m__L3_N67, 
	clk_m__L3_N68, 
	clk_m__L3_N69, 
	clk_m__L3_N7, 
	clk_m__L3_N70, 
	clk_m__L3_N71, 
	clk_m__L3_N72, 
	clk_m__L3_N73, 
	clk_m__L3_N74, 
	clk_m__L3_N75, 
	clk_m__L3_N76, 
	clk_m__L3_N77, 
	clk_m__L3_N78, 
	clk_m__L3_N79, 
	clk_m__L3_N8, 
	clk_m__L3_N80, 
	clk_m__L3_N81, 
	clk_m__L3_N82, 
	clk_m__L3_N83, 
	clk_m__L3_N84, 
	clk_m__L3_N85, 
	clk_m__L3_N86, 
	clk_m__L3_N87, 
	clk_m__L3_N88, 
	clk_m__L3_N89, 
	clk_m__L3_N9, 
	clk_m__L3_N90, 
	clk_m__L3_N91, 
	clk_m__L3_N92, 
	clk_m__L3_N93, 
	clk_m__L3_N94, 
	clk_m__L3_N95, 
	clk_m__L3_N96, 
	clk_m__L3_N97, 
	clk_m__L3_N98, 
	clk_m__L3_N99, 
	clk_m__N0);
   input clk;
   input reset;
   output [15:0] pc_out;
   output [15:0] alu_result;
   input clk_m__L3_N1;
   input clk_m__L3_N10;
   input clk_m__L3_N100;
   input clk_m__L3_N101;
   input clk_m__L3_N102;
   input clk_m__L3_N103;
   input clk_m__L3_N104;
   input clk_m__L3_N105;
   input clk_m__L3_N106;
   input clk_m__L3_N107;
   input clk_m__L3_N108;
   input clk_m__L3_N109;
   input clk_m__L3_N11;
   input clk_m__L3_N110;
   input clk_m__L3_N111;
   input clk_m__L3_N112;
   input clk_m__L3_N113;
   input clk_m__L3_N114;
   input clk_m__L3_N115;
   input clk_m__L3_N116;
   input clk_m__L3_N117;
   input clk_m__L3_N118;
   input clk_m__L3_N119;
   input clk_m__L3_N12;
   input clk_m__L3_N120;
   input clk_m__L3_N121;
   input clk_m__L3_N122;
   input clk_m__L3_N123;
   input clk_m__L3_N124;
   input clk_m__L3_N125;
   input clk_m__L3_N126;
   input clk_m__L3_N127;
   input clk_m__L3_N128;
   input clk_m__L3_N129;
   input clk_m__L3_N13;
   input clk_m__L3_N130;
   input clk_m__L3_N131;
   input clk_m__L3_N132;
   input clk_m__L3_N133;
   input clk_m__L3_N134;
   input clk_m__L3_N135;
   input clk_m__L3_N136;
   input clk_m__L3_N137;
   input clk_m__L3_N138;
   input clk_m__L3_N139;
   input clk_m__L3_N14;
   input clk_m__L3_N140;
   input clk_m__L3_N141;
   input clk_m__L3_N142;
   input clk_m__L3_N143;
   input clk_m__L3_N144;
   input clk_m__L3_N145;
   input clk_m__L3_N146;
   input clk_m__L3_N147;
   input clk_m__L3_N148;
   input clk_m__L3_N149;
   input clk_m__L3_N15;
   input clk_m__L3_N150;
   input clk_m__L3_N151;
   input clk_m__L3_N152;
   input clk_m__L3_N153;
   input clk_m__L3_N154;
   input clk_m__L3_N155;
   input clk_m__L3_N156;
   input clk_m__L3_N157;
   input clk_m__L3_N158;
   input clk_m__L3_N159;
   input clk_m__L3_N16;
   input clk_m__L3_N160;
   input clk_m__L3_N161;
   input clk_m__L3_N162;
   input clk_m__L3_N163;
   input clk_m__L3_N164;
   input clk_m__L3_N165;
   input clk_m__L3_N166;
   input clk_m__L3_N167;
   input clk_m__L3_N168;
   input clk_m__L3_N169;
   input clk_m__L3_N17;
   input clk_m__L3_N170;
   input clk_m__L3_N171;
   input clk_m__L3_N172;
   input clk_m__L3_N173;
   input clk_m__L3_N174;
   input clk_m__L3_N175;
   input clk_m__L3_N176;
   input clk_m__L3_N177;
   input clk_m__L3_N18;
   input clk_m__L3_N19;
   input clk_m__L3_N2;
   input clk_m__L3_N20;
   input clk_m__L3_N21;
   input clk_m__L3_N22;
   input clk_m__L3_N23;
   input clk_m__L3_N24;
   input clk_m__L3_N25;
   input clk_m__L3_N26;
   input clk_m__L3_N27;
   input clk_m__L3_N28;
   input clk_m__L3_N29;
   input clk_m__L3_N3;
   input clk_m__L3_N30;
   input clk_m__L3_N31;
   input clk_m__L3_N32;
   input clk_m__L3_N33;
   input clk_m__L3_N34;
   input clk_m__L3_N35;
   input clk_m__L3_N36;
   input clk_m__L3_N37;
   input clk_m__L3_N38;
   input clk_m__L3_N39;
   input clk_m__L3_N4;
   input clk_m__L3_N40;
   input clk_m__L3_N41;
   input clk_m__L3_N42;
   input clk_m__L3_N43;
   input clk_m__L3_N44;
   input clk_m__L3_N45;
   input clk_m__L3_N46;
   input clk_m__L3_N47;
   input clk_m__L3_N48;
   input clk_m__L3_N49;
   input clk_m__L3_N5;
   input clk_m__L3_N50;
   input clk_m__L3_N51;
   input clk_m__L3_N52;
   input clk_m__L3_N53;
   input clk_m__L3_N54;
   input clk_m__L3_N55;
   input clk_m__L3_N56;
   input clk_m__L3_N57;
   input clk_m__L3_N58;
   input clk_m__L3_N59;
   input clk_m__L3_N6;
   input clk_m__L3_N60;
   input clk_m__L3_N61;
   input clk_m__L3_N62;
   input clk_m__L3_N63;
   input clk_m__L3_N64;
   input clk_m__L3_N65;
   input clk_m__L3_N66;
   input clk_m__L3_N67;
   input clk_m__L3_N68;
   input clk_m__L3_N69;
   input clk_m__L3_N7;
   input clk_m__L3_N70;
   input clk_m__L3_N71;
   input clk_m__L3_N72;
   input clk_m__L3_N73;
   input clk_m__L3_N74;
   input clk_m__L3_N75;
   input clk_m__L3_N76;
   input clk_m__L3_N77;
   input clk_m__L3_N78;
   input clk_m__L3_N79;
   input clk_m__L3_N8;
   input clk_m__L3_N80;
   input clk_m__L3_N81;
   input clk_m__L3_N82;
   input clk_m__L3_N83;
   input clk_m__L3_N84;
   input clk_m__L3_N85;
   input clk_m__L3_N86;
   input clk_m__L3_N87;
   input clk_m__L3_N88;
   input clk_m__L3_N89;
   input clk_m__L3_N9;
   input clk_m__L3_N90;
   input clk_m__L3_N91;
   input clk_m__L3_N92;
   input clk_m__L3_N93;
   input clk_m__L3_N94;
   input clk_m__L3_N95;
   input clk_m__L3_N96;
   input clk_m__L3_N97;
   input clk_m__L3_N98;
   input clk_m__L3_N99;
   input clk_m__N0;

   // Internal wires
   wire FE_PHN4010_pc_next_0_;
   wire FE_PHN3232_pc_next_0_;
   wire FE_PHN3231_pc_next_1_;
   wire FE_PHN99_pc_next_0_;
   wire FE_PHN98_pc_next_1_;
   wire FE_OFN97_n1;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire jump;
   wire branch;
   wire mem_read;
   wire mem_write;
   wire alu_src;
   wire reg_write;
   wire JRControl;
   wire zero_flag;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N67;
   wire N68;
   wire n31;
   wire n35;
   wire n36;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n69;
   wire \add_47/carry[15] ;
   wire \add_47/carry[14] ;
   wire \add_47/carry[13] ;
   wire \add_47/carry[12] ;
   wire \add_47/carry[11] ;
   wire \add_47/carry[10] ;
   wire \add_47/carry[9] ;
   wire \add_47/carry[8] ;
   wire \add_47/carry[7] ;
   wire \add_47/carry[6] ;
   wire \add_47/carry[5] ;
   wire \add_47/carry[4] ;
   wire \add_47/carry[3] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n32;
   wire n33;
   wire n34;
   wire n37;
   wire n68;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire [15:0] pc_next;
   wire [1:0] reg_dst;
   wire [1:0] mem_to_reg;
   wire [1:0] alu_op;
   wire [15:0] reg_write_data;
   wire [15:0] reg_read_data_1;
   wire [15:0] reg_read_data_2;
   wire [2:0] ALU_Control;
   wire [15:0] mem_read_data;

   assign pc_out[0] = N53 ;

   BUFCHD FE_PHC4010_pc_next_0_ (.O(FE_PHN4010_pc_next_0_), 
	.I(FE_PHN99_pc_next_0_));
   BUFCKEHD FE_PHC3232_pc_next_0_ (.O(FE_PHN3232_pc_next_0_), 
	.I(FE_PHN4010_pc_next_0_));
   BUFCHD FE_PHC3231_pc_next_1_ (.O(FE_PHN3231_pc_next_1_), 
	.I(pc_next[1]));
   BUFEHD FE_PHC99_pc_next_0_ (.O(FE_PHN99_pc_next_0_), 
	.I(pc_next[0]));
   BUFCHD FE_PHC98_pc_next_1_ (.O(FE_PHN98_pc_next_1_), 
	.I(FE_PHN3231_pc_next_1_));
   BUFKHD FE_OFC97_n1 (.O(n1), 
	.I(FE_OFN97_n1));
   AO222EHD U14 (.O(reg_write_data[9]), 
	.C2(n4), 
	.C1(N62), 
	.B2(n3), 
	.B1(alu_result[9]), 
	.A2(n31), 
	.A1(mem_read_data[9]));
   AO222EHD U15 (.O(reg_write_data[8]), 
	.C2(n4), 
	.C1(N61), 
	.B2(n3), 
	.B1(alu_result[8]), 
	.A2(n31), 
	.A1(mem_read_data[8]));
   AO222EHD U16 (.O(reg_write_data[7]), 
	.C2(n4), 
	.C1(N60), 
	.B2(n3), 
	.B1(alu_result[7]), 
	.A2(n31), 
	.A1(mem_read_data[7]));
   AO222EHD U17 (.O(reg_write_data[6]), 
	.C2(n4), 
	.C1(N59), 
	.B2(n3), 
	.B1(alu_result[6]), 
	.A2(n31), 
	.A1(mem_read_data[6]));
   AO222EHD U18 (.O(reg_write_data[5]), 
	.C2(n4), 
	.C1(N58), 
	.B2(n3), 
	.B1(alu_result[5]), 
	.A2(n31), 
	.A1(mem_read_data[5]));
   AO222EHD U19 (.O(reg_write_data[4]), 
	.C2(n4), 
	.C1(N57), 
	.B2(n3), 
	.B1(alu_result[4]), 
	.A2(n31), 
	.A1(mem_read_data[4]));
   AO222EHD U20 (.O(reg_write_data[3]), 
	.C2(n4), 
	.C1(N56), 
	.B2(n3), 
	.B1(alu_result[3]), 
	.A2(n31), 
	.A1(mem_read_data[3]));
   AO222EHD U21 (.O(reg_write_data[2]), 
	.C2(n4), 
	.C1(N55), 
	.B2(n3), 
	.B1(alu_result[2]), 
	.A2(n31), 
	.A1(mem_read_data[2]));
   AO222EHD U22 (.O(reg_write_data[1]), 
	.C2(n4), 
	.C1(N54), 
	.B2(n3), 
	.B1(alu_result[1]), 
	.A2(n31), 
	.A1(mem_read_data[1]));
   AO222EHD U23 (.O(reg_write_data[15]), 
	.C2(n4), 
	.C1(N68), 
	.B2(n3), 
	.B1(alu_result[15]), 
	.A2(n31), 
	.A1(mem_read_data[15]));
   AO222EHD U24 (.O(reg_write_data[14]), 
	.C2(n4), 
	.C1(N67), 
	.B2(n3), 
	.B1(alu_result[14]), 
	.A2(n31), 
	.A1(mem_read_data[14]));
   AO222EHD U25 (.O(reg_write_data[13]), 
	.C2(n4), 
	.C1(N66), 
	.B2(n3), 
	.B1(alu_result[13]), 
	.A2(n31), 
	.A1(mem_read_data[13]));
   AO222EHD U26 (.O(reg_write_data[12]), 
	.C2(n4), 
	.C1(N65), 
	.B2(n3), 
	.B1(alu_result[12]), 
	.A2(n31), 
	.A1(mem_read_data[12]));
   AO222EHD U27 (.O(reg_write_data[11]), 
	.C2(n4), 
	.C1(N64), 
	.B2(n3), 
	.B1(alu_result[11]), 
	.A2(n31), 
	.A1(mem_read_data[11]));
   AO222EHD U28 (.O(reg_write_data[10]), 
	.C2(n4), 
	.C1(N63), 
	.B2(n3), 
	.B1(alu_result[10]), 
	.A2(n31), 
	.A1(mem_read_data[10]));
   AO222EHD U29 (.O(reg_write_data[0]), 
	.C2(n4), 
	.C1(N53), 
	.B2(n3), 
	.B1(alu_result[0]), 
	.A2(n31), 
	.A1(mem_read_data[0]));
   OR2B1CHD U117 (.O(n57), 
	.I1(JRControl), 
	.B1(jump));
   instr_mem instrucion_memory (.pc({ pc_out[15],
		pc_out[14],
		pc_out[13],
		pc_out[12],
		pc_out[11],
		pc_out[10],
		pc_out[9],
		pc_out[8],
		pc_out[7],
		pc_out[6],
		pc_out[5],
		pc_out[4],
		pc_out[3],
		pc_out[2],
		pc_out[1],
		N53 }));
   control control_unit (.opcode({ n1,
		n1,
		n1 }), 
	.reset(reset), 
	.reg_dst({ reg_dst[1],
		reg_dst[0] }), 
	.mem_to_reg({ mem_to_reg[1],
		mem_to_reg[0] }), 
	.alu_op({ alu_op[1],
		alu_op[0] }), 
	.jump(jump), 
	.branch(branch), 
	.mem_read(mem_read), 
	.mem_write(mem_write), 
	.alu_src(alu_src), 
	.reg_write(reg_write), 
	.n75(n75));
   register_file reg_file (.clk(clk_m__L3_N122), 
	.rst(reset), 
	.reg_write_en(reg_write), 
	.reg_write_dest({ n2,
		n2,
		n2 }), 
	.reg_write_data({ reg_write_data[15],
		reg_write_data[14],
		reg_write_data[13],
		reg_write_data[12],
		reg_write_data[11],
		reg_write_data[10],
		reg_write_data[9],
		reg_write_data[8],
		reg_write_data[7],
		reg_write_data[6],
		reg_write_data[5],
		reg_write_data[4],
		reg_write_data[3],
		reg_write_data[2],
		reg_write_data[1],
		reg_write_data[0] }), 
	.reg_read_addr_1({ n1,
		n1,
		n1 }), 
	.reg_read_data_1({ reg_read_data_1[15],
		reg_read_data_1[14],
		reg_read_data_1[13],
		reg_read_data_1[12],
		reg_read_data_1[11],
		reg_read_data_1[10],
		reg_read_data_1[9],
		reg_read_data_1[8],
		reg_read_data_1[7],
		reg_read_data_1[6],
		reg_read_data_1[5],
		reg_read_data_1[4],
		reg_read_data_1[3],
		reg_read_data_1[2],
		reg_read_data_1[1],
		reg_read_data_1[0] }), 
	.reg_read_addr_2({ n1,
		n1,
		n1 }), 
	.reg_read_data_2({ reg_read_data_2[15],
		reg_read_data_2[14],
		reg_read_data_2[13],
		reg_read_data_2[12],
		reg_read_data_2[11],
		reg_read_data_2[10],
		reg_read_data_2[9],
		reg_read_data_2[8],
		reg_read_data_2[7],
		reg_read_data_2[6],
		reg_read_data_2[5],
		reg_read_data_2[4],
		reg_read_data_2[3],
		reg_read_data_2[2],
		reg_read_data_2[1],
		reg_read_data_2[0] }), 
	.clk_m__L3_N123(clk_m__L3_N123), 
	.clk_m__L3_N124(clk_m__L3_N124), 
	.clk_m__L3_N126(clk_m__L3_N126), 
	.clk_m__L3_N154(clk_m__L3_N154), 
	.clk_m__L3_N49(clk_m__L3_N49), 
	.clk_m__L3_N50(clk_m__L3_N50), 
	.clk_m__L3_N51(clk_m__L3_N51), 
	.clk_m__L3_N53(clk_m__L3_N53), 
	.clk_m__L3_N54(clk_m__L3_N54), 
	.clk_m__L3_N80(clk_m__L3_N80));
   JR_Control JRControl_unit (.alu_op({ alu_op[1],
		alu_op[0] }), 
	.funct({ n1,
		n1,
		n1,
		n1 }), 
	.JRControl(JRControl));
   ALUControl ALU_Control_unit (.ALU_Control({ ALU_Control[2],
		ALU_Control[1],
		ALU_Control[0] }), 
	.ALUOp({ alu_op[1],
		alu_op[0] }), 
	.Function({ n1,
		n1,
		n1,
		n1 }));
   alu alu_unit (.a({ reg_read_data_1[15],
		reg_read_data_1[14],
		reg_read_data_1[13],
		reg_read_data_1[12],
		reg_read_data_1[11],
		reg_read_data_1[10],
		reg_read_data_1[9],
		reg_read_data_1[8],
		reg_read_data_1[7],
		reg_read_data_1[6],
		reg_read_data_1[5],
		reg_read_data_1[4],
		reg_read_data_1[3],
		reg_read_data_1[2],
		reg_read_data_1[1],
		reg_read_data_1[0] }), 
	.b({ n16,
		n20,
		n18,
		n19,
		n17,
		n15,
		n14,
		n13,
		n12,
		n11,
		n7,
		n5,
		n6,
		n9,
		n8,
		n10 }), 
	.alu_control({ ALU_Control[2],
		ALU_Control[1],
		ALU_Control[0] }), 
	.result({ alu_result[15],
		alu_result[14],
		alu_result[13],
		alu_result[12],
		alu_result[11],
		alu_result[10],
		alu_result[9],
		alu_result[8],
		n76,
		n77,
		n78,
		n79,
		n80,
		n81,
		alu_result[1],
		alu_result[0] }), 
	.zero(zero_flag));
   data_memory datamem (.clk(clk), 
	.mem_access_addr({ alu_result[15],
		alu_result[14],
		alu_result[13],
		alu_result[12],
		alu_result[11],
		alu_result[10],
		alu_result[9],
		alu_result[8],
		alu_result[7],
		alu_result[6],
		alu_result[5],
		alu_result[4],
		alu_result[3],
		alu_result[2],
		alu_result[1],
		alu_result[0] }), 
	.mem_write_data({ reg_read_data_2[15],
		reg_read_data_2[14],
		reg_read_data_2[13],
		reg_read_data_2[12],
		reg_read_data_2[11],
		reg_read_data_2[10],
		reg_read_data_2[9],
		reg_read_data_2[8],
		reg_read_data_2[7],
		reg_read_data_2[6],
		reg_read_data_2[5],
		reg_read_data_2[4],
		reg_read_data_2[3],
		reg_read_data_2[2],
		reg_read_data_2[1],
		reg_read_data_2[0] }), 
	.mem_write_en(mem_write), 
	.mem_read(mem_read), 
	.mem_read_data({ mem_read_data[15],
		mem_read_data[14],
		mem_read_data[13],
		mem_read_data[12],
		mem_read_data[11],
		mem_read_data[10],
		mem_read_data[9],
		mem_read_data[8],
		mem_read_data[7],
		mem_read_data[6],
		mem_read_data[5],
		mem_read_data[4],
		mem_read_data[3],
		mem_read_data[2],
		mem_read_data[1],
		mem_read_data[0] }), 
	.clk_m__L3_N1(clk_m__L3_N1), 
	.clk_m__L3_N10(clk_m__L3_N10), 
	.clk_m__L3_N100(clk_m__L3_N100), 
	.clk_m__L3_N101(clk_m__L3_N101), 
	.clk_m__L3_N102(clk_m__L3_N102), 
	.clk_m__L3_N103(clk_m__L3_N103), 
	.clk_m__L3_N104(clk_m__L3_N104), 
	.clk_m__L3_N105(clk_m__L3_N105), 
	.clk_m__L3_N106(clk_m__L3_N106), 
	.clk_m__L3_N107(clk_m__L3_N107), 
	.clk_m__L3_N108(clk_m__L3_N108), 
	.clk_m__L3_N109(clk_m__L3_N109), 
	.clk_m__L3_N11(clk_m__L3_N11), 
	.clk_m__L3_N110(clk_m__L3_N110), 
	.clk_m__L3_N111(clk_m__L3_N111), 
	.clk_m__L3_N112(clk_m__L3_N112), 
	.clk_m__L3_N113(clk_m__L3_N113), 
	.clk_m__L3_N114(clk_m__L3_N114), 
	.clk_m__L3_N115(clk_m__L3_N115), 
	.clk_m__L3_N116(clk_m__L3_N116), 
	.clk_m__L3_N117(clk_m__L3_N117), 
	.clk_m__L3_N118(clk_m__L3_N118), 
	.clk_m__L3_N119(clk_m__L3_N119), 
	.clk_m__L3_N12(clk_m__L3_N12), 
	.clk_m__L3_N120(clk_m__L3_N120), 
	.clk_m__L3_N121(clk_m__L3_N121), 
	.clk_m__L3_N122(clk_m__L3_N122), 
	.clk_m__L3_N123(clk_m__L3_N123), 
	.clk_m__L3_N124(clk_m__L3_N124), 
	.clk_m__L3_N125(clk_m__L3_N125), 
	.clk_m__L3_N126(clk_m__L3_N126), 
	.clk_m__L3_N127(clk_m__L3_N127), 
	.clk_m__L3_N128(clk_m__L3_N128), 
	.clk_m__L3_N129(clk_m__L3_N129), 
	.clk_m__L3_N13(clk_m__L3_N13), 
	.clk_m__L3_N130(clk_m__L3_N130), 
	.clk_m__L3_N131(clk_m__L3_N131), 
	.clk_m__L3_N132(clk_m__L3_N132), 
	.clk_m__L3_N133(clk_m__L3_N133), 
	.clk_m__L3_N134(clk_m__L3_N134), 
	.clk_m__L3_N135(clk_m__L3_N135), 
	.clk_m__L3_N136(clk_m__L3_N136), 
	.clk_m__L3_N137(clk_m__L3_N137), 
	.clk_m__L3_N138(clk_m__L3_N138), 
	.clk_m__L3_N139(clk_m__L3_N139), 
	.clk_m__L3_N14(clk_m__L3_N14), 
	.clk_m__L3_N140(clk_m__L3_N140), 
	.clk_m__L3_N141(clk_m__L3_N141), 
	.clk_m__L3_N142(clk_m__L3_N142), 
	.clk_m__L3_N143(clk_m__L3_N143), 
	.clk_m__L3_N144(clk_m__L3_N144), 
	.clk_m__L3_N145(clk_m__L3_N145), 
	.clk_m__L3_N146(clk_m__L3_N146), 
	.clk_m__L3_N147(clk_m__L3_N147), 
	.clk_m__L3_N148(clk_m__L3_N148), 
	.clk_m__L3_N149(clk_m__L3_N149), 
	.clk_m__L3_N15(clk_m__L3_N15), 
	.clk_m__L3_N150(clk_m__L3_N150), 
	.clk_m__L3_N151(clk_m__L3_N151), 
	.clk_m__L3_N152(clk_m__L3_N152), 
	.clk_m__L3_N153(clk_m__L3_N153), 
	.clk_m__L3_N154(clk_m__L3_N154), 
	.clk_m__L3_N155(clk_m__L3_N155), 
	.clk_m__L3_N156(clk_m__L3_N156), 
	.clk_m__L3_N157(clk_m__L3_N157), 
	.clk_m__L3_N158(clk_m__L3_N158), 
	.clk_m__L3_N159(clk_m__L3_N159), 
	.clk_m__L3_N16(clk_m__L3_N16), 
	.clk_m__L3_N160(clk_m__L3_N160), 
	.clk_m__L3_N161(clk_m__L3_N161), 
	.clk_m__L3_N162(clk_m__L3_N162), 
	.clk_m__L3_N163(clk_m__L3_N163), 
	.clk_m__L3_N164(clk_m__L3_N164), 
	.clk_m__L3_N165(clk_m__L3_N165), 
	.clk_m__L3_N166(clk_m__L3_N166), 
	.clk_m__L3_N167(clk_m__L3_N167), 
	.clk_m__L3_N168(clk_m__L3_N168), 
	.clk_m__L3_N169(clk_m__L3_N169), 
	.clk_m__L3_N17(clk_m__L3_N17), 
	.clk_m__L3_N170(clk_m__L3_N170), 
	.clk_m__L3_N171(clk_m__L3_N171), 
	.clk_m__L3_N172(clk_m__L3_N172), 
	.clk_m__L3_N173(clk_m__L3_N173), 
	.clk_m__L3_N174(clk_m__L3_N174), 
	.clk_m__L3_N175(clk_m__L3_N175), 
	.clk_m__L3_N176(clk_m__L3_N176), 
	.clk_m__L3_N177(clk_m__L3_N177), 
	.clk_m__L3_N18(clk_m__L3_N18), 
	.clk_m__L3_N19(clk_m__L3_N19), 
	.clk_m__L3_N2(clk_m__L3_N2), 
	.clk_m__L3_N20(clk_m__L3_N20), 
	.clk_m__L3_N21(clk_m__L3_N21), 
	.clk_m__L3_N22(clk_m__L3_N22), 
	.clk_m__L3_N23(clk_m__L3_N23), 
	.clk_m__L3_N24(clk_m__L3_N24), 
	.clk_m__L3_N25(clk_m__L3_N25), 
	.clk_m__L3_N26(clk_m__L3_N26), 
	.clk_m__L3_N27(clk_m__L3_N27), 
	.clk_m__L3_N28(clk_m__L3_N28), 
	.clk_m__L3_N29(clk_m__L3_N29), 
	.clk_m__L3_N3(clk_m__L3_N3), 
	.clk_m__L3_N30(clk_m__L3_N30), 
	.clk_m__L3_N31(clk_m__L3_N31), 
	.clk_m__L3_N32(clk_m__L3_N32), 
	.clk_m__L3_N33(clk_m__L3_N33), 
	.clk_m__L3_N34(clk_m__L3_N34), 
	.clk_m__L3_N35(clk_m__L3_N35), 
	.clk_m__L3_N36(clk_m__L3_N36), 
	.clk_m__L3_N37(clk_m__L3_N37), 
	.clk_m__L3_N38(clk_m__L3_N38), 
	.clk_m__L3_N39(clk_m__L3_N39), 
	.clk_m__L3_N4(clk_m__L3_N4), 
	.clk_m__L3_N40(clk_m__L3_N40), 
	.clk_m__L3_N41(clk_m__L3_N41), 
	.clk_m__L3_N42(clk_m__L3_N42), 
	.clk_m__L3_N43(clk_m__L3_N43), 
	.clk_m__L3_N44(clk_m__L3_N44), 
	.clk_m__L3_N45(clk_m__L3_N45), 
	.clk_m__L3_N46(clk_m__L3_N46), 
	.clk_m__L3_N47(clk_m__L3_N47), 
	.clk_m__L3_N48(clk_m__L3_N48), 
	.clk_m__L3_N49(clk_m__L3_N49), 
	.clk_m__L3_N5(clk_m__L3_N5), 
	.clk_m__L3_N50(clk_m__L3_N50), 
	.clk_m__L3_N52(clk_m__L3_N52), 
	.clk_m__L3_N53(clk_m__L3_N53), 
	.clk_m__L3_N54(clk_m__L3_N54), 
	.clk_m__L3_N55(clk_m__L3_N55), 
	.clk_m__L3_N56(clk_m__L3_N56), 
	.clk_m__L3_N57(clk_m__L3_N57), 
	.clk_m__L3_N58(clk_m__L3_N58), 
	.clk_m__L3_N59(clk_m__L3_N59), 
	.clk_m__L3_N6(clk_m__L3_N6), 
	.clk_m__L3_N60(clk_m__L3_N60), 
	.clk_m__L3_N61(clk_m__L3_N61), 
	.clk_m__L3_N62(clk_m__L3_N62), 
	.clk_m__L3_N63(clk_m__L3_N63), 
	.clk_m__L3_N64(clk_m__L3_N64), 
	.clk_m__L3_N65(clk_m__L3_N65), 
	.clk_m__L3_N66(clk_m__L3_N66), 
	.clk_m__L3_N67(clk_m__L3_N67), 
	.clk_m__L3_N68(clk_m__L3_N68), 
	.clk_m__L3_N69(clk_m__L3_N69), 
	.clk_m__L3_N7(clk_m__L3_N7), 
	.clk_m__L3_N70(clk_m__L3_N70), 
	.clk_m__L3_N71(clk_m__L3_N71), 
	.clk_m__L3_N72(clk_m__L3_N72), 
	.clk_m__L3_N73(clk_m__L3_N73), 
	.clk_m__L3_N74(clk_m__L3_N74), 
	.clk_m__L3_N75(clk_m__L3_N75), 
	.clk_m__L3_N76(clk_m__L3_N76), 
	.clk_m__L3_N77(clk_m__L3_N77), 
	.clk_m__L3_N78(clk_m__L3_N78), 
	.clk_m__L3_N79(clk_m__L3_N79), 
	.clk_m__L3_N8(clk_m__L3_N8), 
	.clk_m__L3_N80(clk_m__L3_N80), 
	.clk_m__L3_N81(clk_m__L3_N81), 
	.clk_m__L3_N82(clk_m__L3_N82), 
	.clk_m__L3_N83(clk_m__L3_N83), 
	.clk_m__L3_N84(clk_m__L3_N84), 
	.clk_m__L3_N85(clk_m__L3_N85), 
	.clk_m__L3_N86(clk_m__L3_N86), 
	.clk_m__L3_N87(clk_m__L3_N87), 
	.clk_m__L3_N88(clk_m__L3_N88), 
	.clk_m__L3_N89(clk_m__L3_N89), 
	.clk_m__L3_N9(clk_m__L3_N9), 
	.clk_m__L3_N90(clk_m__L3_N90), 
	.clk_m__L3_N91(clk_m__L3_N91), 
	.clk_m__L3_N92(clk_m__L3_N92), 
	.clk_m__L3_N93(clk_m__L3_N93), 
	.clk_m__L3_N94(clk_m__L3_N94), 
	.clk_m__L3_N95(clk_m__L3_N95), 
	.clk_m__L3_N96(clk_m__L3_N96), 
	.clk_m__L3_N97(clk_m__L3_N97), 
	.clk_m__L3_N98(clk_m__L3_N98), 
	.clk_m__L3_N99(clk_m__L3_N99), 
	.clk_m__N0(clk_m__N0));
   QDFFRBEHD \pc_current_reg[15]  (.RB(n75), 
	.Q(pc_out[15]), 
	.D(pc_next[15]), 
	.CK(clk_m__L3_N124));
   QDFFRBEHD \pc_current_reg[9]  (.RB(n75), 
	.Q(pc_out[9]), 
	.D(pc_next[9]), 
	.CK(clk_m__L3_N126));
   QDFFRBEHD \pc_current_reg[8]  (.RB(n75), 
	.Q(pc_out[8]), 
	.D(pc_next[8]), 
	.CK(clk_m__L3_N126));
   QDFFRBEHD \pc_current_reg[7]  (.RB(n75), 
	.Q(pc_out[7]), 
	.D(pc_next[7]), 
	.CK(clk_m__L3_N50));
   QDFFRBEHD \pc_current_reg[6]  (.RB(n75), 
	.Q(pc_out[6]), 
	.D(pc_next[6]), 
	.CK(clk_m__L3_N50));
   QDFFRBEHD \pc_current_reg[5]  (.RB(n75), 
	.Q(pc_out[5]), 
	.D(pc_next[5]), 
	.CK(clk_m__L3_N50));
   QDFFRBEHD \pc_current_reg[4]  (.RB(n75), 
	.Q(pc_out[4]), 
	.D(pc_next[4]), 
	.CK(clk_m__L3_N51));
   QDFFRBEHD \pc_current_reg[3]  (.RB(n75), 
	.Q(pc_out[3]), 
	.D(pc_next[3]), 
	.CK(clk_m__L3_N51));
   QDFFRBEHD \pc_current_reg[2]  (.RB(n75), 
	.Q(pc_out[2]), 
	.D(pc_next[2]), 
	.CK(clk_m__L3_N154));
   QDFFRBEHD \pc_current_reg[14]  (.RB(n75), 
	.Q(pc_out[14]), 
	.D(pc_next[14]), 
	.CK(clk_m__L3_N124));
   QDFFRBEHD \pc_current_reg[13]  (.RB(n75), 
	.Q(pc_out[13]), 
	.D(pc_next[13]), 
	.CK(clk_m__L3_N123));
   QDFFRBEHD \pc_current_reg[12]  (.RB(n75), 
	.Q(pc_out[12]), 
	.D(pc_next[12]), 
	.CK(clk_m__L3_N123));
   QDFFRBEHD \pc_current_reg[11]  (.RB(n75), 
	.Q(pc_out[11]), 
	.D(pc_next[11]), 
	.CK(clk_m__L3_N122));
   QDFFRBEHD \pc_current_reg[10]  (.RB(n75), 
	.Q(pc_out[10]), 
	.D(pc_next[10]), 
	.CK(clk_m__L3_N122));
   QDFFRBEHD \pc_current_reg[1]  (.RB(n75), 
	.Q(pc_out[1]), 
	.D(FE_PHN98_pc_next_1_), 
	.CK(clk_m__L3_N51));
   QDFFRBEHD \pc_current_reg[0]  (.RB(n75), 
	.Q(N53), 
	.D(FE_PHN3232_pc_next_0_), 
	.CK(clk_m__L3_N154));
   TIE0KHD U3 (.O(FE_OFN97_n1));
   AN2EHD U4 (.O(n2), 
	.I2(n74), 
	.I1(reg_dst[1]));
   XNR2EHD U5 (.O(n3), 
	.I2(mem_to_reg[1]), 
	.I1(mem_to_reg[0]));
   AN2EHD U6 (.O(n4), 
	.I2(n72), 
	.I1(mem_to_reg[1]));
   INVDHD U7 (.O(n73), 
	.I(alu_src));
   BUFEHD U8 (.O(alu_result[6]), 
	.I(n77));
   BUFEHD U9 (.O(alu_result[7]), 
	.I(n76));
   BUFEHD U10 (.O(alu_result[4]), 
	.I(n79));
   BUFEHD U11 (.O(alu_result[2]), 
	.I(n81));
   BUFEHD U12 (.O(alu_result[5]), 
	.I(n78));
   BUFEHD U13 (.O(alu_result[3]), 
	.I(n80));
   INVDHD U30 (.O(n71), 
	.I(n69));
   AN2EHD U31 (.O(n5), 
	.I2(reg_read_data_2[4]), 
	.I1(n73));
   AN2EHD U32 (.O(n6), 
	.I2(reg_read_data_2[3]), 
	.I1(n73));
   AN2EHD U33 (.O(n7), 
	.I2(reg_read_data_2[5]), 
	.I1(n73));
   AN2EHD U34 (.O(n8), 
	.I2(reg_read_data_2[1]), 
	.I1(n73));
   AN2EHD U35 (.O(n9), 
	.I2(reg_read_data_2[2]), 
	.I1(n73));
   AN2EHD U36 (.O(n10), 
	.I2(reg_read_data_2[0]), 
	.I1(n73));
   AN2EHD U37 (.O(n11), 
	.I2(reg_read_data_2[6]), 
	.I1(n73));
   AN2EHD U38 (.O(n12), 
	.I2(n73), 
	.I1(reg_read_data_2[7]));
   AN2EHD U39 (.O(n13), 
	.I2(n73), 
	.I1(reg_read_data_2[8]));
   AN2EHD U40 (.O(n14), 
	.I2(n73), 
	.I1(reg_read_data_2[9]));
   AN2EHD U41 (.O(n15), 
	.I2(n73), 
	.I1(reg_read_data_2[10]));
   AN2EHD U42 (.O(n16), 
	.I2(n73), 
	.I1(reg_read_data_2[15]));
   AN2EHD U43 (.O(n17), 
	.I2(n73), 
	.I1(reg_read_data_2[11]));
   AN2EHD U44 (.O(n18), 
	.I2(n73), 
	.I1(reg_read_data_2[13]));
   AN2EHD U45 (.O(n19), 
	.I2(n73), 
	.I1(reg_read_data_2[12]));
   AN2EHD U46 (.O(n20), 
	.I2(n73), 
	.I1(reg_read_data_2[14]));
   NR3HHD U48 (.O(n38), 
	.I3(n69), 
	.I2(jump), 
	.I1(JRControl));
   ND3CHD U49 (.O(pc_next[15]), 
	.I3(n34), 
	.I2(n33), 
	.I1(n32));
   ND2DHD U50 (.O(n34), 
	.I2(JRControl), 
	.I1(reg_read_data_1[15]));
   ND2DHD U51 (.O(n33), 
	.I2(n56), 
	.I1(N68));
   ND2DHD U52 (.O(n32), 
	.I2(n38), 
	.I1(N68));
   OAI12CHD U53 (.O(n56), 
	.B2(n71), 
	.B1(JRControl), 
	.A1(n57));
   ND2DHD U54 (.O(n69), 
	.I2(branch), 
	.I1(zero_flag));
   NR3BHD U56 (.O(n39), 
	.I3(n71), 
	.I2(jump), 
	.I1(JRControl));
   ND2DHD U57 (.O(pc_next[10]), 
	.I2(n67), 
	.I1(n66));
   ND2DHD U58 (.O(n67), 
	.I2(n38), 
	.I1(N63));
   AOI22BHD U59 (.O(n66), 
	.B2(JRControl), 
	.B1(reg_read_data_1[10]), 
	.A2(N63), 
	.A1(n39));
   ND2DHD U60 (.O(pc_next[11]), 
	.I2(n65), 
	.I1(n64));
   ND2DHD U61 (.O(n65), 
	.I2(n38), 
	.I1(N64));
   AOI22BHD U62 (.O(n64), 
	.B2(JRControl), 
	.B1(reg_read_data_1[11]), 
	.A2(N64), 
	.A1(n39));
   ND2DHD U63 (.O(pc_next[12]), 
	.I2(n63), 
	.I1(n62));
   ND2DHD U64 (.O(n63), 
	.I2(n38), 
	.I1(N65));
   AOI22BHD U65 (.O(n62), 
	.B2(JRControl), 
	.B1(reg_read_data_1[12]), 
	.A2(N65), 
	.A1(n39));
   ND2DHD U66 (.O(pc_next[13]), 
	.I2(n61), 
	.I1(n60));
   ND2DHD U67 (.O(n61), 
	.I2(n38), 
	.I1(N66));
   AOI22BHD U68 (.O(n60), 
	.B2(JRControl), 
	.B1(reg_read_data_1[13]), 
	.A2(N66), 
	.A1(n39));
   ND2DHD U69 (.O(pc_next[14]), 
	.I2(n59), 
	.I1(n58));
   ND2DHD U70 (.O(n59), 
	.I2(n38), 
	.I1(N67));
   AOI22BHD U71 (.O(n58), 
	.B2(JRControl), 
	.B1(reg_read_data_1[14]), 
	.A2(N67), 
	.A1(n39));
   ND2DHD U72 (.O(pc_next[2]), 
	.I2(n53), 
	.I1(n52));
   ND2DHD U73 (.O(n53), 
	.I2(n38), 
	.I1(N55));
   AOI22BHD U74 (.O(n52), 
	.B2(JRControl), 
	.B1(reg_read_data_1[2]), 
	.A2(N55), 
	.A1(n39));
   ND2DHD U75 (.O(pc_next[3]), 
	.I2(n51), 
	.I1(n50));
   ND2DHD U76 (.O(n51), 
	.I2(n38), 
	.I1(N56));
   AOI22BHD U77 (.O(n50), 
	.B2(JRControl), 
	.B1(reg_read_data_1[3]), 
	.A2(N56), 
	.A1(n39));
   ND2DHD U78 (.O(pc_next[4]), 
	.I2(n49), 
	.I1(n48));
   ND2DHD U79 (.O(n49), 
	.I2(n38), 
	.I1(N57));
   AOI22BHD U80 (.O(n48), 
	.B2(JRControl), 
	.B1(reg_read_data_1[4]), 
	.A2(N57), 
	.A1(n39));
   ND2DHD U81 (.O(pc_next[5]), 
	.I2(n47), 
	.I1(n46));
   ND2DHD U82 (.O(n47), 
	.I2(n38), 
	.I1(N58));
   AOI22BHD U83 (.O(n46), 
	.B2(JRControl), 
	.B1(reg_read_data_1[5]), 
	.A2(N58), 
	.A1(n39));
   ND2DHD U84 (.O(pc_next[6]), 
	.I2(n45), 
	.I1(n44));
   ND2DHD U85 (.O(n45), 
	.I2(n38), 
	.I1(N59));
   AOI22BHD U86 (.O(n44), 
	.B2(JRControl), 
	.B1(reg_read_data_1[6]), 
	.A2(N59), 
	.A1(n39));
   ND2DHD U87 (.O(pc_next[7]), 
	.I2(n43), 
	.I1(n42));
   ND2DHD U88 (.O(n43), 
	.I2(n38), 
	.I1(N60));
   AOI22BHD U89 (.O(n42), 
	.B2(JRControl), 
	.B1(reg_read_data_1[7]), 
	.A2(N60), 
	.A1(n39));
   ND2DHD U90 (.O(pc_next[8]), 
	.I2(n41), 
	.I1(n40));
   ND2DHD U91 (.O(n41), 
	.I2(n38), 
	.I1(N61));
   AOI22BHD U92 (.O(n40), 
	.B2(JRControl), 
	.B1(reg_read_data_1[8]), 
	.A2(N61), 
	.A1(n39));
   ND2DHD U93 (.O(pc_next[9]), 
	.I2(n36), 
	.I1(n35));
   ND2DHD U94 (.O(n36), 
	.I2(n38), 
	.I1(N62));
   AOI22BHD U95 (.O(n35), 
	.B2(JRControl), 
	.B1(reg_read_data_1[9]), 
	.A2(N62), 
	.A1(n39));
   ND2DHD U96 (.O(pc_next[1]), 
	.I2(n55), 
	.I1(n54));
   ND2DHD U97 (.O(n55), 
	.I2(n38), 
	.I1(N54));
   AOI22BHD U98 (.O(n54), 
	.B2(JRControl), 
	.B1(reg_read_data_1[1]), 
	.A2(N54), 
	.A1(n39));
   NR2CHD U100 (.O(n31), 
	.I2(mem_to_reg[1]), 
	.I1(n72));
   INVDHD U101 (.O(n72), 
	.I(mem_to_reg[0]));
   INVDHD U102 (.O(n74), 
	.I(reg_dst[0]));
   ND3CHD U103 (.O(pc_next[0]), 
	.I3(n70), 
	.I2(n68), 
	.I1(n37));
   ND2DHD U104 (.O(n70), 
	.I2(JRControl), 
	.I1(reg_read_data_1[0]));
   ND2DHD U105 (.O(n37), 
	.I2(N53), 
	.I1(n39));
   ND2DHD U106 (.O(n68), 
	.I2(n38), 
	.I1(N53));
   INVDHD U108 (.O(N54), 
	.I(pc_out[1]));
   INVDHD U109 (.O(n75), 
	.I(reset));
   XOR2CHD U110 (.O(N68), 
	.I2(\add_47/carry[15] ), 
	.I1(pc_out[15]));
   AN2CHD U111 (.O(\add_47/carry[15] ), 
	.I2(\add_47/carry[14] ), 
	.I1(pc_out[14]));
   XOR2CHD U112 (.O(N67), 
	.I2(\add_47/carry[14] ), 
	.I1(pc_out[14]));
   AN2CHD U113 (.O(\add_47/carry[14] ), 
	.I2(\add_47/carry[13] ), 
	.I1(pc_out[13]));
   XOR2CHD U114 (.O(N66), 
	.I2(\add_47/carry[13] ), 
	.I1(pc_out[13]));
   AN2CHD U115 (.O(\add_47/carry[13] ), 
	.I2(\add_47/carry[12] ), 
	.I1(pc_out[12]));
   XOR2CHD U116 (.O(N65), 
	.I2(\add_47/carry[12] ), 
	.I1(pc_out[12]));
   AN2CHD U118 (.O(\add_47/carry[12] ), 
	.I2(\add_47/carry[11] ), 
	.I1(pc_out[11]));
   XOR2CHD U119 (.O(N64), 
	.I2(\add_47/carry[11] ), 
	.I1(pc_out[11]));
   AN2CHD U120 (.O(\add_47/carry[11] ), 
	.I2(\add_47/carry[10] ), 
	.I1(pc_out[10]));
   XOR2CHD U121 (.O(N63), 
	.I2(\add_47/carry[10] ), 
	.I1(pc_out[10]));
   AN2CHD U122 (.O(\add_47/carry[10] ), 
	.I2(\add_47/carry[9] ), 
	.I1(pc_out[9]));
   XOR2CHD U123 (.O(N62), 
	.I2(\add_47/carry[9] ), 
	.I1(pc_out[9]));
   AN2CHD U124 (.O(\add_47/carry[9] ), 
	.I2(\add_47/carry[8] ), 
	.I1(pc_out[8]));
   XOR2CHD U125 (.O(N61), 
	.I2(\add_47/carry[8] ), 
	.I1(pc_out[8]));
   AN2CHD U126 (.O(\add_47/carry[8] ), 
	.I2(\add_47/carry[7] ), 
	.I1(pc_out[7]));
   XOR2CHD U127 (.O(N60), 
	.I2(\add_47/carry[7] ), 
	.I1(pc_out[7]));
   AN2CHD U128 (.O(\add_47/carry[7] ), 
	.I2(\add_47/carry[6] ), 
	.I1(pc_out[6]));
   XOR2CHD U129 (.O(N59), 
	.I2(\add_47/carry[6] ), 
	.I1(pc_out[6]));
   AN2CHD U130 (.O(\add_47/carry[6] ), 
	.I2(\add_47/carry[5] ), 
	.I1(pc_out[5]));
   XOR2CHD U131 (.O(N58), 
	.I2(\add_47/carry[5] ), 
	.I1(pc_out[5]));
   AN2CHD U132 (.O(\add_47/carry[5] ), 
	.I2(\add_47/carry[4] ), 
	.I1(pc_out[4]));
   XOR2CHD U133 (.O(N57), 
	.I2(\add_47/carry[4] ), 
	.I1(pc_out[4]));
   AN2CHD U134 (.O(\add_47/carry[4] ), 
	.I2(\add_47/carry[3] ), 
	.I1(pc_out[3]));
   XOR2CHD U135 (.O(N56), 
	.I2(\add_47/carry[3] ), 
	.I1(pc_out[3]));
   AN2CHD U136 (.O(\add_47/carry[3] ), 
	.I2(pc_out[1]), 
	.I1(pc_out[2]));
   XOR2CHD U137 (.O(N55), 
	.I2(pc_out[1]), 
	.I1(pc_out[2]));
endmodule

module mips (
	vdd, 
	vddio, 
	gnd, 
	vss, 
	clk, 
	reset, 
	pc_out, 
	alu_result);
   inout vdd;
   inout vddio;
   inout gnd;
   inout vss;
   input clk;
   input reset;
   output [15:0] pc_out;
   output [15:0] alu_result;

   // Internal wires
   wire clk_m__N0;
   wire clk_m__L3_N177;
   wire clk_m__L3_N176;
   wire clk_m__L3_N175;
   wire clk_m__L3_N174;
   wire clk_m__L3_N173;
   wire clk_m__L3_N172;
   wire clk_m__L3_N171;
   wire clk_m__L3_N170;
   wire clk_m__L3_N169;
   wire clk_m__L3_N168;
   wire clk_m__L3_N167;
   wire clk_m__L3_N166;
   wire clk_m__L3_N165;
   wire clk_m__L3_N164;
   wire clk_m__L3_N163;
   wire clk_m__L3_N162;
   wire clk_m__L3_N161;
   wire clk_m__L3_N160;
   wire clk_m__L3_N159;
   wire clk_m__L3_N158;
   wire clk_m__L3_N157;
   wire clk_m__L3_N156;
   wire clk_m__L3_N155;
   wire clk_m__L3_N154;
   wire clk_m__L3_N153;
   wire clk_m__L3_N152;
   wire clk_m__L3_N151;
   wire clk_m__L3_N150;
   wire clk_m__L3_N149;
   wire clk_m__L3_N148;
   wire clk_m__L3_N147;
   wire clk_m__L3_N146;
   wire clk_m__L3_N145;
   wire clk_m__L3_N144;
   wire clk_m__L3_N143;
   wire clk_m__L3_N142;
   wire clk_m__L3_N141;
   wire clk_m__L3_N140;
   wire clk_m__L3_N139;
   wire clk_m__L3_N138;
   wire clk_m__L3_N137;
   wire clk_m__L3_N136;
   wire clk_m__L3_N135;
   wire clk_m__L3_N134;
   wire clk_m__L3_N133;
   wire clk_m__L3_N132;
   wire clk_m__L3_N131;
   wire clk_m__L3_N130;
   wire clk_m__L3_N129;
   wire clk_m__L3_N128;
   wire clk_m__L3_N127;
   wire clk_m__L3_N126;
   wire clk_m__L3_N125;
   wire clk_m__L3_N124;
   wire clk_m__L3_N123;
   wire clk_m__L3_N122;
   wire clk_m__L3_N121;
   wire clk_m__L3_N120;
   wire clk_m__L3_N119;
   wire clk_m__L3_N118;
   wire clk_m__L3_N117;
   wire clk_m__L3_N116;
   wire clk_m__L3_N115;
   wire clk_m__L3_N114;
   wire clk_m__L3_N113;
   wire clk_m__L3_N112;
   wire clk_m__L3_N111;
   wire clk_m__L3_N110;
   wire clk_m__L3_N109;
   wire clk_m__L3_N108;
   wire clk_m__L3_N107;
   wire clk_m__L3_N106;
   wire clk_m__L3_N105;
   wire clk_m__L3_N104;
   wire clk_m__L3_N103;
   wire clk_m__L3_N102;
   wire clk_m__L3_N101;
   wire clk_m__L3_N100;
   wire clk_m__L3_N99;
   wire clk_m__L3_N98;
   wire clk_m__L3_N97;
   wire clk_m__L3_N96;
   wire clk_m__L3_N95;
   wire clk_m__L3_N94;
   wire clk_m__L3_N93;
   wire clk_m__L3_N92;
   wire clk_m__L3_N91;
   wire clk_m__L3_N90;
   wire clk_m__L3_N89;
   wire clk_m__L3_N88;
   wire clk_m__L3_N87;
   wire clk_m__L3_N86;
   wire clk_m__L3_N85;
   wire clk_m__L3_N84;
   wire clk_m__L3_N83;
   wire clk_m__L3_N82;
   wire clk_m__L3_N81;
   wire clk_m__L3_N80;
   wire clk_m__L3_N79;
   wire clk_m__L3_N78;
   wire clk_m__L3_N77;
   wire clk_m__L3_N76;
   wire clk_m__L3_N75;
   wire clk_m__L3_N74;
   wire clk_m__L3_N73;
   wire clk_m__L3_N72;
   wire clk_m__L3_N71;
   wire clk_m__L3_N70;
   wire clk_m__L3_N69;
   wire clk_m__L3_N68;
   wire clk_m__L3_N67;
   wire clk_m__L3_N66;
   wire clk_m__L3_N65;
   wire clk_m__L3_N64;
   wire clk_m__L3_N63;
   wire clk_m__L3_N62;
   wire clk_m__L3_N61;
   wire clk_m__L3_N60;
   wire clk_m__L3_N59;
   wire clk_m__L3_N58;
   wire clk_m__L3_N57;
   wire clk_m__L3_N56;
   wire clk_m__L3_N55;
   wire clk_m__L3_N54;
   wire clk_m__L3_N53;
   wire clk_m__L3_N52;
   wire clk_m__L3_N51;
   wire clk_m__L3_N50;
   wire clk_m__L3_N49;
   wire clk_m__L3_N48;
   wire clk_m__L3_N47;
   wire clk_m__L3_N46;
   wire clk_m__L3_N45;
   wire clk_m__L3_N44;
   wire clk_m__L3_N43;
   wire clk_m__L3_N42;
   wire clk_m__L3_N41;
   wire clk_m__L3_N40;
   wire clk_m__L3_N39;
   wire clk_m__L3_N38;
   wire clk_m__L3_N37;
   wire clk_m__L3_N36;
   wire clk_m__L3_N35;
   wire clk_m__L3_N34;
   wire clk_m__L3_N33;
   wire clk_m__L3_N32;
   wire clk_m__L3_N31;
   wire clk_m__L3_N30;
   wire clk_m__L3_N29;
   wire clk_m__L3_N28;
   wire clk_m__L3_N27;
   wire clk_m__L3_N26;
   wire clk_m__L3_N25;
   wire clk_m__L3_N24;
   wire clk_m__L3_N23;
   wire clk_m__L3_N22;
   wire clk_m__L3_N21;
   wire clk_m__L3_N20;
   wire clk_m__L3_N19;
   wire clk_m__L3_N18;
   wire clk_m__L3_N17;
   wire clk_m__L3_N16;
   wire clk_m__L3_N15;
   wire clk_m__L3_N14;
   wire clk_m__L3_N13;
   wire clk_m__L3_N12;
   wire clk_m__L3_N11;
   wire clk_m__L3_N10;
   wire clk_m__L3_N9;
   wire clk_m__L3_N8;
   wire clk_m__L3_N7;
   wire clk_m__L3_N6;
   wire clk_m__L3_N5;
   wire clk_m__L3_N4;
   wire clk_m__L3_N3;
   wire clk_m__L3_N2;
   wire clk_m__L3_N1;
   wire clk_m__L3_N0;
   wire clk_m__L2_N17;
   wire clk_m__L2_N16;
   wire clk_m__L2_N15;
   wire clk_m__L2_N14;
   wire clk_m__L2_N13;
   wire clk_m__L2_N12;
   wire clk_m__L2_N11;
   wire clk_m__L2_N10;
   wire clk_m__L2_N9;
   wire clk_m__L2_N8;
   wire clk_m__L2_N7;
   wire clk_m__L2_N6;
   wire clk_m__L2_N5;
   wire clk_m__L2_N4;
   wire clk_m__L2_N3;
   wire clk_m__L2_N2;
   wire clk_m__L2_N1;
   wire clk_m__L2_N0;
   wire clk_m__L1_N5;
   wire clk_m__L1_N4;
   wire clk_m__L1_N3;
   wire clk_m__L1_N2;
   wire clk_m__L1_N1;
   wire clk_m__L1_N0;
   wire FE_OFN96_n1;
   wire clk_m;
   wire reset_m;
   wire n1;
   wire n2;
   wire [15:0] pc_out_m;
   wire [15:0] alu_result_m;

   BUFCKGHD clk_m__I0 (.O(clk_m__N0), 
	.I(clk_m__L2_N10));
   BUFCKGHD clk_m__L3_I177 (.O(clk_m__L3_N177), 
	.I(clk_m__L2_N17));
   BUFCKHHD clk_m__L3_I176 (.O(clk_m__L3_N176), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I175 (.O(clk_m__L3_N175), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I174 (.O(clk_m__L3_N174), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I173 (.O(clk_m__L3_N173), 
	.I(clk_m__L2_N17));
   BUFCKHHD clk_m__L3_I172 (.O(clk_m__L3_N172), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I171 (.O(clk_m__L3_N171), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I170 (.O(clk_m__L3_N170), 
	.I(clk_m__L2_N17));
   BUFCKHHD clk_m__L3_I169 (.O(clk_m__L3_N169), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I168 (.O(clk_m__L3_N168), 
	.I(clk_m__L2_N17));
   BUFCKGHD clk_m__L3_I167 (.O(clk_m__L3_N167), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I166 (.O(clk_m__L3_N166), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I165 (.O(clk_m__L3_N165), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I164 (.O(clk_m__L3_N164), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I163 (.O(clk_m__L3_N163), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I162 (.O(clk_m__L3_N162), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I161 (.O(clk_m__L3_N161), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I160 (.O(clk_m__L3_N160), 
	.I(clk_m__L2_N16));
   BUFCKHHD clk_m__L3_I159 (.O(clk_m__L3_N159), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I158 (.O(clk_m__L3_N158), 
	.I(clk_m__L2_N16));
   BUFCKGHD clk_m__L3_I157 (.O(clk_m__L3_N157), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I156 (.O(clk_m__L3_N156), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I155 (.O(clk_m__L3_N155), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I154 (.O(clk_m__L3_N154), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I153 (.O(clk_m__L3_N153), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I152 (.O(clk_m__L3_N152), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I151 (.O(clk_m__L3_N151), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I150 (.O(clk_m__L3_N150), 
	.I(clk_m__L2_N15));
   BUFCKHHD clk_m__L3_I149 (.O(clk_m__L3_N149), 
	.I(clk_m__L2_N15));
   BUFCKGHD clk_m__L3_I148 (.O(clk_m__L3_N148), 
	.I(clk_m__L2_N15));
   BUFCKHHD clk_m__L3_I147 (.O(clk_m__L3_N147), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I146 (.O(clk_m__L3_N146), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I145 (.O(clk_m__L3_N145), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I144 (.O(clk_m__L3_N144), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I143 (.O(clk_m__L3_N143), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I142 (.O(clk_m__L3_N142), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I141 (.O(clk_m__L3_N141), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I140 (.O(clk_m__L3_N140), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I139 (.O(clk_m__L3_N139), 
	.I(clk_m__L2_N14));
   BUFCKHHD clk_m__L3_I138 (.O(clk_m__L3_N138), 
	.I(clk_m__L2_N14));
   BUFCKGHD clk_m__L3_I137 (.O(clk_m__L3_N137), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I136 (.O(clk_m__L3_N136), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I135 (.O(clk_m__L3_N135), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I134 (.O(clk_m__L3_N134), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I133 (.O(clk_m__L3_N133), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I132 (.O(clk_m__L3_N132), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I131 (.O(clk_m__L3_N131), 
	.I(clk_m__L2_N13));
   BUFCKHHD clk_m__L3_I130 (.O(clk_m__L3_N130), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I129 (.O(clk_m__L3_N129), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I128 (.O(clk_m__L3_N128), 
	.I(clk_m__L2_N13));
   BUFCKGHD clk_m__L3_I127 (.O(clk_m__L3_N127), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I126 (.O(clk_m__L3_N126), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I125 (.O(clk_m__L3_N125), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I124 (.O(clk_m__L3_N124), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I123 (.O(clk_m__L3_N123), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I122 (.O(clk_m__L3_N122), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I121 (.O(clk_m__L3_N121), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I120 (.O(clk_m__L3_N120), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I119 (.O(clk_m__L3_N119), 
	.I(clk_m__L2_N12));
   BUFCKHHD clk_m__L3_I118 (.O(clk_m__L3_N118), 
	.I(clk_m__L2_N12));
   BUFCKGHD clk_m__L3_I117 (.O(clk_m__L3_N117), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I116 (.O(clk_m__L3_N116), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I115 (.O(clk_m__L3_N115), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I114 (.O(clk_m__L3_N114), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I113 (.O(clk_m__L3_N113), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I112 (.O(clk_m__L3_N112), 
	.I(clk_m__L2_N11));
   BUFCKGHD clk_m__L3_I111 (.O(clk_m__L3_N111), 
	.I(clk_m__L2_N11));
   BUFCKHHD clk_m__L3_I110 (.O(clk_m__L3_N110), 
	.I(clk_m__L2_N11));
   BUFCKHHD clk_m__L3_I109 (.O(clk_m__L3_N109), 
	.I(clk_m__L2_N11));
   BUFCKHHD clk_m__L3_I108 (.O(clk_m__L3_N108), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I107 (.O(clk_m__L3_N107), 
	.I(clk_m__L2_N10));
   BUFCKGHD clk_m__L3_I106 (.O(clk_m__L3_N106), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I105 (.O(clk_m__L3_N105), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I104 (.O(clk_m__L3_N104), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I103 (.O(clk_m__L3_N103), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I102 (.O(clk_m__L3_N102), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I101 (.O(clk_m__L3_N101), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I100 (.O(clk_m__L3_N100), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I99 (.O(clk_m__L3_N99), 
	.I(clk_m__L2_N10));
   BUFCKHHD clk_m__L3_I98 (.O(clk_m__L3_N98), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I97 (.O(clk_m__L3_N97), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I96 (.O(clk_m__L3_N96), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I95 (.O(clk_m__L3_N95), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I94 (.O(clk_m__L3_N94), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I93 (.O(clk_m__L3_N93), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I92 (.O(clk_m__L3_N92), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I91 (.O(clk_m__L3_N91), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I90 (.O(clk_m__L3_N90), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I89 (.O(clk_m__L3_N89), 
	.I(clk_m__L2_N9));
   BUFCKHHD clk_m__L3_I88 (.O(clk_m__L3_N88), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I87 (.O(clk_m__L3_N87), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I86 (.O(clk_m__L3_N86), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I85 (.O(clk_m__L3_N85), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I84 (.O(clk_m__L3_N84), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I83 (.O(clk_m__L3_N83), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I82 (.O(clk_m__L3_N82), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I81 (.O(clk_m__L3_N81), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I80 (.O(clk_m__L3_N80), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I79 (.O(clk_m__L3_N79), 
	.I(clk_m__L2_N8));
   BUFCKHHD clk_m__L3_I78 (.O(clk_m__L3_N78), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I77 (.O(clk_m__L3_N77), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I76 (.O(clk_m__L3_N76), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I75 (.O(clk_m__L3_N75), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I74 (.O(clk_m__L3_N74), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I73 (.O(clk_m__L3_N73), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I72 (.O(clk_m__L3_N72), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I71 (.O(clk_m__L3_N71), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I70 (.O(clk_m__L3_N70), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I69 (.O(clk_m__L3_N69), 
	.I(clk_m__L2_N7));
   BUFCKHHD clk_m__L3_I68 (.O(clk_m__L3_N68), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I67 (.O(clk_m__L3_N67), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I66 (.O(clk_m__L3_N66), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I65 (.O(clk_m__L3_N65), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I64 (.O(clk_m__L3_N64), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I63 (.O(clk_m__L3_N63), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I62 (.O(clk_m__L3_N62), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I61 (.O(clk_m__L3_N61), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I60 (.O(clk_m__L3_N60), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I59 (.O(clk_m__L3_N59), 
	.I(clk_m__L2_N6));
   BUFCKHHD clk_m__L3_I58 (.O(clk_m__L3_N58), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I57 (.O(clk_m__L3_N57), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I56 (.O(clk_m__L3_N56), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I55 (.O(clk_m__L3_N55), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I54 (.O(clk_m__L3_N54), 
	.I(clk_m__L2_N5));
   BUFCKHHD clk_m__L3_I53 (.O(clk_m__L3_N53), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I52 (.O(clk_m__L3_N52), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I51 (.O(clk_m__L3_N51), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I50 (.O(clk_m__L3_N50), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I49 (.O(clk_m__L3_N49), 
	.I(clk_m__L2_N5));
   BUFCKGHD clk_m__L3_I48 (.O(clk_m__L3_N48), 
	.I(clk_m__L2_N4));
   BUFCKGHD clk_m__L3_I47 (.O(clk_m__L3_N47), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I46 (.O(clk_m__L3_N46), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I45 (.O(clk_m__L3_N45), 
	.I(clk_m__L2_N4));
   BUFCKGHD clk_m__L3_I44 (.O(clk_m__L3_N44), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I43 (.O(clk_m__L3_N43), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I42 (.O(clk_m__L3_N42), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I41 (.O(clk_m__L3_N41), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I40 (.O(clk_m__L3_N40), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I39 (.O(clk_m__L3_N39), 
	.I(clk_m__L2_N4));
   BUFCKHHD clk_m__L3_I38 (.O(clk_m__L3_N38), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I37 (.O(clk_m__L3_N37), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I36 (.O(clk_m__L3_N36), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I35 (.O(clk_m__L3_N35), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I34 (.O(clk_m__L3_N34), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I33 (.O(clk_m__L3_N33), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I32 (.O(clk_m__L3_N32), 
	.I(clk_m__L2_N3));
   BUFCKGHD clk_m__L3_I31 (.O(clk_m__L3_N31), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I30 (.O(clk_m__L3_N30), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I29 (.O(clk_m__L3_N29), 
	.I(clk_m__L2_N3));
   BUFCKHHD clk_m__L3_I28 (.O(clk_m__L3_N28), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I27 (.O(clk_m__L3_N27), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I26 (.O(clk_m__L3_N26), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I25 (.O(clk_m__L3_N25), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I24 (.O(clk_m__L3_N24), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I23 (.O(clk_m__L3_N23), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I22 (.O(clk_m__L3_N22), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I21 (.O(clk_m__L3_N21), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I20 (.O(clk_m__L3_N20), 
	.I(clk_m__L2_N2));
   BUFCKHHD clk_m__L3_I19 (.O(clk_m__L3_N19), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I18 (.O(clk_m__L3_N18), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I17 (.O(clk_m__L3_N17), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I16 (.O(clk_m__L3_N16), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I15 (.O(clk_m__L3_N15), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I14 (.O(clk_m__L3_N14), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I13 (.O(clk_m__L3_N13), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I12 (.O(clk_m__L3_N12), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I11 (.O(clk_m__L3_N11), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I10 (.O(clk_m__L3_N10), 
	.I(clk_m__L2_N1));
   BUFCKHHD clk_m__L3_I9 (.O(clk_m__L3_N9), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I8 (.O(clk_m__L3_N8), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I7 (.O(clk_m__L3_N7), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I6 (.O(clk_m__L3_N6), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I5 (.O(clk_m__L3_N5), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I4 (.O(clk_m__L3_N4), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I3 (.O(clk_m__L3_N3), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I2 (.O(clk_m__L3_N2), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I1 (.O(clk_m__L3_N1), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L3_I0 (.O(clk_m__L3_N0), 
	.I(clk_m__L2_N0));
   BUFCKHHD clk_m__L2_I17 (.O(clk_m__L2_N17), 
	.I(clk_m__L1_N5));
   BUFCKHHD clk_m__L2_I16 (.O(clk_m__L2_N16), 
	.I(clk_m__L1_N5));
   BUFCKHHD clk_m__L2_I15 (.O(clk_m__L2_N15), 
	.I(clk_m__L1_N5));
   BUFCKHHD clk_m__L2_I14 (.O(clk_m__L2_N14), 
	.I(clk_m__L1_N4));
   BUFCKHHD clk_m__L2_I13 (.O(clk_m__L2_N13), 
	.I(clk_m__L1_N4));
   BUFCKHHD clk_m__L2_I12 (.O(clk_m__L2_N12), 
	.I(clk_m__L1_N4));
   BUFCKHHD clk_m__L2_I11 (.O(clk_m__L2_N11), 
	.I(clk_m__L1_N3));
   BUFCKHHD clk_m__L2_I10 (.O(clk_m__L2_N10), 
	.I(clk_m__L1_N3));
   BUFCKHHD clk_m__L2_I9 (.O(clk_m__L2_N9), 
	.I(clk_m__L1_N3));
   BUFCKHHD clk_m__L2_I8 (.O(clk_m__L2_N8), 
	.I(clk_m__L1_N2));
   BUFCKHHD clk_m__L2_I7 (.O(clk_m__L2_N7), 
	.I(clk_m__L1_N2));
   BUFCKHHD clk_m__L2_I6 (.O(clk_m__L2_N6), 
	.I(clk_m__L1_N2));
   BUFCKHHD clk_m__L2_I5 (.O(clk_m__L2_N5), 
	.I(clk_m__L1_N1));
   BUFCKHHD clk_m__L2_I4 (.O(clk_m__L2_N4), 
	.I(clk_m__L1_N1));
   BUFCKHHD clk_m__L2_I3 (.O(clk_m__L2_N3), 
	.I(clk_m__L1_N1));
   BUFCKHHD clk_m__L2_I2 (.O(clk_m__L2_N2), 
	.I(clk_m__L1_N0));
   BUFCKHHD clk_m__L2_I1 (.O(clk_m__L2_N1), 
	.I(clk_m__L1_N0));
   BUFCKHHD clk_m__L2_I0 (.O(clk_m__L2_N0), 
	.I(clk_m__L1_N0));
   BUFCKHHD clk_m__L1_I5 (.O(clk_m__L1_N5), 
	.I(clk_m));
   BUFCKGHD clk_m__L1_I4 (.O(clk_m__L1_N4), 
	.I(clk_m));
   BUFCKHHD clk_m__L1_I3 (.O(clk_m__L1_N3), 
	.I(clk_m));
   BUFCKHHD clk_m__L1_I2 (.O(clk_m__L1_N2), 
	.I(clk_m));
   BUFCKGHD clk_m__L1_I1 (.O(clk_m__L1_N1), 
	.I(clk_m));
   BUFCKHHD clk_m__L1_I0 (.O(clk_m__L1_N0), 
	.I(clk_m));
   BUFCKIHD FE_OFC96_n1 (.O(FE_OFN96_n1), 
	.I(n1));
   XMHA in1 (.SMT(n1), 
	.PU(n1), 
	.PD(n1), 
	.O(clk_m), 
	.I(clk));
   XMHA in2 (.SMT(n1), 
	.PU(n1), 
	.PD(n1), 
	.O(reset_m), 
	.I(reset));
   YA28SHA out1 (.SR(n1), 
	.O(pc_out[0]), 
	.I(pc_out_m[0]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out2 (.SR(n1), 
	.O(pc_out[1]), 
	.I(pc_out_m[1]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out3 (.SR(n1), 
	.O(pc_out[2]), 
	.I(pc_out_m[2]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out4 (.SR(n1), 
	.O(pc_out[3]), 
	.I(pc_out_m[3]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out5 (.SR(n1), 
	.O(pc_out[4]), 
	.I(pc_out_m[4]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out6 (.SR(FE_OFN96_n1), 
	.O(pc_out[5]), 
	.I(pc_out_m[5]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out7 (.SR(FE_OFN96_n1), 
	.O(pc_out[6]), 
	.I(pc_out_m[6]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out8 (.SR(n1), 
	.O(pc_out[7]), 
	.I(pc_out_m[7]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out9 (.SR(n1), 
	.O(pc_out[8]), 
	.I(pc_out_m[8]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out10 (.SR(n1), 
	.O(pc_out[9]), 
	.I(pc_out_m[9]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out11 (.SR(n1), 
	.O(pc_out[10]), 
	.I(pc_out_m[10]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out12 (.SR(n1), 
	.O(pc_out[11]), 
	.I(pc_out_m[11]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out13 (.SR(n1), 
	.O(pc_out[12]), 
	.I(pc_out_m[12]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out14 (.SR(n1), 
	.O(pc_out[13]), 
	.I(pc_out_m[13]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out15 (.SR(n1), 
	.O(pc_out[14]), 
	.I(pc_out_m[14]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out16 (.SR(n1), 
	.O(pc_out[15]), 
	.I(pc_out_m[15]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out17 (.SR(n1), 
	.O(alu_result[0]), 
	.I(alu_result_m[0]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out18 (.SR(n1), 
	.O(alu_result[1]), 
	.I(alu_result_m[1]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out19 (.SR(n1), 
	.O(alu_result[2]), 
	.I(alu_result_m[2]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out20 (.SR(n1), 
	.O(alu_result[3]), 
	.I(alu_result_m[3]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out21 (.SR(n1), 
	.O(alu_result[4]), 
	.I(alu_result_m[4]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out22 (.SR(n1), 
	.O(alu_result[5]), 
	.I(alu_result_m[5]), 
	.E4(n1), 
	.E2(n1), 
	.E(n2));
   YA28SHA out23 (.SR(FE_OFN96_n1), 
	.O(alu_result[6]), 
	.I(alu_result_m[6]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out24 (.SR(FE_OFN96_n1), 
	.O(alu_result[7]), 
	.I(alu_result_m[7]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out25 (.SR(FE_OFN96_n1), 
	.O(alu_result[8]), 
	.I(alu_result_m[8]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out26 (.SR(FE_OFN96_n1), 
	.O(alu_result[9]), 
	.I(alu_result_m[9]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out27 (.SR(FE_OFN96_n1), 
	.O(alu_result[10]), 
	.I(alu_result_m[10]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out28 (.SR(FE_OFN96_n1), 
	.O(alu_result[11]), 
	.I(alu_result_m[11]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out29 (.SR(FE_OFN96_n1), 
	.O(alu_result[12]), 
	.I(alu_result_m[12]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out30 (.SR(FE_OFN96_n1), 
	.O(alu_result[13]), 
	.I(alu_result_m[13]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out31 (.SR(FE_OFN96_n1), 
	.O(alu_result[14]), 
	.I(alu_result_m[14]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   YA28SHA out32 (.SR(FE_OFN96_n1), 
	.O(alu_result[15]), 
	.I(alu_result_m[15]), 
	.E4(FE_OFN96_n1), 
	.E2(FE_OFN96_n1), 
	.E(n2));
   VCCKHA pwr_1 (.VCC(vdd));
   VCCKHA pwr_2 (.VCC(vdd));
   VCCKHA pwr_3 (.VCC(vdd));
   VCCKHA pwr_4 (.VCC(vdd));
   VCC3IHA pwr_5 (.VCC3I(vddio));
   VCC3IHA pwr_6 (.VCC3I(vddio));
   VCC3IHA pwr_7 (.VCC3I(vddio));
   VCC3IHA pwr_8 (.VCC3I(vddio));
   GND3IHA gnd_1 (.GND3I(vss));
   GND3IHA gnd_2 (.GND3I(vss));
   GND3IHA gnd_3 (.GND3I(vss));
   GND3IHA gnd_4 (.GND3I(vss));
   GNDKHA gnd_5 (.GND(gnd));
   GNDKHA gnd_6 (.GND(gnd));
   GNDKHA gnd_7 (.GND(gnd));
   GNDKHA gnd_8 (.GND(gnd));
   CORNERHA corner_1 ();
   CORNERHA corner_2 ();
   CORNERHA corner_3 ();
   CORNERHA corner_4 ();
   mips_16 mips_core (.clk(clk_m__L3_N0), 
	.reset(reset_m), 
	.pc_out({ pc_out_m[15],
		pc_out_m[14],
		pc_out_m[13],
		pc_out_m[12],
		pc_out_m[11],
		pc_out_m[10],
		pc_out_m[9],
		pc_out_m[8],
		pc_out_m[7],
		pc_out_m[6],
		pc_out_m[5],
		pc_out_m[4],
		pc_out_m[3],
		pc_out_m[2],
		pc_out_m[1],
		pc_out_m[0] }), 
	.alu_result({ alu_result_m[15],
		alu_result_m[14],
		alu_result_m[13],
		alu_result_m[12],
		alu_result_m[11],
		alu_result_m[10],
		alu_result_m[9],
		alu_result_m[8],
		alu_result_m[7],
		alu_result_m[6],
		alu_result_m[5],
		alu_result_m[4],
		alu_result_m[3],
		alu_result_m[2],
		alu_result_m[1],
		alu_result_m[0] }), 
	.clk_m__L3_N1(clk_m__L3_N1), 
	.clk_m__L3_N10(clk_m__L3_N10), 
	.clk_m__L3_N100(clk_m__L3_N100), 
	.clk_m__L3_N101(clk_m__L3_N101), 
	.clk_m__L3_N102(clk_m__L3_N102), 
	.clk_m__L3_N103(clk_m__L3_N103), 
	.clk_m__L3_N104(clk_m__L3_N104), 
	.clk_m__L3_N105(clk_m__L3_N105), 
	.clk_m__L3_N106(clk_m__L3_N106), 
	.clk_m__L3_N107(clk_m__L3_N107), 
	.clk_m__L3_N108(clk_m__L3_N108), 
	.clk_m__L3_N109(clk_m__L3_N109), 
	.clk_m__L3_N11(clk_m__L3_N11), 
	.clk_m__L3_N110(clk_m__L3_N110), 
	.clk_m__L3_N111(clk_m__L3_N111), 
	.clk_m__L3_N112(clk_m__L3_N112), 
	.clk_m__L3_N113(clk_m__L3_N113), 
	.clk_m__L3_N114(clk_m__L3_N114), 
	.clk_m__L3_N115(clk_m__L3_N115), 
	.clk_m__L3_N116(clk_m__L3_N116), 
	.clk_m__L3_N117(clk_m__L3_N117), 
	.clk_m__L3_N118(clk_m__L3_N118), 
	.clk_m__L3_N119(clk_m__L3_N119), 
	.clk_m__L3_N12(clk_m__L3_N12), 
	.clk_m__L3_N120(clk_m__L3_N120), 
	.clk_m__L3_N121(clk_m__L3_N121), 
	.clk_m__L3_N122(clk_m__L3_N122), 
	.clk_m__L3_N123(clk_m__L3_N123), 
	.clk_m__L3_N124(clk_m__L3_N124), 
	.clk_m__L3_N125(clk_m__L3_N125), 
	.clk_m__L3_N126(clk_m__L3_N126), 
	.clk_m__L3_N127(clk_m__L3_N127), 
	.clk_m__L3_N128(clk_m__L3_N128), 
	.clk_m__L3_N129(clk_m__L3_N129), 
	.clk_m__L3_N13(clk_m__L3_N13), 
	.clk_m__L3_N130(clk_m__L3_N130), 
	.clk_m__L3_N131(clk_m__L3_N131), 
	.clk_m__L3_N132(clk_m__L3_N132), 
	.clk_m__L3_N133(clk_m__L3_N133), 
	.clk_m__L3_N134(clk_m__L3_N134), 
	.clk_m__L3_N135(clk_m__L3_N135), 
	.clk_m__L3_N136(clk_m__L3_N136), 
	.clk_m__L3_N137(clk_m__L3_N137), 
	.clk_m__L3_N138(clk_m__L3_N138), 
	.clk_m__L3_N139(clk_m__L3_N139), 
	.clk_m__L3_N14(clk_m__L3_N14), 
	.clk_m__L3_N140(clk_m__L3_N140), 
	.clk_m__L3_N141(clk_m__L3_N141), 
	.clk_m__L3_N142(clk_m__L3_N142), 
	.clk_m__L3_N143(clk_m__L3_N143), 
	.clk_m__L3_N144(clk_m__L3_N144), 
	.clk_m__L3_N145(clk_m__L3_N145), 
	.clk_m__L3_N146(clk_m__L3_N146), 
	.clk_m__L3_N147(clk_m__L3_N147), 
	.clk_m__L3_N148(clk_m__L3_N148), 
	.clk_m__L3_N149(clk_m__L3_N149), 
	.clk_m__L3_N15(clk_m__L3_N15), 
	.clk_m__L3_N150(clk_m__L3_N150), 
	.clk_m__L3_N151(clk_m__L3_N151), 
	.clk_m__L3_N152(clk_m__L3_N152), 
	.clk_m__L3_N153(clk_m__L3_N153), 
	.clk_m__L3_N154(clk_m__L3_N154), 
	.clk_m__L3_N155(clk_m__L3_N155), 
	.clk_m__L3_N156(clk_m__L3_N156), 
	.clk_m__L3_N157(clk_m__L3_N157), 
	.clk_m__L3_N158(clk_m__L3_N158), 
	.clk_m__L3_N159(clk_m__L3_N159), 
	.clk_m__L3_N16(clk_m__L3_N16), 
	.clk_m__L3_N160(clk_m__L3_N160), 
	.clk_m__L3_N161(clk_m__L3_N161), 
	.clk_m__L3_N162(clk_m__L3_N162), 
	.clk_m__L3_N163(clk_m__L3_N163), 
	.clk_m__L3_N164(clk_m__L3_N164), 
	.clk_m__L3_N165(clk_m__L3_N165), 
	.clk_m__L3_N166(clk_m__L3_N166), 
	.clk_m__L3_N167(clk_m__L3_N167), 
	.clk_m__L3_N168(clk_m__L3_N168), 
	.clk_m__L3_N169(clk_m__L3_N169), 
	.clk_m__L3_N17(clk_m__L3_N17), 
	.clk_m__L3_N170(clk_m__L3_N170), 
	.clk_m__L3_N171(clk_m__L3_N171), 
	.clk_m__L3_N172(clk_m__L3_N172), 
	.clk_m__L3_N173(clk_m__L3_N173), 
	.clk_m__L3_N174(clk_m__L3_N174), 
	.clk_m__L3_N175(clk_m__L3_N175), 
	.clk_m__L3_N176(clk_m__L3_N176), 
	.clk_m__L3_N177(clk_m__L3_N177), 
	.clk_m__L3_N18(clk_m__L3_N18), 
	.clk_m__L3_N19(clk_m__L3_N19), 
	.clk_m__L3_N2(clk_m__L3_N2), 
	.clk_m__L3_N20(clk_m__L3_N20), 
	.clk_m__L3_N21(clk_m__L3_N21), 
	.clk_m__L3_N22(clk_m__L3_N22), 
	.clk_m__L3_N23(clk_m__L3_N23), 
	.clk_m__L3_N24(clk_m__L3_N24), 
	.clk_m__L3_N25(clk_m__L3_N25), 
	.clk_m__L3_N26(clk_m__L3_N26), 
	.clk_m__L3_N27(clk_m__L3_N27), 
	.clk_m__L3_N28(clk_m__L3_N28), 
	.clk_m__L3_N29(clk_m__L3_N29), 
	.clk_m__L3_N3(clk_m__L3_N3), 
	.clk_m__L3_N30(clk_m__L3_N30), 
	.clk_m__L3_N31(clk_m__L3_N31), 
	.clk_m__L3_N32(clk_m__L3_N32), 
	.clk_m__L3_N33(clk_m__L3_N33), 
	.clk_m__L3_N34(clk_m__L3_N34), 
	.clk_m__L3_N35(clk_m__L3_N35), 
	.clk_m__L3_N36(clk_m__L3_N36), 
	.clk_m__L3_N37(clk_m__L3_N37), 
	.clk_m__L3_N38(clk_m__L3_N38), 
	.clk_m__L3_N39(clk_m__L3_N39), 
	.clk_m__L3_N4(clk_m__L3_N4), 
	.clk_m__L3_N40(clk_m__L3_N40), 
	.clk_m__L3_N41(clk_m__L3_N41), 
	.clk_m__L3_N42(clk_m__L3_N42), 
	.clk_m__L3_N43(clk_m__L3_N43), 
	.clk_m__L3_N44(clk_m__L3_N44), 
	.clk_m__L3_N45(clk_m__L3_N45), 
	.clk_m__L3_N46(clk_m__L3_N46), 
	.clk_m__L3_N47(clk_m__L3_N47), 
	.clk_m__L3_N48(clk_m__L3_N48), 
	.clk_m__L3_N49(clk_m__L3_N49), 
	.clk_m__L3_N5(clk_m__L3_N5), 
	.clk_m__L3_N50(clk_m__L3_N50), 
	.clk_m__L3_N51(clk_m__L3_N51), 
	.clk_m__L3_N52(clk_m__L3_N52), 
	.clk_m__L3_N53(clk_m__L3_N53), 
	.clk_m__L3_N54(clk_m__L3_N54), 
	.clk_m__L3_N55(clk_m__L3_N55), 
	.clk_m__L3_N56(clk_m__L3_N56), 
	.clk_m__L3_N57(clk_m__L3_N57), 
	.clk_m__L3_N58(clk_m__L3_N58), 
	.clk_m__L3_N59(clk_m__L3_N59), 
	.clk_m__L3_N6(clk_m__L3_N6), 
	.clk_m__L3_N60(clk_m__L3_N60), 
	.clk_m__L3_N61(clk_m__L3_N61), 
	.clk_m__L3_N62(clk_m__L3_N62), 
	.clk_m__L3_N63(clk_m__L3_N63), 
	.clk_m__L3_N64(clk_m__L3_N64), 
	.clk_m__L3_N65(clk_m__L3_N65), 
	.clk_m__L3_N66(clk_m__L3_N66), 
	.clk_m__L3_N67(clk_m__L3_N67), 
	.clk_m__L3_N68(clk_m__L3_N68), 
	.clk_m__L3_N69(clk_m__L3_N69), 
	.clk_m__L3_N7(clk_m__L3_N7), 
	.clk_m__L3_N70(clk_m__L3_N70), 
	.clk_m__L3_N71(clk_m__L3_N71), 
	.clk_m__L3_N72(clk_m__L3_N72), 
	.clk_m__L3_N73(clk_m__L3_N73), 
	.clk_m__L3_N74(clk_m__L3_N74), 
	.clk_m__L3_N75(clk_m__L3_N75), 
	.clk_m__L3_N76(clk_m__L3_N76), 
	.clk_m__L3_N77(clk_m__L3_N77), 
	.clk_m__L3_N78(clk_m__L3_N78), 
	.clk_m__L3_N79(clk_m__L3_N79), 
	.clk_m__L3_N8(clk_m__L3_N8), 
	.clk_m__L3_N80(clk_m__L3_N80), 
	.clk_m__L3_N81(clk_m__L3_N81), 
	.clk_m__L3_N82(clk_m__L3_N82), 
	.clk_m__L3_N83(clk_m__L3_N83), 
	.clk_m__L3_N84(clk_m__L3_N84), 
	.clk_m__L3_N85(clk_m__L3_N85), 
	.clk_m__L3_N86(clk_m__L3_N86), 
	.clk_m__L3_N87(clk_m__L3_N87), 
	.clk_m__L3_N88(clk_m__L3_N88), 
	.clk_m__L3_N89(clk_m__L3_N89), 
	.clk_m__L3_N9(clk_m__L3_N9), 
	.clk_m__L3_N90(clk_m__L3_N90), 
	.clk_m__L3_N91(clk_m__L3_N91), 
	.clk_m__L3_N92(clk_m__L3_N92), 
	.clk_m__L3_N93(clk_m__L3_N93), 
	.clk_m__L3_N94(clk_m__L3_N94), 
	.clk_m__L3_N95(clk_m__L3_N95), 
	.clk_m__L3_N96(clk_m__L3_N96), 
	.clk_m__L3_N97(clk_m__L3_N97), 
	.clk_m__L3_N98(clk_m__L3_N98), 
	.clk_m__L3_N99(clk_m__L3_N99), 
	.clk_m__N0(clk_m__N0));
   TIE1DHD U3 (.O(n2));
   TIE0DHD U4 (.O(n1));
endmodule

