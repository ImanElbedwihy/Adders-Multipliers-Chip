/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu May  6 00:00:30 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1554889499 */

module CLA_adder(A, B, Cin, Sum, Cout, overflow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]Sum;
   output Cout;
   output overflow;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;

   OAI21_X1_LVT i_0_0_0 (.A(n_0_0_2), .B1(n_0_0_3), .B2(n_0_0_1), .ZN(Cout));
   AND2_X1_LVT i_0_0_1 (.A1(n_0_0_1), .A2(n_0_0_0), .ZN(overflow));
   XNOR2_X1_LVT i_0_0_2 (.A(A[31]), .B(n_0_0_3), .ZN(n_0_0_0));
   XOR2_X1_LVT i_0_0_3 (.A(Cin), .B(n_0_0_94), .Z(Sum[0]));
   XNOR2_X1_LVT i_0_0_4 (.A(n_0_0_93), .B(n_0_0_91), .ZN(Sum[1]));
   XNOR2_X1_LVT i_0_0_5 (.A(n_0_0_90), .B(n_0_0_88), .ZN(Sum[2]));
   XNOR2_X1_LVT i_0_0_6 (.A(n_0_0_87), .B(n_0_0_85), .ZN(Sum[3]));
   XNOR2_X1_LVT i_0_0_7 (.A(n_0_0_84), .B(n_0_0_82), .ZN(Sum[4]));
   XNOR2_X1_LVT i_0_0_8 (.A(n_0_0_81), .B(n_0_0_79), .ZN(Sum[5]));
   XNOR2_X1_LVT i_0_0_9 (.A(n_0_0_78), .B(n_0_0_76), .ZN(Sum[6]));
   XNOR2_X1_LVT i_0_0_10 (.A(n_0_0_75), .B(n_0_0_73), .ZN(Sum[7]));
   XNOR2_X1_LVT i_0_0_11 (.A(n_0_0_72), .B(n_0_0_70), .ZN(Sum[8]));
   XNOR2_X1_LVT i_0_0_12 (.A(n_0_0_69), .B(n_0_0_67), .ZN(Sum[9]));
   XNOR2_X1_LVT i_0_0_13 (.A(n_0_0_66), .B(n_0_0_64), .ZN(Sum[10]));
   XNOR2_X1_LVT i_0_0_14 (.A(n_0_0_63), .B(n_0_0_61), .ZN(Sum[11]));
   XNOR2_X1_LVT i_0_0_15 (.A(n_0_0_60), .B(n_0_0_58), .ZN(Sum[12]));
   XNOR2_X1_LVT i_0_0_16 (.A(n_0_0_57), .B(n_0_0_55), .ZN(Sum[13]));
   XNOR2_X1_LVT i_0_0_17 (.A(n_0_0_54), .B(n_0_0_52), .ZN(Sum[14]));
   XNOR2_X1_LVT i_0_0_18 (.A(n_0_0_51), .B(n_0_0_49), .ZN(Sum[15]));
   XNOR2_X1_LVT i_0_0_19 (.A(n_0_0_48), .B(n_0_0_46), .ZN(Sum[16]));
   XNOR2_X1_LVT i_0_0_20 (.A(n_0_0_45), .B(n_0_0_43), .ZN(Sum[17]));
   XNOR2_X1_LVT i_0_0_21 (.A(n_0_0_42), .B(n_0_0_40), .ZN(Sum[18]));
   XNOR2_X1_LVT i_0_0_22 (.A(n_0_0_39), .B(n_0_0_37), .ZN(Sum[19]));
   XNOR2_X1_LVT i_0_0_23 (.A(n_0_0_36), .B(n_0_0_34), .ZN(Sum[20]));
   XNOR2_X1_LVT i_0_0_24 (.A(n_0_0_33), .B(n_0_0_31), .ZN(Sum[21]));
   XNOR2_X1_LVT i_0_0_25 (.A(n_0_0_30), .B(n_0_0_28), .ZN(Sum[22]));
   XNOR2_X1_LVT i_0_0_26 (.A(n_0_0_27), .B(n_0_0_25), .ZN(Sum[23]));
   XNOR2_X1_LVT i_0_0_27 (.A(n_0_0_24), .B(n_0_0_22), .ZN(Sum[24]));
   XNOR2_X1_LVT i_0_0_28 (.A(n_0_0_21), .B(n_0_0_19), .ZN(Sum[25]));
   XNOR2_X1_LVT i_0_0_29 (.A(n_0_0_18), .B(n_0_0_16), .ZN(Sum[26]));
   XNOR2_X1_LVT i_0_0_30 (.A(n_0_0_15), .B(n_0_0_13), .ZN(Sum[27]));
   XNOR2_X1_LVT i_0_0_31 (.A(n_0_0_12), .B(n_0_0_10), .ZN(Sum[28]));
   XNOR2_X1_LVT i_0_0_32 (.A(n_0_0_9), .B(n_0_0_7), .ZN(Sum[29]));
   XNOR2_X1_LVT i_0_0_33 (.A(n_0_0_6), .B(n_0_0_4), .ZN(Sum[30]));
   XOR2_X1_LVT i_0_0_34 (.A(n_0_0_3), .B(n_0_0_1), .Z(Sum[31]));
   OAI21_X1_LVT i_0_0_35 (.A(n_0_0_2), .B1(B[31]), .B2(A[31]), .ZN(n_0_0_1));
   NAND2_X1_LVT i_0_0_36 (.A1(B[31]), .A2(A[31]), .ZN(n_0_0_2));
   AOI22_X1_LVT i_0_0_37 (.A1(B[30]), .A2(A[30]), .B1(n_0_0_5), .B2(n_0_0_4), 
      .ZN(n_0_0_3));
   XOR2_X1_LVT i_0_0_38 (.A(B[30]), .B(A[30]), .Z(n_0_0_4));
   INV_X1_LVT i_0_0_39 (.A(n_0_0_6), .ZN(n_0_0_5));
   AOI22_X1_LVT i_0_0_40 (.A1(B[29]), .A2(A[29]), .B1(n_0_0_8), .B2(n_0_0_7), 
      .ZN(n_0_0_6));
   XOR2_X1_LVT i_0_0_41 (.A(B[29]), .B(A[29]), .Z(n_0_0_7));
   INV_X1_LVT i_0_0_42 (.A(n_0_0_9), .ZN(n_0_0_8));
   AOI22_X1_LVT i_0_0_43 (.A1(B[28]), .A2(A[28]), .B1(n_0_0_11), .B2(n_0_0_10), 
      .ZN(n_0_0_9));
   XOR2_X1_LVT i_0_0_44 (.A(B[28]), .B(A[28]), .Z(n_0_0_10));
   INV_X1_LVT i_0_0_45 (.A(n_0_0_12), .ZN(n_0_0_11));
   AOI22_X1_LVT i_0_0_46 (.A1(B[27]), .A2(A[27]), .B1(n_0_0_14), .B2(n_0_0_13), 
      .ZN(n_0_0_12));
   XOR2_X1_LVT i_0_0_47 (.A(B[27]), .B(A[27]), .Z(n_0_0_13));
   INV_X1_LVT i_0_0_48 (.A(n_0_0_15), .ZN(n_0_0_14));
   AOI22_X1_LVT i_0_0_49 (.A1(B[26]), .A2(A[26]), .B1(n_0_0_17), .B2(n_0_0_16), 
      .ZN(n_0_0_15));
   XOR2_X1_LVT i_0_0_50 (.A(B[26]), .B(A[26]), .Z(n_0_0_16));
   INV_X1_LVT i_0_0_51 (.A(n_0_0_18), .ZN(n_0_0_17));
   AOI22_X1_LVT i_0_0_52 (.A1(B[25]), .A2(A[25]), .B1(n_0_0_20), .B2(n_0_0_19), 
      .ZN(n_0_0_18));
   XOR2_X1_LVT i_0_0_53 (.A(B[25]), .B(A[25]), .Z(n_0_0_19));
   INV_X1_LVT i_0_0_54 (.A(n_0_0_21), .ZN(n_0_0_20));
   AOI22_X1_LVT i_0_0_55 (.A1(B[24]), .A2(A[24]), .B1(n_0_0_23), .B2(n_0_0_22), 
      .ZN(n_0_0_21));
   XOR2_X1_LVT i_0_0_56 (.A(B[24]), .B(A[24]), .Z(n_0_0_22));
   INV_X1_LVT i_0_0_57 (.A(n_0_0_24), .ZN(n_0_0_23));
   AOI22_X1_LVT i_0_0_58 (.A1(B[23]), .A2(A[23]), .B1(n_0_0_26), .B2(n_0_0_25), 
      .ZN(n_0_0_24));
   XOR2_X1_LVT i_0_0_59 (.A(B[23]), .B(A[23]), .Z(n_0_0_25));
   INV_X1_LVT i_0_0_60 (.A(n_0_0_27), .ZN(n_0_0_26));
   AOI22_X1_LVT i_0_0_61 (.A1(B[22]), .A2(A[22]), .B1(n_0_0_29), .B2(n_0_0_28), 
      .ZN(n_0_0_27));
   XOR2_X1_LVT i_0_0_62 (.A(B[22]), .B(A[22]), .Z(n_0_0_28));
   INV_X1_LVT i_0_0_63 (.A(n_0_0_30), .ZN(n_0_0_29));
   AOI22_X1_LVT i_0_0_64 (.A1(B[21]), .A2(A[21]), .B1(n_0_0_32), .B2(n_0_0_31), 
      .ZN(n_0_0_30));
   XOR2_X1_LVT i_0_0_65 (.A(B[21]), .B(A[21]), .Z(n_0_0_31));
   INV_X1_LVT i_0_0_66 (.A(n_0_0_33), .ZN(n_0_0_32));
   AOI22_X1_LVT i_0_0_67 (.A1(B[20]), .A2(A[20]), .B1(n_0_0_35), .B2(n_0_0_34), 
      .ZN(n_0_0_33));
   XOR2_X1_LVT i_0_0_68 (.A(B[20]), .B(A[20]), .Z(n_0_0_34));
   INV_X1_LVT i_0_0_69 (.A(n_0_0_36), .ZN(n_0_0_35));
   AOI22_X1_LVT i_0_0_70 (.A1(B[19]), .A2(A[19]), .B1(n_0_0_38), .B2(n_0_0_37), 
      .ZN(n_0_0_36));
   XOR2_X1_LVT i_0_0_71 (.A(B[19]), .B(A[19]), .Z(n_0_0_37));
   INV_X1_LVT i_0_0_72 (.A(n_0_0_39), .ZN(n_0_0_38));
   AOI22_X1_LVT i_0_0_73 (.A1(B[18]), .A2(A[18]), .B1(n_0_0_41), .B2(n_0_0_40), 
      .ZN(n_0_0_39));
   XOR2_X1_LVT i_0_0_74 (.A(B[18]), .B(A[18]), .Z(n_0_0_40));
   INV_X1_LVT i_0_0_75 (.A(n_0_0_42), .ZN(n_0_0_41));
   AOI22_X1_LVT i_0_0_76 (.A1(B[17]), .A2(A[17]), .B1(n_0_0_44), .B2(n_0_0_43), 
      .ZN(n_0_0_42));
   XOR2_X1_LVT i_0_0_77 (.A(B[17]), .B(A[17]), .Z(n_0_0_43));
   INV_X1_LVT i_0_0_78 (.A(n_0_0_45), .ZN(n_0_0_44));
   AOI22_X1_LVT i_0_0_79 (.A1(B[16]), .A2(A[16]), .B1(n_0_0_47), .B2(n_0_0_46), 
      .ZN(n_0_0_45));
   XOR2_X1_LVT i_0_0_80 (.A(B[16]), .B(A[16]), .Z(n_0_0_46));
   INV_X1_LVT i_0_0_81 (.A(n_0_0_48), .ZN(n_0_0_47));
   AOI22_X1_LVT i_0_0_82 (.A1(B[15]), .A2(A[15]), .B1(n_0_0_50), .B2(n_0_0_49), 
      .ZN(n_0_0_48));
   XOR2_X1_LVT i_0_0_83 (.A(B[15]), .B(A[15]), .Z(n_0_0_49));
   INV_X1_LVT i_0_0_84 (.A(n_0_0_51), .ZN(n_0_0_50));
   AOI22_X1_LVT i_0_0_85 (.A1(B[14]), .A2(A[14]), .B1(n_0_0_53), .B2(n_0_0_52), 
      .ZN(n_0_0_51));
   XOR2_X1_LVT i_0_0_86 (.A(B[14]), .B(A[14]), .Z(n_0_0_52));
   INV_X1_LVT i_0_0_87 (.A(n_0_0_54), .ZN(n_0_0_53));
   AOI22_X1_LVT i_0_0_88 (.A1(B[13]), .A2(A[13]), .B1(n_0_0_56), .B2(n_0_0_55), 
      .ZN(n_0_0_54));
   XOR2_X1_LVT i_0_0_89 (.A(B[13]), .B(A[13]), .Z(n_0_0_55));
   INV_X1_LVT i_0_0_90 (.A(n_0_0_57), .ZN(n_0_0_56));
   AOI22_X1_LVT i_0_0_91 (.A1(B[12]), .A2(A[12]), .B1(n_0_0_59), .B2(n_0_0_58), 
      .ZN(n_0_0_57));
   XOR2_X1_LVT i_0_0_92 (.A(B[12]), .B(A[12]), .Z(n_0_0_58));
   INV_X1_LVT i_0_0_93 (.A(n_0_0_60), .ZN(n_0_0_59));
   AOI22_X1_LVT i_0_0_94 (.A1(B[11]), .A2(A[11]), .B1(n_0_0_62), .B2(n_0_0_61), 
      .ZN(n_0_0_60));
   XOR2_X1_LVT i_0_0_95 (.A(B[11]), .B(A[11]), .Z(n_0_0_61));
   INV_X1_LVT i_0_0_96 (.A(n_0_0_63), .ZN(n_0_0_62));
   AOI22_X1_LVT i_0_0_97 (.A1(B[10]), .A2(A[10]), .B1(n_0_0_65), .B2(n_0_0_64), 
      .ZN(n_0_0_63));
   XOR2_X1_LVT i_0_0_98 (.A(B[10]), .B(A[10]), .Z(n_0_0_64));
   INV_X1_LVT i_0_0_99 (.A(n_0_0_66), .ZN(n_0_0_65));
   AOI22_X1_LVT i_0_0_100 (.A1(B[9]), .A2(A[9]), .B1(n_0_0_68), .B2(n_0_0_67), 
      .ZN(n_0_0_66));
   XOR2_X1_LVT i_0_0_101 (.A(B[9]), .B(A[9]), .Z(n_0_0_67));
   INV_X1_LVT i_0_0_102 (.A(n_0_0_69), .ZN(n_0_0_68));
   AOI22_X1_LVT i_0_0_103 (.A1(B[8]), .A2(A[8]), .B1(n_0_0_71), .B2(n_0_0_70), 
      .ZN(n_0_0_69));
   XOR2_X1_LVT i_0_0_104 (.A(B[8]), .B(A[8]), .Z(n_0_0_70));
   INV_X1_LVT i_0_0_105 (.A(n_0_0_72), .ZN(n_0_0_71));
   AOI22_X1_LVT i_0_0_106 (.A1(B[7]), .A2(A[7]), .B1(n_0_0_74), .B2(n_0_0_73), 
      .ZN(n_0_0_72));
   XOR2_X1_LVT i_0_0_107 (.A(B[7]), .B(A[7]), .Z(n_0_0_73));
   INV_X1_LVT i_0_0_108 (.A(n_0_0_75), .ZN(n_0_0_74));
   AOI22_X1_LVT i_0_0_109 (.A1(B[6]), .A2(A[6]), .B1(n_0_0_77), .B2(n_0_0_76), 
      .ZN(n_0_0_75));
   XOR2_X1_LVT i_0_0_110 (.A(B[6]), .B(A[6]), .Z(n_0_0_76));
   INV_X1_LVT i_0_0_111 (.A(n_0_0_78), .ZN(n_0_0_77));
   AOI22_X1_LVT i_0_0_112 (.A1(B[5]), .A2(A[5]), .B1(n_0_0_80), .B2(n_0_0_79), 
      .ZN(n_0_0_78));
   XOR2_X1_LVT i_0_0_113 (.A(B[5]), .B(A[5]), .Z(n_0_0_79));
   INV_X1_LVT i_0_0_114 (.A(n_0_0_81), .ZN(n_0_0_80));
   AOI22_X1_LVT i_0_0_115 (.A1(B[4]), .A2(A[4]), .B1(n_0_0_83), .B2(n_0_0_82), 
      .ZN(n_0_0_81));
   XOR2_X1_LVT i_0_0_116 (.A(B[4]), .B(A[4]), .Z(n_0_0_82));
   INV_X1_LVT i_0_0_117 (.A(n_0_0_84), .ZN(n_0_0_83));
   AOI22_X1_LVT i_0_0_118 (.A1(B[3]), .A2(A[3]), .B1(n_0_0_86), .B2(n_0_0_85), 
      .ZN(n_0_0_84));
   XOR2_X1_LVT i_0_0_119 (.A(B[3]), .B(A[3]), .Z(n_0_0_85));
   INV_X1_LVT i_0_0_120 (.A(n_0_0_87), .ZN(n_0_0_86));
   AOI22_X1_LVT i_0_0_121 (.A1(B[2]), .A2(A[2]), .B1(n_0_0_89), .B2(n_0_0_88), 
      .ZN(n_0_0_87));
   XOR2_X1_LVT i_0_0_122 (.A(B[2]), .B(A[2]), .Z(n_0_0_88));
   INV_X1_LVT i_0_0_123 (.A(n_0_0_90), .ZN(n_0_0_89));
   AOI22_X1_LVT i_0_0_124 (.A1(B[1]), .A2(A[1]), .B1(n_0_0_92), .B2(n_0_0_91), 
      .ZN(n_0_0_90));
   XOR2_X1_LVT i_0_0_125 (.A(B[1]), .B(A[1]), .Z(n_0_0_91));
   INV_X1_LVT i_0_0_126 (.A(n_0_0_93), .ZN(n_0_0_92));
   AOI22_X1_LVT i_0_0_127 (.A1(B[0]), .A2(A[0]), .B1(Cin), .B2(n_0_0_94), 
      .ZN(n_0_0_93));
   XOR2_X1_LVT i_0_0_128 (.A(B[0]), .B(A[0]), .Z(n_0_0_94));
endmodule
